
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_ALU_N64 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   FUNCRL, FUNCRR);
attribute ENUM_ENCODING of TYPE_OP : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001";
   
   -- Declarations for conversion functions.
   function TYPE_OP_to_std_logic_vector(arg : in TYPE_OP) return 
               std_logic_vector;

end CONV_PACK_ALU_N64;

package body CONV_PACK_ALU_N64 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_to_std_logic_vector(arg : in TYPE_OP) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when FUNCRL => return "1000";
         when FUNCRR => return "1001";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_ALU_N64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_N64.all;

entity ALU_N64_DW01_cmp2_0 is

   port( A, B : in std_logic_vector (63 downto 0);  LEQ, TC : in std_logic;  
         LT_LE, GE_GT : out std_logic);

end ALU_N64_DW01_cmp2_0;

architecture SYN_rpl of ALU_N64_DW01_cmp2_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B(2), ZN => n125);
   U2 : INV_X1 port map( A => n191, ZN => n63);
   U3 : INV_X1 port map( A => B(4), ZN => n123);
   U4 : INV_X1 port map( A => B(3), ZN => n124);
   U5 : INV_X1 port map( A => B(6), ZN => n121);
   U6 : INV_X1 port map( A => B(5), ZN => n122);
   U7 : INV_X1 port map( A => B(8), ZN => n119);
   U8 : INV_X1 port map( A => B(7), ZN => n120);
   U9 : INV_X1 port map( A => B(9), ZN => n118);
   U10 : INV_X1 port map( A => B(10), ZN => n117);
   U11 : INV_X1 port map( A => B(12), ZN => n115);
   U12 : INV_X1 port map( A => B(11), ZN => n116);
   U13 : INV_X1 port map( A => B(14), ZN => n113);
   U14 : INV_X1 port map( A => B(13), ZN => n114);
   U15 : INV_X1 port map( A => B(16), ZN => n111);
   U16 : INV_X1 port map( A => B(15), ZN => n112);
   U17 : INV_X1 port map( A => B(18), ZN => n109);
   U18 : INV_X1 port map( A => B(17), ZN => n110);
   U19 : INV_X1 port map( A => B(20), ZN => n107);
   U20 : INV_X1 port map( A => B(19), ZN => n108);
   U21 : INV_X1 port map( A => B(22), ZN => n105);
   U22 : INV_X1 port map( A => B(21), ZN => n106);
   U23 : INV_X1 port map( A => B(24), ZN => n103);
   U24 : INV_X1 port map( A => B(23), ZN => n104);
   U25 : INV_X1 port map( A => B(26), ZN => n101);
   U26 : INV_X1 port map( A => B(25), ZN => n102);
   U27 : INV_X1 port map( A => B(28), ZN => n99);
   U28 : INV_X1 port map( A => B(27), ZN => n100);
   U29 : INV_X1 port map( A => B(30), ZN => n97);
   U30 : INV_X1 port map( A => B(29), ZN => n98);
   U31 : INV_X1 port map( A => B(32), ZN => n95);
   U32 : INV_X1 port map( A => B(31), ZN => n96);
   U33 : INV_X1 port map( A => B(34), ZN => n93);
   U34 : INV_X1 port map( A => B(33), ZN => n94);
   U35 : INV_X1 port map( A => B(36), ZN => n91);
   U36 : INV_X1 port map( A => B(35), ZN => n92);
   U37 : INV_X1 port map( A => B(38), ZN => n89);
   U38 : INV_X1 port map( A => B(37), ZN => n90);
   U39 : INV_X1 port map( A => B(40), ZN => n87);
   U40 : INV_X1 port map( A => B(39), ZN => n88);
   U41 : INV_X1 port map( A => B(42), ZN => n85);
   U42 : INV_X1 port map( A => B(41), ZN => n86);
   U43 : INV_X1 port map( A => B(44), ZN => n83);
   U44 : INV_X1 port map( A => B(43), ZN => n84);
   U45 : INV_X1 port map( A => B(46), ZN => n81);
   U46 : INV_X1 port map( A => B(45), ZN => n82);
   U47 : INV_X1 port map( A => B(48), ZN => n79);
   U48 : INV_X1 port map( A => B(47), ZN => n80);
   U49 : INV_X1 port map( A => B(50), ZN => n77);
   U50 : INV_X1 port map( A => B(49), ZN => n78);
   U51 : INV_X1 port map( A => B(52), ZN => n75);
   U52 : INV_X1 port map( A => B(51), ZN => n76);
   U53 : INV_X1 port map( A => B(54), ZN => n73);
   U54 : INV_X1 port map( A => B(53), ZN => n74);
   U55 : INV_X1 port map( A => B(56), ZN => n71);
   U56 : INV_X1 port map( A => B(55), ZN => n72);
   U57 : INV_X1 port map( A => B(58), ZN => n69);
   U58 : INV_X1 port map( A => B(57), ZN => n70);
   U59 : INV_X1 port map( A => B(60), ZN => n67);
   U60 : INV_X1 port map( A => B(59), ZN => n68);
   U61 : INV_X1 port map( A => B(61), ZN => n66);
   U62 : INV_X1 port map( A => A(61), ZN => n2);
   U63 : INV_X1 port map( A => B(0), ZN => n126);
   U64 : INV_X1 port map( A => B(63), ZN => n64);
   U65 : INV_X1 port map( A => A(63), ZN => n1);
   U66 : INV_X1 port map( A => B(62), ZN => n65);
   U67 : INV_X1 port map( A => A(2), ZN => n61);
   U68 : INV_X1 port map( A => A(4), ZN => n59);
   U69 : INV_X1 port map( A => A(6), ZN => n57);
   U70 : INV_X1 port map( A => A(8), ZN => n55);
   U71 : INV_X1 port map( A => A(10), ZN => n53);
   U72 : INV_X1 port map( A => A(12), ZN => n51);
   U73 : INV_X1 port map( A => A(14), ZN => n49);
   U74 : INV_X1 port map( A => A(16), ZN => n47);
   U75 : INV_X1 port map( A => A(18), ZN => n45);
   U76 : INV_X1 port map( A => A(20), ZN => n43);
   U77 : INV_X1 port map( A => A(22), ZN => n41);
   U78 : INV_X1 port map( A => A(24), ZN => n39);
   U79 : INV_X1 port map( A => A(26), ZN => n37);
   U80 : INV_X1 port map( A => A(28), ZN => n35);
   U81 : INV_X1 port map( A => A(30), ZN => n33);
   U82 : INV_X1 port map( A => A(32), ZN => n31);
   U83 : INV_X1 port map( A => A(34), ZN => n29);
   U84 : INV_X1 port map( A => A(36), ZN => n27);
   U85 : INV_X1 port map( A => A(38), ZN => n25);
   U86 : INV_X1 port map( A => A(40), ZN => n23);
   U87 : INV_X1 port map( A => A(42), ZN => n21);
   U88 : INV_X1 port map( A => A(44), ZN => n19);
   U89 : INV_X1 port map( A => A(46), ZN => n17);
   U90 : INV_X1 port map( A => A(48), ZN => n15);
   U91 : INV_X1 port map( A => A(50), ZN => n13);
   U92 : INV_X1 port map( A => A(52), ZN => n11);
   U93 : INV_X1 port map( A => A(54), ZN => n9);
   U94 : INV_X1 port map( A => A(56), ZN => n7);
   U95 : INV_X1 port map( A => A(58), ZN => n5);
   U96 : INV_X1 port map( A => A(60), ZN => n3);
   U97 : INV_X1 port map( A => A(1), ZN => n62);
   U98 : INV_X1 port map( A => A(3), ZN => n60);
   U99 : INV_X1 port map( A => A(5), ZN => n58);
   U100 : INV_X1 port map( A => A(7), ZN => n56);
   U101 : INV_X1 port map( A => A(9), ZN => n54);
   U102 : INV_X1 port map( A => A(11), ZN => n52);
   U103 : INV_X1 port map( A => A(13), ZN => n50);
   U104 : INV_X1 port map( A => A(15), ZN => n48);
   U105 : INV_X1 port map( A => A(17), ZN => n46);
   U106 : INV_X1 port map( A => A(19), ZN => n44);
   U107 : INV_X1 port map( A => A(21), ZN => n42);
   U108 : INV_X1 port map( A => A(23), ZN => n40);
   U109 : INV_X1 port map( A => A(25), ZN => n38);
   U110 : INV_X1 port map( A => A(27), ZN => n36);
   U111 : INV_X1 port map( A => A(29), ZN => n34);
   U112 : INV_X1 port map( A => A(31), ZN => n32);
   U113 : INV_X1 port map( A => A(33), ZN => n30);
   U114 : INV_X1 port map( A => A(35), ZN => n28);
   U115 : INV_X1 port map( A => A(37), ZN => n26);
   U116 : INV_X1 port map( A => A(39), ZN => n24);
   U117 : INV_X1 port map( A => A(41), ZN => n22);
   U118 : INV_X1 port map( A => A(43), ZN => n20);
   U119 : INV_X1 port map( A => A(45), ZN => n18);
   U120 : INV_X1 port map( A => A(47), ZN => n16);
   U121 : INV_X1 port map( A => A(49), ZN => n14);
   U122 : INV_X1 port map( A => A(51), ZN => n12);
   U123 : INV_X1 port map( A => A(53), ZN => n10);
   U124 : INV_X1 port map( A => A(55), ZN => n8);
   U125 : INV_X1 port map( A => A(57), ZN => n6);
   U126 : INV_X1 port map( A => A(59), ZN => n4);
   U127 : OAI21_X1 port map( B1 => A(63), B2 => n64, A => n127, ZN => LT_LE);
   U128 : OAI22_X1 port map( A1 => n128, A2 => n129, B1 => B(63), B2 => n1, ZN 
                           => n127);
   U129 : AOI221_X1 port map( B1 => A(62), B2 => n65, C1 => A(61), C2 => n66, A
                           => n130, ZN => n129);
   U130 : AOI221_X1 port map( B1 => B(61), B2 => n2, C1 => B(60), C2 => n3, A 
                           => n131, ZN => n130);
   U131 : AOI221_X1 port map( B1 => A(60), B2 => n67, C1 => A(59), C2 => n68, A
                           => n132, ZN => n131);
   U132 : AOI221_X1 port map( B1 => B(59), B2 => n4, C1 => B(58), C2 => n5, A 
                           => n133, ZN => n132);
   U133 : AOI221_X1 port map( B1 => A(58), B2 => n69, C1 => A(57), C2 => n70, A
                           => n134, ZN => n133);
   U134 : AOI221_X1 port map( B1 => B(57), B2 => n6, C1 => B(56), C2 => n7, A 
                           => n135, ZN => n134);
   U135 : AOI221_X1 port map( B1 => A(56), B2 => n71, C1 => A(55), C2 => n72, A
                           => n136, ZN => n135);
   U136 : AOI221_X1 port map( B1 => B(55), B2 => n8, C1 => B(54), C2 => n9, A 
                           => n137, ZN => n136);
   U137 : AOI221_X1 port map( B1 => A(54), B2 => n73, C1 => A(53), C2 => n74, A
                           => n138, ZN => n137);
   U138 : AOI221_X1 port map( B1 => B(53), B2 => n10, C1 => B(52), C2 => n11, A
                           => n139, ZN => n138);
   U139 : AOI221_X1 port map( B1 => A(52), B2 => n75, C1 => A(51), C2 => n76, A
                           => n140, ZN => n139);
   U140 : AOI221_X1 port map( B1 => B(51), B2 => n12, C1 => B(50), C2 => n13, A
                           => n141, ZN => n140);
   U141 : AOI221_X1 port map( B1 => A(50), B2 => n77, C1 => A(49), C2 => n78, A
                           => n142, ZN => n141);
   U142 : AOI221_X1 port map( B1 => B(49), B2 => n14, C1 => B(48), C2 => n15, A
                           => n143, ZN => n142);
   U143 : AOI221_X1 port map( B1 => A(48), B2 => n79, C1 => A(47), C2 => n80, A
                           => n144, ZN => n143);
   U144 : AOI221_X1 port map( B1 => B(47), B2 => n16, C1 => B(46), C2 => n17, A
                           => n145, ZN => n144);
   U145 : AOI221_X1 port map( B1 => A(46), B2 => n81, C1 => A(45), C2 => n82, A
                           => n146, ZN => n145);
   U146 : AOI221_X1 port map( B1 => B(45), B2 => n18, C1 => B(44), C2 => n19, A
                           => n147, ZN => n146);
   U147 : AOI221_X1 port map( B1 => A(44), B2 => n83, C1 => A(43), C2 => n84, A
                           => n148, ZN => n147);
   U148 : AOI221_X1 port map( B1 => B(43), B2 => n20, C1 => B(42), C2 => n21, A
                           => n149, ZN => n148);
   U149 : AOI221_X1 port map( B1 => A(42), B2 => n85, C1 => A(41), C2 => n86, A
                           => n150, ZN => n149);
   U150 : AOI221_X1 port map( B1 => B(41), B2 => n22, C1 => B(40), C2 => n23, A
                           => n151, ZN => n150);
   U151 : AOI221_X1 port map( B1 => A(40), B2 => n87, C1 => A(39), C2 => n88, A
                           => n152, ZN => n151);
   U152 : AOI221_X1 port map( B1 => B(39), B2 => n24, C1 => B(38), C2 => n25, A
                           => n153, ZN => n152);
   U153 : AOI221_X1 port map( B1 => A(38), B2 => n89, C1 => A(37), C2 => n90, A
                           => n154, ZN => n153);
   U154 : AOI221_X1 port map( B1 => B(37), B2 => n26, C1 => B(36), C2 => n27, A
                           => n155, ZN => n154);
   U155 : AOI221_X1 port map( B1 => A(36), B2 => n91, C1 => A(35), C2 => n92, A
                           => n156, ZN => n155);
   U156 : AOI221_X1 port map( B1 => B(35), B2 => n28, C1 => B(34), C2 => n29, A
                           => n157, ZN => n156);
   U157 : AOI221_X1 port map( B1 => A(34), B2 => n93, C1 => A(33), C2 => n94, A
                           => n158, ZN => n157);
   U158 : AOI221_X1 port map( B1 => B(33), B2 => n30, C1 => B(32), C2 => n31, A
                           => n159, ZN => n158);
   U159 : AOI221_X1 port map( B1 => A(32), B2 => n95, C1 => A(31), C2 => n96, A
                           => n160, ZN => n159);
   U160 : AOI221_X1 port map( B1 => B(31), B2 => n32, C1 => B(30), C2 => n33, A
                           => n161, ZN => n160);
   U161 : AOI221_X1 port map( B1 => A(30), B2 => n97, C1 => A(29), C2 => n98, A
                           => n162, ZN => n161);
   U162 : AOI221_X1 port map( B1 => B(29), B2 => n34, C1 => B(28), C2 => n35, A
                           => n163, ZN => n162);
   U163 : AOI221_X1 port map( B1 => A(28), B2 => n99, C1 => A(27), C2 => n100, 
                           A => n164, ZN => n163);
   U164 : AOI221_X1 port map( B1 => B(27), B2 => n36, C1 => B(26), C2 => n37, A
                           => n165, ZN => n164);
   U165 : AOI221_X1 port map( B1 => A(26), B2 => n101, C1 => A(25), C2 => n102,
                           A => n166, ZN => n165);
   U166 : AOI221_X1 port map( B1 => B(25), B2 => n38, C1 => B(24), C2 => n39, A
                           => n167, ZN => n166);
   U167 : AOI221_X1 port map( B1 => A(24), B2 => n103, C1 => A(23), C2 => n104,
                           A => n168, ZN => n167);
   U168 : AOI221_X1 port map( B1 => B(23), B2 => n40, C1 => B(22), C2 => n41, A
                           => n169, ZN => n168);
   U169 : AOI221_X1 port map( B1 => A(22), B2 => n105, C1 => A(21), C2 => n106,
                           A => n170, ZN => n169);
   U170 : AOI221_X1 port map( B1 => B(21), B2 => n42, C1 => B(20), C2 => n43, A
                           => n171, ZN => n170);
   U171 : AOI221_X1 port map( B1 => A(20), B2 => n107, C1 => A(19), C2 => n108,
                           A => n172, ZN => n171);
   U172 : AOI221_X1 port map( B1 => B(19), B2 => n44, C1 => B(18), C2 => n45, A
                           => n173, ZN => n172);
   U173 : AOI221_X1 port map( B1 => A(18), B2 => n109, C1 => A(17), C2 => n110,
                           A => n174, ZN => n173);
   U174 : AOI221_X1 port map( B1 => B(17), B2 => n46, C1 => B(16), C2 => n47, A
                           => n175, ZN => n174);
   U175 : AOI221_X1 port map( B1 => A(16), B2 => n111, C1 => A(15), C2 => n112,
                           A => n176, ZN => n175);
   U176 : AOI221_X1 port map( B1 => B(15), B2 => n48, C1 => B(14), C2 => n49, A
                           => n177, ZN => n176);
   U177 : AOI221_X1 port map( B1 => A(14), B2 => n113, C1 => A(13), C2 => n114,
                           A => n178, ZN => n177);
   U178 : AOI221_X1 port map( B1 => B(13), B2 => n50, C1 => B(12), C2 => n51, A
                           => n179, ZN => n178);
   U179 : AOI221_X1 port map( B1 => A(12), B2 => n115, C1 => A(11), C2 => n116,
                           A => n180, ZN => n179);
   U180 : AOI221_X1 port map( B1 => B(11), B2 => n52, C1 => B(10), C2 => n53, A
                           => n181, ZN => n180);
   U181 : AOI221_X1 port map( B1 => A(9), B2 => n118, C1 => A(10), C2 => n117, 
                           A => n182, ZN => n181);
   U182 : AOI221_X1 port map( B1 => B(9), B2 => n54, C1 => B(8), C2 => n55, A 
                           => n183, ZN => n182);
   U183 : AOI221_X1 port map( B1 => A(8), B2 => n119, C1 => A(7), C2 => n120, A
                           => n184, ZN => n183);
   U184 : AOI221_X1 port map( B1 => B(7), B2 => n56, C1 => B(6), C2 => n57, A 
                           => n185, ZN => n184);
   U185 : AOI221_X1 port map( B1 => A(6), B2 => n121, C1 => A(5), C2 => n122, A
                           => n186, ZN => n185);
   U186 : AOI221_X1 port map( B1 => B(5), B2 => n58, C1 => B(4), C2 => n59, A 
                           => n187, ZN => n186);
   U187 : AOI221_X1 port map( B1 => A(4), B2 => n123, C1 => A(3), C2 => n124, A
                           => n188, ZN => n187);
   U188 : AOI221_X1 port map( B1 => B(3), B2 => n60, C1 => B(2), C2 => n61, A 
                           => n189, ZN => n188);
   U189 : AOI221_X1 port map( B1 => A(2), B2 => n125, C1 => A(1), C2 => n63, A 
                           => n190, ZN => n189);
   U190 : AOI21_X1 port map( B1 => n191, B2 => n62, A => B(1), ZN => n190);
   U191 : NOR2_X1 port map( A1 => n126, A2 => A(0), ZN => n191);
   U192 : NOR2_X1 port map( A1 => A(62), A2 => n65, ZN => n128);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_N64.all;

entity ALU_N64_DW01_add_0 is

   port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (61 downto 0);  CO : out std_logic);

end ALU_N64_DW01_add_0;

architecture SYN_cla of ALU_N64_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_61_port, SUM_60_port, SUM_59_port, SUM_58_port, SUM_57_port, 
      SUM_56_port, SUM_55_port, SUM_54_port, SUM_53_port, SUM_52_port, 
      SUM_51_port, SUM_50_port, SUM_49_port, SUM_48_port, SUM_47_port, 
      SUM_46_port, SUM_45_port, SUM_44_port, SUM_43_port, SUM_42_port, 
      SUM_41_port, SUM_40_port, SUM_39_port, SUM_38_port, SUM_37_port, 
      SUM_36_port, SUM_35_port, SUM_34_port, SUM_33_port, SUM_32_port, n1, n2, 
      SUM_31_port, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172 : std_logic;

begin
   SUM <= ( SUM_61_port, SUM_60_port, SUM_59_port, SUM_58_port, SUM_57_port, 
      SUM_56_port, SUM_55_port, SUM_54_port, SUM_53_port, SUM_52_port, 
      SUM_51_port, SUM_50_port, SUM_49_port, SUM_48_port, SUM_47_port, 
      SUM_46_port, SUM_45_port, SUM_44_port, SUM_43_port, SUM_42_port, 
      SUM_41_port, SUM_40_port, SUM_39_port, SUM_38_port, SUM_37_port, 
      SUM_36_port, SUM_35_port, SUM_34_port, SUM_33_port, SUM_32_port, 
      SUM_31_port, A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), 
      A(22), A(21), A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), 
      A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1)
      , A(0) );
   
   U2 : OR2_X1 port map( A1 => B(31), A2 => A(31), ZN => n1);
   U3 : OR2_X1 port map( A1 => n105, A2 => n106, ZN => n2);
   U4 : INV_X1 port map( A => n78, ZN => n13);
   U5 : INV_X1 port map( A => n70, ZN => n11);
   U6 : INV_X1 port map( A => n62, ZN => n9);
   U7 : INV_X1 port map( A => n54, ZN => n7);
   U8 : INV_X1 port map( A => n46, ZN => n5);
   U9 : INV_X1 port map( A => n86, ZN => n15);
   U10 : INV_X1 port map( A => n154, ZN => n36);
   U11 : INV_X1 port map( A => n146, ZN => n31);
   U12 : INV_X1 port map( A => n133, ZN => n27);
   U13 : INV_X1 port map( A => n155, ZN => n35);
   U14 : INV_X1 port map( A => n142, ZN => n30);
   U15 : INV_X1 port map( A => n88, ZN => n16);
   U16 : INV_X1 port map( A => n80, ZN => n14);
   U17 : INV_X1 port map( A => n72, ZN => n12);
   U18 : INV_X1 port map( A => n64, ZN => n10);
   U19 : INV_X1 port map( A => n56, ZN => n8);
   U20 : INV_X1 port map( A => n48, ZN => n6);
   U21 : INV_X1 port map( A => n40, ZN => n4);
   U22 : INV_X1 port map( A => n139, ZN => n28);
   U23 : INV_X1 port map( A => n99, ZN => n20);
   U24 : INV_X1 port map( A => n94, ZN => n18);
   U25 : INV_X1 port map( A => n145, ZN => n29);
   U26 : INV_X1 port map( A => n125, ZN => n25);
   U27 : INV_X1 port map( A => n167, ZN => n34);
   U28 : INV_X1 port map( A => n131, ZN => n24);
   U29 : INV_X1 port map( A => n172, ZN => n38);
   U30 : INV_X1 port map( A => n116, ZN => n21);
   U31 : INV_X1 port map( A => n111, ZN => n19);
   U32 : INV_X1 port map( A => n91, ZN => n17);
   U33 : INV_X1 port map( A => n157, ZN => n33);
   U34 : INV_X1 port map( A => n120, ZN => n23);
   U35 : INV_X1 port map( A => n119, ZN => n22);
   U36 : INV_X1 port map( A => n135, ZN => n26);
   U37 : INV_X1 port map( A => n162, ZN => n37);
   U38 : INV_X1 port map( A => n143, ZN => n32);
   U39 : AND2_X1 port map( A1 => n1, A2 => n172, ZN => SUM_31_port);
   U40 : XOR2_X1 port map( A => n39, B => B(61), Z => SUM_61_port);
   U41 : OAI21_X1 port map( B1 => n40, B2 => n41, A => n42, ZN => n39);
   U42 : XOR2_X1 port map( A => n43, B => n41, Z => SUM_60_port);
   U43 : AOI21_X1 port map( B1 => n5, B2 => n44, A => n45, ZN => n41);
   U44 : NAND2_X1 port map( A1 => n4, A2 => n42, ZN => n43);
   U45 : NAND2_X1 port map( A1 => B(60), A2 => A(60), ZN => n42);
   U46 : NOR2_X1 port map( A1 => B(60), A2 => A(60), ZN => n40);
   U47 : XOR2_X1 port map( A => n44, B => n47, Z => SUM_59_port);
   U48 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => n47);
   U49 : NOR2_X1 port map( A1 => B(59), A2 => A(59), ZN => n46);
   U50 : AND2_X1 port map( A1 => B(59), A2 => A(59), ZN => n45);
   U51 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => n44);
   U52 : XOR2_X1 port map( A => n51, B => n49, Z => SUM_58_port);
   U53 : AOI21_X1 port map( B1 => n7, B2 => n52, A => n53, ZN => n49);
   U54 : NAND2_X1 port map( A1 => n6, A2 => n50, ZN => n51);
   U55 : NAND2_X1 port map( A1 => B(58), A2 => A(58), ZN => n50);
   U56 : NOR2_X1 port map( A1 => B(58), A2 => A(58), ZN => n48);
   U57 : XOR2_X1 port map( A => n52, B => n55, Z => SUM_57_port);
   U58 : NOR2_X1 port map( A1 => n53, A2 => n54, ZN => n55);
   U59 : NOR2_X1 port map( A1 => B(57), A2 => A(57), ZN => n54);
   U60 : AND2_X1 port map( A1 => B(57), A2 => A(57), ZN => n53);
   U61 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n52);
   U62 : XOR2_X1 port map( A => n59, B => n57, Z => SUM_56_port);
   U63 : AOI21_X1 port map( B1 => n9, B2 => n60, A => n61, ZN => n57);
   U64 : NAND2_X1 port map( A1 => n8, A2 => n58, ZN => n59);
   U65 : NAND2_X1 port map( A1 => B(56), A2 => A(56), ZN => n58);
   U66 : NOR2_X1 port map( A1 => B(56), A2 => A(56), ZN => n56);
   U67 : XOR2_X1 port map( A => n60, B => n63, Z => SUM_55_port);
   U68 : NOR2_X1 port map( A1 => n61, A2 => n62, ZN => n63);
   U69 : NOR2_X1 port map( A1 => B(55), A2 => A(55), ZN => n62);
   U70 : AND2_X1 port map( A1 => B(55), A2 => A(55), ZN => n61);
   U71 : OAI21_X1 port map( B1 => n64, B2 => n65, A => n66, ZN => n60);
   U72 : XOR2_X1 port map( A => n67, B => n65, Z => SUM_54_port);
   U73 : AOI21_X1 port map( B1 => n11, B2 => n68, A => n69, ZN => n65);
   U74 : NAND2_X1 port map( A1 => n10, A2 => n66, ZN => n67);
   U75 : NAND2_X1 port map( A1 => B(54), A2 => A(54), ZN => n66);
   U76 : NOR2_X1 port map( A1 => B(54), A2 => A(54), ZN => n64);
   U77 : XOR2_X1 port map( A => n68, B => n71, Z => SUM_53_port);
   U78 : NOR2_X1 port map( A1 => n69, A2 => n70, ZN => n71);
   U79 : NOR2_X1 port map( A1 => B(53), A2 => A(53), ZN => n70);
   U80 : AND2_X1 port map( A1 => B(53), A2 => A(53), ZN => n69);
   U81 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n68);
   U82 : XOR2_X1 port map( A => n75, B => n73, Z => SUM_52_port);
   U83 : AOI21_X1 port map( B1 => n13, B2 => n76, A => n77, ZN => n73);
   U84 : NAND2_X1 port map( A1 => n12, A2 => n74, ZN => n75);
   U85 : NAND2_X1 port map( A1 => B(52), A2 => A(52), ZN => n74);
   U86 : NOR2_X1 port map( A1 => B(52), A2 => A(52), ZN => n72);
   U87 : XOR2_X1 port map( A => n76, B => n79, Z => SUM_51_port);
   U88 : NOR2_X1 port map( A1 => n77, A2 => n78, ZN => n79);
   U89 : NOR2_X1 port map( A1 => B(51), A2 => A(51), ZN => n78);
   U90 : AND2_X1 port map( A1 => B(51), A2 => A(51), ZN => n77);
   U91 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => n76);
   U92 : XOR2_X1 port map( A => n83, B => n81, Z => SUM_50_port);
   U93 : AOI21_X1 port map( B1 => n15, B2 => n84, A => n85, ZN => n81);
   U94 : NAND2_X1 port map( A1 => n14, A2 => n82, ZN => n83);
   U95 : NAND2_X1 port map( A1 => B(50), A2 => A(50), ZN => n82);
   U96 : NOR2_X1 port map( A1 => B(50), A2 => A(50), ZN => n80);
   U97 : XOR2_X1 port map( A => n84, B => n87, Z => SUM_49_port);
   U98 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n87);
   U99 : NOR2_X1 port map( A1 => B(49), A2 => A(49), ZN => n86);
   U100 : AND2_X1 port map( A1 => B(49), A2 => A(49), ZN => n85);
   U101 : OAI21_X1 port map( B1 => n88, B2 => n17, A => n89, ZN => n84);
   U102 : XOR2_X1 port map( A => n90, B => n17, Z => SUM_48_port);
   U103 : OAI21_X1 port map( B1 => n92, B2 => n93, A => n94, ZN => n91);
   U104 : AOI21_X1 port map( B1 => n95, B2 => n19, A => n96, ZN => n93);
   U105 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n95);
   U106 : AOI21_X1 port map( B1 => n100, B2 => n21, A => n101, ZN => n98);
   U107 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n22, ZN => n100);
   U108 : AOI221_X1 port map( B1 => n104, B2 => n105, C1 => n106, C2 => n104, A
                           => n107, ZN => n102);
   U109 : NAND2_X1 port map( A1 => n16, A2 => n89, ZN => n90);
   U110 : NAND2_X1 port map( A1 => B(48), A2 => A(48), ZN => n89);
   U111 : NOR2_X1 port map( A1 => B(48), A2 => A(48), ZN => n88);
   U112 : XNOR2_X1 port map( A => n108, B => n109, ZN => SUM_47_port);
   U113 : NOR2_X1 port map( A1 => n18, A2 => n92, ZN => n109);
   U114 : NOR2_X1 port map( A1 => B(47), A2 => A(47), ZN => n92);
   U115 : NAND2_X1 port map( A1 => B(47), A2 => A(47), ZN => n94);
   U116 : AOI21_X1 port map( B1 => n19, B2 => n110, A => n96, ZN => n108);
   U117 : XOR2_X1 port map( A => n110, B => n112, Z => SUM_46_port);
   U118 : NOR2_X1 port map( A1 => n96, A2 => n111, ZN => n112);
   U119 : NOR2_X1 port map( A1 => B(46), A2 => A(46), ZN => n111);
   U120 : AND2_X1 port map( A1 => B(46), A2 => A(46), ZN => n96);
   U121 : OAI21_X1 port map( B1 => n97, B2 => n113, A => n99, ZN => n110);
   U122 : XNOR2_X1 port map( A => n113, B => n114, ZN => SUM_45_port);
   U123 : NOR2_X1 port map( A1 => n20, A2 => n97, ZN => n114);
   U124 : NOR2_X1 port map( A1 => B(45), A2 => A(45), ZN => n97);
   U125 : NAND2_X1 port map( A1 => B(45), A2 => A(45), ZN => n99);
   U126 : AOI21_X1 port map( B1 => n21, B2 => n115, A => n101, ZN => n113);
   U127 : XOR2_X1 port map( A => n115, B => n117, Z => SUM_44_port);
   U128 : NOR2_X1 port map( A1 => n101, A2 => n116, ZN => n117);
   U129 : NOR2_X1 port map( A1 => B(44), A2 => A(44), ZN => n116);
   U130 : AND2_X1 port map( A1 => B(44), A2 => A(44), ZN => n101);
   U131 : OAI21_X1 port map( B1 => n118, B2 => n103, A => n22, ZN => n115);
   U132 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => n119);
   U133 : AOI21_X1 port map( B1 => n123, B2 => n24, A => n124, ZN => n121);
   U134 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n123);
   U135 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n103);
   U136 : XOR2_X1 port map( A => n128, B => n129, Z => SUM_43_port);
   U137 : AOI21_X1 port map( B1 => n130, B2 => n24, A => n124, ZN => n129);
   U138 : NAND2_X1 port map( A1 => n23, A2 => n122, ZN => n128);
   U139 : NAND2_X1 port map( A1 => B(43), A2 => A(43), ZN => n122);
   U140 : NOR2_X1 port map( A1 => B(43), A2 => A(43), ZN => n120);
   U141 : XOR2_X1 port map( A => n130, B => n132, Z => SUM_42_port);
   U142 : NOR2_X1 port map( A1 => n124, A2 => n131, ZN => n132);
   U143 : NOR2_X1 port map( A1 => B(42), A2 => A(42), ZN => n131);
   U144 : AND2_X1 port map( A1 => B(42), A2 => A(42), ZN => n124);
   U145 : OAI21_X1 port map( B1 => n125, B2 => n27, A => n127, ZN => n130);
   U146 : XNOR2_X1 port map( A => n134, B => n133, ZN => SUM_41_port);
   U147 : OAI21_X1 port map( B1 => n135, B2 => n118, A => n126, ZN => n133);
   U148 : NAND2_X1 port map( A1 => n25, A2 => n127, ZN => n134);
   U149 : NAND2_X1 port map( A1 => B(41), A2 => A(41), ZN => n127);
   U150 : NOR2_X1 port map( A1 => B(41), A2 => A(41), ZN => n125);
   U151 : XNOR2_X1 port map( A => n118, B => n136, ZN => SUM_40_port);
   U152 : AND2_X1 port map( A1 => n126, A2 => n26, ZN => n136);
   U153 : NOR2_X1 port map( A1 => B(40), A2 => A(40), ZN => n135);
   U154 : NAND2_X1 port map( A1 => B(40), A2 => A(40), ZN => n126);
   U155 : AOI21_X1 port map( B1 => n2, B2 => n104, A => n107, ZN => n118);
   U156 : OAI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n107);
   U157 : AOI21_X1 port map( B1 => n140, B2 => n29, A => n141, ZN => n138);
   U158 : OAI21_X1 port map( B1 => n142, B2 => n143, A => n144, ZN => n140);
   U159 : NOR4_X1 port map( A1 => n137, A2 => n145, A3 => n142, A4 => n146, ZN 
                           => n104);
   U160 : XNOR2_X1 port map( A => n147, B => n148, ZN => SUM_39_port);
   U161 : NOR2_X1 port map( A1 => n28, A2 => n137, ZN => n148);
   U162 : NOR2_X1 port map( A1 => B(39), A2 => A(39), ZN => n137);
   U163 : NAND2_X1 port map( A1 => B(39), A2 => A(39), ZN => n139);
   U164 : AOI21_X1 port map( B1 => n29, B2 => n149, A => n141, ZN => n147);
   U165 : XOR2_X1 port map( A => n149, B => n150, Z => SUM_38_port);
   U166 : NOR2_X1 port map( A1 => n141, A2 => n145, ZN => n150);
   U167 : NOR2_X1 port map( A1 => B(38), A2 => A(38), ZN => n145);
   U168 : AND2_X1 port map( A1 => B(38), A2 => A(38), ZN => n141);
   U169 : OAI21_X1 port map( B1 => n142, B2 => n151, A => n144, ZN => n149);
   U170 : XOR2_X1 port map( A => n152, B => n151, Z => SUM_37_port);
   U171 : AOI21_X1 port map( B1 => n31, B2 => n2, A => n32, ZN => n151);
   U172 : NAND2_X1 port map( A1 => n30, A2 => n144, ZN => n152);
   U173 : NAND2_X1 port map( A1 => B(37), A2 => A(37), ZN => n144);
   U174 : NOR2_X1 port map( A1 => B(37), A2 => A(37), ZN => n142);
   U175 : XOR2_X1 port map( A => n2, B => n153, Z => SUM_36_port);
   U176 : NOR2_X1 port map( A1 => n32, A2 => n146, ZN => n153);
   U177 : NOR2_X1 port map( A1 => B(36), A2 => A(36), ZN => n146);
   U178 : NAND2_X1 port map( A1 => B(36), A2 => A(36), ZN => n143);
   U179 : NOR4_X1 port map( A1 => n172, A2 => n154, A3 => n155, A4 => n156, ZN 
                           => n106);
   U180 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n156);
   U181 : OAI21_X1 port map( B1 => n157, B2 => n158, A => n159, ZN => n105);
   U182 : AOI21_X1 port map( B1 => n160, B2 => n34, A => n161, ZN => n158);
   U183 : OAI21_X1 port map( B1 => n155, B2 => n162, A => n163, ZN => n160);
   U184 : XOR2_X1 port map( A => n164, B => n165, Z => SUM_35_port);
   U185 : AOI21_X1 port map( B1 => n166, B2 => n34, A => n161, ZN => n165);
   U186 : NAND2_X1 port map( A1 => n33, A2 => n159, ZN => n164);
   U187 : NAND2_X1 port map( A1 => B(35), A2 => A(35), ZN => n159);
   U188 : NOR2_X1 port map( A1 => B(35), A2 => A(35), ZN => n157);
   U189 : XOR2_X1 port map( A => n166, B => n168, Z => SUM_34_port);
   U190 : NOR2_X1 port map( A1 => n161, A2 => n167, ZN => n168);
   U191 : NOR2_X1 port map( A1 => B(34), A2 => A(34), ZN => n167);
   U192 : AND2_X1 port map( A1 => B(34), A2 => A(34), ZN => n161);
   U193 : OAI21_X1 port map( B1 => n155, B2 => n169, A => n163, ZN => n166);
   U194 : XOR2_X1 port map( A => n170, B => n169, Z => SUM_33_port);
   U195 : AOI21_X1 port map( B1 => n36, B2 => n38, A => n37, ZN => n169);
   U196 : NAND2_X1 port map( A1 => n35, A2 => n163, ZN => n170);
   U197 : NAND2_X1 port map( A1 => B(33), A2 => A(33), ZN => n163);
   U198 : NOR2_X1 port map( A1 => B(33), A2 => A(33), ZN => n155);
   U199 : XOR2_X1 port map( A => n38, B => n171, Z => SUM_32_port);
   U200 : NOR2_X1 port map( A1 => n37, A2 => n154, ZN => n171);
   U201 : NOR2_X1 port map( A1 => B(32), A2 => A(32), ZN => n154);
   U202 : NAND2_X1 port map( A1 => B(32), A2 => A(32), ZN => n162);
   U203 : NAND2_X1 port map( A1 => B(31), A2 => A(31), ZN => n172);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_N64.all;

entity ALU_N64_DW02_mult_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (63 downto 0));

end ALU_N64_DW02_mult_0;

architecture SYN_csa of ALU_N64_DW02_mult_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N64_DW01_add_0
      port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (61 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_31_31_port, ab_31_30_port, ab_31_29_port, 
      ab_31_28_port, ab_31_27_port, ab_31_26_port, ab_31_25_port, ab_31_24_port
      , ab_31_23_port, ab_31_22_port, ab_31_21_port, ab_31_20_port, 
      ab_31_19_port, ab_31_18_port, ab_31_17_port, ab_31_16_port, ab_31_15_port
      , ab_31_14_port, ab_31_13_port, ab_31_12_port, ab_31_11_port, 
      ab_31_10_port, ab_31_9_port, ab_31_8_port, ab_31_7_port, ab_31_6_port, 
      ab_31_5_port, ab_31_4_port, ab_31_3_port, ab_31_2_port, ab_31_1_port, 
      ab_31_0_port, ab_30_31_port, ab_30_30_port, ab_30_29_port, ab_30_28_port,
      ab_30_27_port, ab_30_26_port, ab_30_25_port, ab_30_24_port, ab_30_23_port
      , ab_30_22_port, ab_30_21_port, ab_30_20_port, ab_30_19_port, 
      ab_30_18_port, ab_30_17_port, ab_30_16_port, ab_30_15_port, ab_30_14_port
      , ab_30_13_port, ab_30_12_port, ab_30_11_port, ab_30_10_port, 
      ab_30_9_port, ab_30_8_port, ab_30_7_port, ab_30_6_port, ab_30_5_port, 
      ab_30_4_port, ab_30_3_port, ab_30_2_port, ab_30_1_port, ab_30_0_port, 
      ab_29_31_port, ab_29_30_port, ab_29_29_port, ab_29_28_port, ab_29_27_port
      , ab_29_26_port, ab_29_25_port, ab_29_24_port, ab_29_23_port, 
      ab_29_22_port, ab_29_21_port, ab_29_20_port, ab_29_19_port, ab_29_18_port
      , ab_29_17_port, ab_29_16_port, ab_29_15_port, ab_29_14_port, 
      ab_29_13_port, ab_29_12_port, ab_29_11_port, ab_29_10_port, ab_29_9_port,
      ab_29_8_port, ab_29_7_port, ab_29_6_port, ab_29_5_port, ab_29_4_port, 
      ab_29_3_port, ab_29_2_port, ab_29_1_port, ab_29_0_port, ab_28_31_port, 
      ab_28_30_port, ab_28_29_port, ab_28_28_port, ab_28_27_port, ab_28_26_port
      , ab_28_25_port, ab_28_24_port, ab_28_23_port, ab_28_22_port, 
      ab_28_21_port, ab_28_20_port, ab_28_19_port, ab_28_18_port, ab_28_17_port
      , ab_28_16_port, ab_28_15_port, ab_28_14_port, ab_28_13_port, 
      ab_28_12_port, ab_28_11_port, ab_28_10_port, ab_28_9_port, ab_28_8_port, 
      ab_28_7_port, ab_28_6_port, ab_28_5_port, ab_28_4_port, ab_28_3_port, 
      ab_28_2_port, ab_28_1_port, ab_28_0_port, ab_27_31_port, ab_27_30_port, 
      ab_27_29_port, ab_27_28_port, ab_27_27_port, ab_27_26_port, ab_27_25_port
      , ab_27_24_port, ab_27_23_port, ab_27_22_port, ab_27_21_port, 
      ab_27_20_port, ab_27_19_port, ab_27_18_port, ab_27_17_port, ab_27_16_port
      , ab_27_15_port, ab_27_14_port, ab_27_13_port, ab_27_12_port, 
      ab_27_11_port, ab_27_10_port, ab_27_9_port, ab_27_8_port, ab_27_7_port, 
      ab_27_6_port, ab_27_5_port, ab_27_4_port, ab_27_3_port, ab_27_2_port, 
      ab_27_1_port, ab_27_0_port, ab_26_31_port, ab_26_30_port, ab_26_29_port, 
      ab_26_28_port, ab_26_27_port, ab_26_26_port, ab_26_25_port, ab_26_24_port
      , ab_26_23_port, ab_26_22_port, ab_26_21_port, ab_26_20_port, 
      ab_26_19_port, ab_26_18_port, ab_26_17_port, ab_26_16_port, ab_26_15_port
      , ab_26_14_port, ab_26_13_port, ab_26_12_port, ab_26_11_port, 
      ab_26_10_port, ab_26_9_port, ab_26_8_port, ab_26_7_port, ab_26_6_port, 
      ab_26_5_port, ab_26_4_port, ab_26_3_port, ab_26_2_port, ab_26_1_port, 
      ab_26_0_port, ab_25_31_port, ab_25_30_port, ab_25_29_port, ab_25_28_port,
      ab_25_27_port, ab_25_26_port, ab_25_25_port, ab_25_24_port, ab_25_23_port
      , ab_25_22_port, ab_25_21_port, ab_25_20_port, ab_25_19_port, 
      ab_25_18_port, ab_25_17_port, ab_25_16_port, ab_25_15_port, ab_25_14_port
      , ab_25_13_port, ab_25_12_port, ab_25_11_port, ab_25_10_port, 
      ab_25_9_port, ab_25_8_port, ab_25_7_port, ab_25_6_port, ab_25_5_port, 
      ab_25_4_port, ab_25_3_port, ab_25_2_port, ab_25_1_port, ab_25_0_port, 
      ab_24_31_port, ab_24_30_port, ab_24_29_port, ab_24_28_port, ab_24_27_port
      , ab_24_26_port, ab_24_25_port, ab_24_24_port, ab_24_23_port, 
      ab_24_22_port, ab_24_21_port, ab_24_20_port, ab_24_19_port, ab_24_18_port
      , ab_24_17_port, ab_24_16_port, ab_24_15_port, ab_24_14_port, 
      ab_24_13_port, ab_24_12_port, ab_24_11_port, ab_24_10_port, ab_24_9_port,
      ab_24_8_port, ab_24_7_port, ab_24_6_port, ab_24_5_port, ab_24_4_port, 
      ab_24_3_port, ab_24_2_port, ab_24_1_port, ab_24_0_port, ab_23_31_port, 
      ab_23_30_port, ab_23_29_port, ab_23_28_port, ab_23_27_port, ab_23_26_port
      , ab_23_25_port, ab_23_24_port, ab_23_23_port, ab_23_22_port, 
      ab_23_21_port, ab_23_20_port, ab_23_19_port, ab_23_18_port, ab_23_17_port
      , ab_23_16_port, ab_23_15_port, ab_23_14_port, ab_23_13_port, 
      ab_23_12_port, ab_23_11_port, ab_23_10_port, ab_23_9_port, ab_23_8_port, 
      ab_23_7_port, ab_23_6_port, ab_23_5_port, ab_23_4_port, ab_23_3_port, 
      ab_23_2_port, ab_23_1_port, ab_23_0_port, ab_22_31_port, ab_22_30_port, 
      ab_22_29_port, ab_22_28_port, ab_22_27_port, ab_22_26_port, ab_22_25_port
      , ab_22_24_port, ab_22_23_port, ab_22_22_port, ab_22_21_port, 
      ab_22_20_port, ab_22_19_port, ab_22_18_port, ab_22_17_port, ab_22_16_port
      , ab_22_15_port, ab_22_14_port, ab_22_13_port, ab_22_12_port, 
      ab_22_11_port, ab_22_10_port, ab_22_9_port, ab_22_8_port, ab_22_7_port, 
      ab_22_6_port, ab_22_5_port, ab_22_4_port, ab_22_3_port, ab_22_2_port, 
      ab_22_1_port, ab_22_0_port, ab_21_31_port, ab_21_30_port, ab_21_29_port, 
      ab_21_28_port, ab_21_27_port, ab_21_26_port, ab_21_25_port, ab_21_24_port
      , ab_21_23_port, ab_21_22_port, ab_21_21_port, ab_21_20_port, 
      ab_21_19_port, ab_21_18_port, ab_21_17_port, ab_21_16_port, ab_21_15_port
      , ab_21_14_port, ab_21_13_port, ab_21_12_port, ab_21_11_port, 
      ab_21_10_port, ab_21_9_port, ab_21_8_port, ab_21_7_port, ab_21_6_port, 
      ab_21_5_port, ab_21_4_port, ab_21_3_port, ab_21_2_port, ab_21_1_port, 
      ab_21_0_port, ab_20_31_port, ab_20_30_port, ab_20_29_port, ab_20_28_port,
      ab_20_27_port, ab_20_26_port, ab_20_25_port, ab_20_24_port, ab_20_23_port
      , ab_20_22_port, ab_20_21_port, ab_20_20_port, ab_20_19_port, 
      ab_20_18_port, ab_20_17_port, ab_20_16_port, ab_20_15_port, ab_20_14_port
      , ab_20_13_port, ab_20_12_port, ab_20_11_port, ab_20_10_port, 
      ab_20_9_port, ab_20_8_port, ab_20_7_port, ab_20_6_port, ab_20_5_port, 
      ab_20_4_port, ab_20_3_port, ab_20_2_port, ab_20_1_port, ab_20_0_port, 
      ab_19_31_port, ab_19_30_port, ab_19_29_port, ab_19_28_port, ab_19_27_port
      , ab_19_26_port, ab_19_25_port, ab_19_24_port, ab_19_23_port, 
      ab_19_22_port, ab_19_21_port, ab_19_20_port, ab_19_19_port, ab_19_18_port
      , ab_19_17_port, ab_19_16_port, ab_19_15_port, ab_19_14_port, 
      ab_19_13_port, ab_19_12_port, ab_19_11_port, ab_19_10_port, ab_19_9_port,
      ab_19_8_port, ab_19_7_port, ab_19_6_port, ab_19_5_port, ab_19_4_port, 
      ab_19_3_port, ab_19_2_port, ab_19_1_port, ab_19_0_port, ab_18_31_port, 
      ab_18_30_port, ab_18_29_port, ab_18_28_port, ab_18_27_port, ab_18_26_port
      , ab_18_25_port, ab_18_24_port, ab_18_23_port, ab_18_22_port, 
      ab_18_21_port, ab_18_20_port, ab_18_19_port, ab_18_18_port, ab_18_17_port
      , ab_18_16_port, ab_18_15_port, ab_18_14_port, ab_18_13_port, 
      ab_18_12_port, ab_18_11_port, ab_18_10_port, ab_18_9_port, ab_18_8_port, 
      ab_18_7_port, ab_18_6_port, ab_18_5_port, ab_18_4_port, ab_18_3_port, 
      ab_18_2_port, ab_18_1_port, ab_18_0_port, ab_17_31_port, ab_17_30_port, 
      ab_17_29_port, ab_17_28_port, ab_17_27_port, ab_17_26_port, ab_17_25_port
      , ab_17_24_port, ab_17_23_port, ab_17_22_port, ab_17_21_port, 
      ab_17_20_port, ab_17_19_port, ab_17_18_port, ab_17_17_port, ab_17_16_port
      , ab_17_15_port, ab_17_14_port, ab_17_13_port, ab_17_12_port, 
      ab_17_11_port, ab_17_10_port, ab_17_9_port, ab_17_8_port, ab_17_7_port, 
      ab_17_6_port, ab_17_5_port, ab_17_4_port, ab_17_3_port, ab_17_2_port, 
      ab_17_1_port, ab_17_0_port, ab_16_31_port, ab_16_30_port, ab_16_29_port, 
      ab_16_28_port, ab_16_27_port, ab_16_26_port, ab_16_25_port, ab_16_24_port
      , ab_16_23_port, ab_16_22_port, ab_16_21_port, ab_16_20_port, 
      ab_16_19_port, ab_16_18_port, ab_16_17_port, ab_16_16_port, ab_16_15_port
      , ab_16_14_port, ab_16_13_port, ab_16_12_port, ab_16_11_port, 
      ab_16_10_port, ab_16_9_port, ab_16_8_port, ab_16_7_port, ab_16_6_port, 
      ab_16_5_port, ab_16_4_port, ab_16_3_port, ab_16_2_port, ab_16_1_port, 
      ab_16_0_port, ab_15_31_port, ab_15_30_port, ab_15_29_port, ab_15_28_port,
      ab_15_27_port, ab_15_26_port, ab_15_25_port, ab_15_24_port, ab_15_23_port
      , ab_15_22_port, ab_15_21_port, ab_15_20_port, ab_15_19_port, 
      ab_15_18_port, ab_15_17_port, ab_15_16_port, ab_15_15_port, ab_15_14_port
      , ab_15_13_port, ab_15_12_port, ab_15_11_port, ab_15_10_port, 
      ab_15_9_port, ab_15_8_port, ab_15_7_port, ab_15_6_port, ab_15_5_port, 
      ab_15_4_port, ab_15_3_port, ab_15_2_port, ab_15_1_port, ab_15_0_port, 
      ab_14_31_port, ab_14_30_port, ab_14_29_port, ab_14_28_port, ab_14_27_port
      , ab_14_26_port, ab_14_25_port, ab_14_24_port, ab_14_23_port, 
      ab_14_22_port, ab_14_21_port, ab_14_20_port, ab_14_19_port, ab_14_18_port
      , ab_14_17_port, ab_14_16_port, ab_14_15_port, ab_14_14_port, 
      ab_14_13_port, ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port,
      ab_14_8_port, ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, 
      ab_14_3_port, ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_31_port, 
      ab_13_30_port, ab_13_29_port, ab_13_28_port, ab_13_27_port, ab_13_26_port
      , ab_13_25_port, ab_13_24_port, ab_13_23_port, ab_13_22_port, 
      ab_13_21_port, ab_13_20_port, ab_13_19_port, ab_13_18_port, ab_13_17_port
      , ab_13_16_port, ab_13_15_port, ab_13_14_port, ab_13_13_port, 
      ab_13_12_port, ab_13_11_port, ab_13_10_port, ab_13_9_port, ab_13_8_port, 
      ab_13_7_port, ab_13_6_port, ab_13_5_port, ab_13_4_port, ab_13_3_port, 
      ab_13_2_port, ab_13_1_port, ab_13_0_port, ab_12_31_port, ab_12_30_port, 
      ab_12_29_port, ab_12_28_port, ab_12_27_port, ab_12_26_port, ab_12_25_port
      , ab_12_24_port, ab_12_23_port, ab_12_22_port, ab_12_21_port, 
      ab_12_20_port, ab_12_19_port, ab_12_18_port, ab_12_17_port, ab_12_16_port
      , ab_12_15_port, ab_12_14_port, ab_12_13_port, ab_12_12_port, 
      ab_12_11_port, ab_12_10_port, ab_12_9_port, ab_12_8_port, ab_12_7_port, 
      ab_12_6_port, ab_12_5_port, ab_12_4_port, ab_12_3_port, ab_12_2_port, 
      ab_12_1_port, ab_12_0_port, ab_11_31_port, ab_11_30_port, ab_11_29_port, 
      ab_11_28_port, ab_11_27_port, ab_11_26_port, ab_11_25_port, ab_11_24_port
      , ab_11_23_port, ab_11_22_port, ab_11_21_port, ab_11_20_port, 
      ab_11_19_port, ab_11_18_port, ab_11_17_port, ab_11_16_port, ab_11_15_port
      , ab_11_14_port, ab_11_13_port, ab_11_12_port, ab_11_11_port, 
      ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, ab_11_6_port, 
      ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, ab_11_1_port, 
      ab_11_0_port, ab_10_31_port, ab_10_30_port, ab_10_29_port, ab_10_28_port,
      ab_10_27_port, ab_10_26_port, ab_10_25_port, ab_10_24_port, ab_10_23_port
      , ab_10_22_port, ab_10_21_port, ab_10_20_port, ab_10_19_port, 
      ab_10_18_port, ab_10_17_port, ab_10_16_port, ab_10_15_port, ab_10_14_port
      , ab_10_13_port, ab_10_12_port, ab_10_11_port, ab_10_10_port, 
      ab_10_9_port, ab_10_8_port, ab_10_7_port, ab_10_6_port, ab_10_5_port, 
      ab_10_4_port, ab_10_3_port, ab_10_2_port, ab_10_1_port, ab_10_0_port, 
      ab_9_31_port, ab_9_30_port, ab_9_29_port, ab_9_28_port, ab_9_27_port, 
      ab_9_26_port, ab_9_25_port, ab_9_24_port, ab_9_23_port, ab_9_22_port, 
      ab_9_21_port, ab_9_20_port, ab_9_19_port, ab_9_18_port, ab_9_17_port, 
      ab_9_16_port, ab_9_15_port, ab_9_14_port, ab_9_13_port, ab_9_12_port, 
      ab_9_11_port, ab_9_10_port, ab_9_9_port, ab_9_8_port, ab_9_7_port, 
      ab_9_6_port, ab_9_5_port, ab_9_4_port, ab_9_3_port, ab_9_2_port, 
      ab_9_1_port, ab_9_0_port, ab_8_31_port, ab_8_30_port, ab_8_29_port, 
      ab_8_28_port, ab_8_27_port, ab_8_26_port, ab_8_25_port, ab_8_24_port, 
      ab_8_23_port, ab_8_22_port, ab_8_21_port, ab_8_20_port, ab_8_19_port, 
      ab_8_18_port, ab_8_17_port, ab_8_16_port, ab_8_15_port, ab_8_14_port, 
      ab_8_13_port, ab_8_12_port, ab_8_11_port, ab_8_10_port, ab_8_9_port, 
      ab_8_8_port, ab_8_7_port, ab_8_6_port, ab_8_5_port, ab_8_4_port, 
      ab_8_3_port, ab_8_2_port, ab_8_1_port, ab_8_0_port, ab_7_31_port, 
      ab_7_30_port, ab_7_29_port, ab_7_28_port, ab_7_27_port, ab_7_26_port, 
      ab_7_25_port, ab_7_24_port, ab_7_23_port, ab_7_22_port, ab_7_21_port, 
      ab_7_20_port, ab_7_19_port, ab_7_18_port, ab_7_17_port, ab_7_16_port, 
      ab_7_15_port, ab_7_14_port, ab_7_13_port, ab_7_12_port, ab_7_11_port, 
      ab_7_10_port, ab_7_9_port, ab_7_8_port, ab_7_7_port, ab_7_6_port, 
      ab_7_5_port, ab_7_4_port, ab_7_3_port, ab_7_2_port, ab_7_1_port, 
      ab_7_0_port, ab_6_31_port, ab_6_30_port, ab_6_29_port, ab_6_28_port, 
      ab_6_27_port, ab_6_26_port, ab_6_25_port, ab_6_24_port, ab_6_23_port, 
      ab_6_22_port, ab_6_21_port, ab_6_20_port, ab_6_19_port, ab_6_18_port, 
      ab_6_17_port, ab_6_16_port, ab_6_15_port, ab_6_14_port, ab_6_13_port, 
      ab_6_12_port, ab_6_11_port, ab_6_10_port, ab_6_9_port, ab_6_8_port, 
      ab_6_7_port, ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, 
      ab_6_2_port, ab_6_1_port, ab_6_0_port, ab_5_31_port, ab_5_30_port, 
      ab_5_29_port, ab_5_28_port, ab_5_27_port, ab_5_26_port, ab_5_25_port, 
      ab_5_24_port, ab_5_23_port, ab_5_22_port, ab_5_21_port, ab_5_20_port, 
      ab_5_19_port, ab_5_18_port, ab_5_17_port, ab_5_16_port, ab_5_15_port, 
      ab_5_14_port, ab_5_13_port, ab_5_12_port, ab_5_11_port, ab_5_10_port, 
      ab_5_9_port, ab_5_8_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_31_port, ab_4_30_port, ab_4_29_port, ab_4_28_port, ab_4_27_port, 
      ab_4_26_port, ab_4_25_port, ab_4_24_port, ab_4_23_port, ab_4_22_port, 
      ab_4_21_port, ab_4_20_port, ab_4_19_port, ab_4_18_port, ab_4_17_port, 
      ab_4_16_port, ab_4_15_port, ab_4_14_port, ab_4_13_port, ab_4_12_port, 
      ab_4_11_port, ab_4_10_port, ab_4_9_port, ab_4_8_port, ab_4_7_port, 
      ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, ab_4_2_port, 
      ab_4_1_port, ab_4_0_port, ab_3_31_port, ab_3_30_port, ab_3_29_port, 
      ab_3_28_port, ab_3_27_port, ab_3_26_port, ab_3_25_port, ab_3_24_port, 
      ab_3_23_port, ab_3_22_port, ab_3_21_port, ab_3_20_port, ab_3_19_port, 
      ab_3_18_port, ab_3_17_port, ab_3_16_port, ab_3_15_port, ab_3_14_port, 
      ab_3_13_port, ab_3_12_port, ab_3_11_port, ab_3_10_port, ab_3_9_port, 
      ab_3_8_port, ab_3_7_port, ab_3_6_port, ab_3_5_port, ab_3_4_port, 
      ab_3_3_port, ab_3_2_port, ab_3_1_port, ab_3_0_port, ab_2_31_port, 
      ab_2_30_port, ab_2_29_port, ab_2_28_port, ab_2_27_port, ab_2_26_port, 
      ab_2_25_port, ab_2_24_port, ab_2_23_port, ab_2_22_port, ab_2_21_port, 
      ab_2_20_port, ab_2_19_port, ab_2_18_port, ab_2_17_port, ab_2_16_port, 
      ab_2_15_port, ab_2_14_port, ab_2_13_port, ab_2_12_port, ab_2_11_port, 
      ab_2_10_port, ab_2_9_port, ab_2_8_port, ab_2_7_port, ab_2_6_port, 
      ab_2_5_port, ab_2_4_port, ab_2_3_port, ab_2_2_port, ab_2_1_port, 
      ab_2_0_port, ab_1_31_port, ab_1_30_port, ab_1_29_port, ab_1_28_port, 
      ab_1_27_port, ab_1_26_port, ab_1_25_port, ab_1_24_port, ab_1_23_port, 
      ab_1_22_port, ab_1_21_port, ab_1_20_port, ab_1_19_port, ab_1_18_port, 
      ab_1_17_port, ab_1_16_port, ab_1_15_port, ab_1_14_port, ab_1_13_port, 
      ab_1_12_port, ab_1_11_port, ab_1_10_port, ab_1_9_port, ab_1_8_port, 
      ab_1_7_port, ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, 
      ab_1_2_port, ab_1_1_port, ab_1_0_port, ab_0_31_port, ab_0_30_port, 
      ab_0_29_port, ab_0_28_port, ab_0_27_port, ab_0_26_port, ab_0_25_port, 
      ab_0_24_port, ab_0_23_port, ab_0_22_port, ab_0_21_port, ab_0_20_port, 
      ab_0_19_port, ab_0_18_port, ab_0_17_port, ab_0_16_port, ab_0_15_port, 
      ab_0_14_port, ab_0_13_port, ab_0_12_port, ab_0_11_port, ab_0_10_port, 
      ab_0_9_port, ab_0_8_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_15_30_port, 
      CARRYB_15_29_port, CARRYB_15_28_port, CARRYB_15_27_port, 
      CARRYB_15_26_port, CARRYB_15_25_port, CARRYB_15_24_port, 
      CARRYB_15_23_port, CARRYB_15_22_port, CARRYB_15_21_port, 
      CARRYB_15_20_port, CARRYB_15_19_port, CARRYB_15_18_port, 
      CARRYB_15_17_port, CARRYB_15_16_port, CARRYB_15_15_port, 
      CARRYB_15_14_port, CARRYB_15_13_port, CARRYB_15_12_port, 
      CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port, CARRYB_15_8_port,
      CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port, CARRYB_15_4_port, 
      CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_1_port, CARRYB_15_0_port, 
      CARRYB_14_30_port, CARRYB_14_29_port, CARRYB_14_28_port, 
      CARRYB_14_27_port, CARRYB_14_26_port, CARRYB_14_25_port, 
      CARRYB_14_24_port, CARRYB_14_23_port, CARRYB_14_22_port, 
      CARRYB_14_21_port, CARRYB_14_20_port, CARRYB_14_19_port, 
      CARRYB_14_18_port, CARRYB_14_17_port, CARRYB_14_16_port, 
      CARRYB_14_15_port, CARRYB_14_14_port, CARRYB_14_13_port, 
      CARRYB_14_12_port, CARRYB_14_11_port, CARRYB_14_10_port, CARRYB_14_9_port
      , CARRYB_14_8_port, CARRYB_14_7_port, CARRYB_14_6_port, CARRYB_14_5_port,
      CARRYB_14_4_port, CARRYB_14_3_port, CARRYB_14_2_port, CARRYB_14_1_port, 
      CARRYB_14_0_port, CARRYB_13_30_port, CARRYB_13_29_port, CARRYB_13_28_port
      , CARRYB_13_27_port, CARRYB_13_26_port, CARRYB_13_25_port, 
      CARRYB_13_24_port, CARRYB_13_23_port, CARRYB_13_22_port, 
      CARRYB_13_21_port, CARRYB_13_20_port, CARRYB_13_19_port, 
      CARRYB_13_18_port, CARRYB_13_17_port, CARRYB_13_16_port, 
      CARRYB_13_15_port, CARRYB_13_14_port, CARRYB_13_13_port, 
      CARRYB_13_12_port, CARRYB_13_11_port, CARRYB_13_10_port, CARRYB_13_9_port
      , CARRYB_13_8_port, CARRYB_13_7_port, CARRYB_13_6_port, CARRYB_13_5_port,
      CARRYB_13_4_port, CARRYB_13_3_port, CARRYB_13_2_port, CARRYB_13_1_port, 
      CARRYB_13_0_port, CARRYB_12_30_port, CARRYB_12_29_port, CARRYB_12_28_port
      , CARRYB_12_27_port, CARRYB_12_26_port, CARRYB_12_25_port, 
      CARRYB_12_24_port, CARRYB_12_23_port, CARRYB_12_22_port, 
      CARRYB_12_21_port, CARRYB_12_20_port, CARRYB_12_19_port, 
      CARRYB_12_18_port, CARRYB_12_17_port, CARRYB_12_16_port, 
      CARRYB_12_15_port, CARRYB_12_14_port, CARRYB_12_13_port, 
      CARRYB_12_12_port, CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port
      , CARRYB_12_8_port, CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port,
      CARRYB_12_4_port, CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, 
      CARRYB_12_0_port, CARRYB_11_30_port, CARRYB_11_29_port, CARRYB_11_28_port
      , CARRYB_11_27_port, CARRYB_11_26_port, CARRYB_11_25_port, 
      CARRYB_11_24_port, CARRYB_11_23_port, CARRYB_11_22_port, 
      CARRYB_11_21_port, CARRYB_11_20_port, CARRYB_11_19_port, 
      CARRYB_11_18_port, CARRYB_11_17_port, CARRYB_11_16_port, 
      CARRYB_11_15_port, CARRYB_11_14_port, CARRYB_11_13_port, 
      CARRYB_11_12_port, CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port
      , CARRYB_11_8_port, CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_5_port,
      CARRYB_11_4_port, CARRYB_11_3_port, CARRYB_11_2_port, CARRYB_11_1_port, 
      CARRYB_11_0_port, CARRYB_10_30_port, CARRYB_10_29_port, CARRYB_10_28_port
      , CARRYB_10_27_port, CARRYB_10_26_port, CARRYB_10_25_port, 
      CARRYB_10_24_port, CARRYB_10_23_port, CARRYB_10_22_port, 
      CARRYB_10_21_port, CARRYB_10_20_port, CARRYB_10_19_port, 
      CARRYB_10_18_port, CARRYB_10_17_port, CARRYB_10_16_port, 
      CARRYB_10_15_port, CARRYB_10_14_port, CARRYB_10_13_port, 
      CARRYB_10_12_port, CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port
      , CARRYB_10_8_port, CARRYB_10_7_port, CARRYB_10_6_port, CARRYB_10_5_port,
      CARRYB_10_4_port, CARRYB_10_3_port, CARRYB_10_2_port, CARRYB_10_1_port, 
      CARRYB_10_0_port, CARRYB_9_30_port, CARRYB_9_29_port, CARRYB_9_28_port, 
      CARRYB_9_27_port, CARRYB_9_26_port, CARRYB_9_25_port, CARRYB_9_24_port, 
      CARRYB_9_23_port, CARRYB_9_22_port, CARRYB_9_21_port, CARRYB_9_20_port, 
      CARRYB_9_19_port, CARRYB_9_18_port, CARRYB_9_17_port, CARRYB_9_16_port, 
      CARRYB_9_15_port, CARRYB_9_14_port, CARRYB_9_13_port, CARRYB_9_12_port, 
      CARRYB_9_11_port, CARRYB_9_10_port, CARRYB_9_9_port, CARRYB_9_8_port, 
      CARRYB_9_7_port, CARRYB_9_6_port, CARRYB_9_5_port, CARRYB_9_4_port, 
      CARRYB_9_3_port, CARRYB_9_2_port, CARRYB_9_1_port, CARRYB_9_0_port, 
      CARRYB_8_30_port, CARRYB_8_29_port, CARRYB_8_28_port, CARRYB_8_27_port, 
      CARRYB_8_26_port, CARRYB_8_25_port, CARRYB_8_24_port, CARRYB_8_23_port, 
      CARRYB_8_22_port, CARRYB_8_21_port, CARRYB_8_20_port, CARRYB_8_19_port, 
      CARRYB_8_18_port, CARRYB_8_17_port, CARRYB_8_16_port, CARRYB_8_15_port, 
      CARRYB_8_14_port, CARRYB_8_13_port, CARRYB_8_12_port, CARRYB_8_11_port, 
      CARRYB_8_10_port, CARRYB_8_9_port, CARRYB_8_8_port, CARRYB_8_7_port, 
      CARRYB_8_6_port, CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, 
      CARRYB_8_2_port, CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_30_port, 
      CARRYB_7_29_port, CARRYB_7_28_port, CARRYB_7_27_port, CARRYB_7_26_port, 
      CARRYB_7_25_port, CARRYB_7_24_port, CARRYB_7_23_port, CARRYB_7_22_port, 
      CARRYB_7_21_port, CARRYB_7_20_port, CARRYB_7_19_port, CARRYB_7_18_port, 
      CARRYB_7_17_port, CARRYB_7_16_port, CARRYB_7_15_port, CARRYB_7_14_port, 
      CARRYB_7_13_port, CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, 
      CARRYB_7_9_port, CARRYB_7_8_port, CARRYB_7_7_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_30_port, CARRYB_6_29_port, 
      CARRYB_6_28_port, CARRYB_6_27_port, CARRYB_6_26_port, CARRYB_6_25_port, 
      CARRYB_6_24_port, CARRYB_6_23_port, CARRYB_6_22_port, CARRYB_6_21_port, 
      CARRYB_6_20_port, CARRYB_6_19_port, CARRYB_6_18_port, CARRYB_6_17_port, 
      CARRYB_6_16_port, CARRYB_6_15_port, CARRYB_6_14_port, CARRYB_6_13_port, 
      CARRYB_6_12_port, CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, 
      CARRYB_6_8_port, CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_30_port, CARRYB_5_29_port, CARRYB_5_28_port, 
      CARRYB_5_27_port, CARRYB_5_26_port, CARRYB_5_25_port, CARRYB_5_24_port, 
      CARRYB_5_23_port, CARRYB_5_22_port, CARRYB_5_21_port, CARRYB_5_20_port, 
      CARRYB_5_19_port, CARRYB_5_18_port, CARRYB_5_17_port, CARRYB_5_16_port, 
      CARRYB_5_15_port, CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, 
      CARRYB_5_11_port, CARRYB_5_10_port, CARRYB_5_9_port, CARRYB_5_8_port, 
      CARRYB_5_7_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_30_port, CARRYB_4_29_port, CARRYB_4_28_port, CARRYB_4_27_port, 
      CARRYB_4_26_port, CARRYB_4_25_port, CARRYB_4_24_port, CARRYB_4_23_port, 
      CARRYB_4_22_port, CARRYB_4_21_port, CARRYB_4_20_port, CARRYB_4_19_port, 
      CARRYB_4_18_port, CARRYB_4_17_port, CARRYB_4_16_port, CARRYB_4_15_port, 
      CARRYB_4_14_port, CARRYB_4_13_port, CARRYB_4_12_port, CARRYB_4_11_port, 
      CARRYB_4_10_port, CARRYB_4_9_port, CARRYB_4_8_port, CARRYB_4_7_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_30_port, 
      CARRYB_3_29_port, CARRYB_3_28_port, CARRYB_3_27_port, CARRYB_3_26_port, 
      CARRYB_3_25_port, CARRYB_3_24_port, CARRYB_3_23_port, CARRYB_3_22_port, 
      CARRYB_3_21_port, CARRYB_3_20_port, CARRYB_3_19_port, CARRYB_3_18_port, 
      CARRYB_3_17_port, CARRYB_3_16_port, CARRYB_3_15_port, CARRYB_3_14_port, 
      CARRYB_3_13_port, CARRYB_3_12_port, CARRYB_3_11_port, CARRYB_3_10_port, 
      CARRYB_3_9_port, CARRYB_3_8_port, CARRYB_3_7_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_30_port, CARRYB_2_29_port, 
      CARRYB_2_28_port, CARRYB_2_27_port, CARRYB_2_26_port, CARRYB_2_25_port, 
      CARRYB_2_24_port, CARRYB_2_23_port, CARRYB_2_22_port, CARRYB_2_21_port, 
      CARRYB_2_20_port, CARRYB_2_19_port, CARRYB_2_18_port, CARRYB_2_17_port, 
      CARRYB_2_16_port, CARRYB_2_15_port, CARRYB_2_14_port, CARRYB_2_13_port, 
      CARRYB_2_12_port, CARRYB_2_11_port, CARRYB_2_10_port, CARRYB_2_9_port, 
      CARRYB_2_8_port, CARRYB_2_7_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_15_30_port, SUMB_15_29_port, SUMB_15_28_port, 
      SUMB_15_27_port, SUMB_15_26_port, SUMB_15_25_port, SUMB_15_24_port, 
      SUMB_15_23_port, SUMB_15_22_port, SUMB_15_21_port, SUMB_15_20_port, 
      SUMB_15_19_port, SUMB_15_18_port, SUMB_15_17_port, SUMB_15_16_port, 
      SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, SUMB_15_12_port, 
      SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, SUMB_15_8_port, 
      SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, SUMB_15_4_port, 
      SUMB_15_3_port, SUMB_15_2_port, SUMB_15_1_port, SUMB_14_30_port, 
      SUMB_14_29_port, SUMB_14_28_port, SUMB_14_27_port, SUMB_14_26_port, 
      SUMB_14_25_port, SUMB_14_24_port, SUMB_14_23_port, SUMB_14_22_port, 
      SUMB_14_21_port, SUMB_14_20_port, SUMB_14_19_port, SUMB_14_18_port, 
      SUMB_14_17_port, SUMB_14_16_port, SUMB_14_15_port, SUMB_14_14_port, 
      SUMB_14_13_port, SUMB_14_12_port, SUMB_14_11_port, SUMB_14_10_port, 
      SUMB_14_9_port, SUMB_14_8_port, SUMB_14_7_port, SUMB_14_6_port, 
      SUMB_14_5_port, SUMB_14_4_port, SUMB_14_3_port, SUMB_14_2_port, 
      SUMB_14_1_port, SUMB_13_30_port, SUMB_13_29_port, SUMB_13_28_port, 
      SUMB_13_27_port, SUMB_13_26_port, SUMB_13_25_port, SUMB_13_24_port, 
      SUMB_13_23_port, SUMB_13_22_port, SUMB_13_21_port, SUMB_13_20_port, 
      SUMB_13_19_port, SUMB_13_18_port, SUMB_13_17_port, SUMB_13_16_port, 
      SUMB_13_15_port, SUMB_13_14_port, SUMB_13_13_port, SUMB_13_12_port, 
      SUMB_13_11_port, SUMB_13_10_port, SUMB_13_9_port, SUMB_13_8_port, 
      SUMB_13_7_port, SUMB_13_6_port, SUMB_13_5_port, SUMB_13_4_port, 
      SUMB_13_3_port, SUMB_13_2_port, SUMB_13_1_port, SUMB_12_30_port, 
      SUMB_12_29_port, SUMB_12_28_port, SUMB_12_27_port, SUMB_12_26_port, 
      SUMB_12_25_port, SUMB_12_24_port, SUMB_12_23_port, SUMB_12_22_port, 
      SUMB_12_21_port, SUMB_12_20_port, SUMB_12_19_port, SUMB_12_18_port, 
      SUMB_12_17_port, SUMB_12_16_port, SUMB_12_15_port, SUMB_12_14_port, 
      SUMB_12_13_port, SUMB_12_12_port, SUMB_12_11_port, SUMB_12_10_port, 
      SUMB_12_9_port, SUMB_12_8_port, SUMB_12_7_port, SUMB_12_6_port, 
      SUMB_12_5_port, SUMB_12_4_port, SUMB_12_3_port, SUMB_12_2_port, 
      SUMB_12_1_port, SUMB_11_30_port, SUMB_11_29_port, SUMB_11_28_port, 
      SUMB_11_27_port, SUMB_11_26_port, SUMB_11_25_port, SUMB_11_24_port, 
      SUMB_11_23_port, SUMB_11_22_port, SUMB_11_21_port, SUMB_11_20_port, 
      SUMB_11_19_port, SUMB_11_18_port, SUMB_11_17_port, SUMB_11_16_port, 
      SUMB_11_15_port, SUMB_11_14_port, SUMB_11_13_port, SUMB_11_12_port, 
      SUMB_11_11_port, SUMB_11_10_port, SUMB_11_9_port, SUMB_11_8_port, 
      SUMB_11_7_port, SUMB_11_6_port, SUMB_11_5_port, SUMB_11_4_port, 
      SUMB_11_3_port, SUMB_11_2_port, SUMB_11_1_port, SUMB_10_30_port, 
      SUMB_10_29_port, SUMB_10_28_port, SUMB_10_27_port, SUMB_10_26_port, 
      SUMB_10_25_port, SUMB_10_24_port, SUMB_10_23_port, SUMB_10_22_port, 
      SUMB_10_21_port, SUMB_10_20_port, SUMB_10_19_port, SUMB_10_18_port, 
      SUMB_10_17_port, SUMB_10_16_port, SUMB_10_15_port, SUMB_10_14_port, 
      SUMB_10_13_port, SUMB_10_12_port, SUMB_10_11_port, SUMB_10_10_port, 
      SUMB_10_9_port, SUMB_10_8_port, SUMB_10_7_port, SUMB_10_6_port, 
      SUMB_10_5_port, SUMB_10_4_port, SUMB_10_3_port, SUMB_10_2_port, 
      SUMB_10_1_port, SUMB_9_30_port, SUMB_9_29_port, SUMB_9_28_port, 
      SUMB_9_27_port, SUMB_9_26_port, SUMB_9_25_port, SUMB_9_24_port, 
      SUMB_9_23_port, SUMB_9_22_port, SUMB_9_21_port, SUMB_9_20_port, 
      SUMB_9_19_port, SUMB_9_18_port, SUMB_9_17_port, SUMB_9_16_port, 
      SUMB_9_15_port, SUMB_9_14_port, SUMB_9_13_port, SUMB_9_12_port, 
      SUMB_9_11_port, SUMB_9_10_port, SUMB_9_9_port, SUMB_9_8_port, 
      SUMB_9_7_port, SUMB_9_6_port, SUMB_9_5_port, SUMB_9_4_port, SUMB_9_3_port
      , SUMB_9_2_port, SUMB_9_1_port, SUMB_8_30_port, SUMB_8_29_port, 
      SUMB_8_28_port, SUMB_8_27_port, SUMB_8_26_port, SUMB_8_25_port, 
      SUMB_8_24_port, SUMB_8_23_port, SUMB_8_22_port, SUMB_8_21_port, 
      SUMB_8_20_port, SUMB_8_19_port, SUMB_8_18_port, SUMB_8_17_port, 
      SUMB_8_16_port, SUMB_8_15_port, SUMB_8_14_port, SUMB_8_13_port, 
      SUMB_8_12_port, SUMB_8_11_port, SUMB_8_10_port, SUMB_8_9_port, 
      SUMB_8_8_port, SUMB_8_7_port, SUMB_8_6_port, SUMB_8_5_port, SUMB_8_4_port
      , SUMB_8_3_port, SUMB_8_2_port, SUMB_8_1_port, SUMB_7_30_port, 
      SUMB_7_29_port, SUMB_7_28_port, SUMB_7_27_port, SUMB_7_26_port, 
      SUMB_7_25_port, SUMB_7_24_port, SUMB_7_23_port, SUMB_7_22_port, 
      SUMB_7_21_port, SUMB_7_20_port, SUMB_7_19_port, SUMB_7_18_port, 
      SUMB_7_17_port, SUMB_7_16_port, SUMB_7_15_port, SUMB_7_14_port, 
      SUMB_7_13_port, SUMB_7_12_port, SUMB_7_11_port, SUMB_7_10_port, 
      SUMB_7_9_port, SUMB_7_8_port, SUMB_7_7_port, SUMB_7_6_port, SUMB_7_5_port
      , SUMB_7_4_port, SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, 
      SUMB_6_30_port, SUMB_6_29_port, SUMB_6_28_port, SUMB_6_27_port, 
      SUMB_6_26_port, SUMB_6_25_port, SUMB_6_24_port, SUMB_6_23_port, 
      SUMB_6_22_port, SUMB_6_21_port, SUMB_6_20_port, SUMB_6_19_port, 
      SUMB_6_18_port, SUMB_6_17_port, SUMB_6_16_port, SUMB_6_15_port, 
      SUMB_6_14_port, SUMB_6_13_port, SUMB_6_12_port, SUMB_6_11_port, 
      SUMB_6_10_port, SUMB_6_9_port, SUMB_6_8_port, SUMB_6_7_port, 
      SUMB_6_6_port, SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port
      , SUMB_6_1_port, SUMB_5_30_port, SUMB_5_29_port, SUMB_5_28_port, 
      SUMB_5_27_port, SUMB_5_26_port, SUMB_5_25_port, SUMB_5_24_port, 
      SUMB_5_23_port, SUMB_5_22_port, SUMB_5_21_port, SUMB_5_20_port, 
      SUMB_5_19_port, SUMB_5_18_port, SUMB_5_17_port, SUMB_5_16_port, 
      SUMB_5_15_port, SUMB_5_14_port, SUMB_5_13_port, SUMB_5_12_port, 
      SUMB_5_11_port, SUMB_5_10_port, SUMB_5_9_port, SUMB_5_8_port, 
      SUMB_5_7_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_30_port, SUMB_4_29_port, 
      SUMB_4_28_port, SUMB_4_27_port, SUMB_4_26_port, SUMB_4_25_port, 
      SUMB_4_24_port, SUMB_4_23_port, SUMB_4_22_port, SUMB_4_21_port, 
      SUMB_4_20_port, SUMB_4_19_port, SUMB_4_18_port, SUMB_4_17_port, 
      SUMB_4_16_port, SUMB_4_15_port, SUMB_4_14_port, SUMB_4_13_port, 
      SUMB_4_12_port, SUMB_4_11_port, SUMB_4_10_port, SUMB_4_9_port, 
      SUMB_4_8_port, SUMB_4_7_port, SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port
      , SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_30_port, 
      SUMB_3_29_port, SUMB_3_28_port, SUMB_3_27_port, SUMB_3_26_port, 
      SUMB_3_25_port, SUMB_3_24_port, SUMB_3_23_port, SUMB_3_22_port, 
      SUMB_3_21_port, SUMB_3_20_port, SUMB_3_19_port, SUMB_3_18_port, 
      SUMB_3_17_port, SUMB_3_16_port, SUMB_3_15_port, SUMB_3_14_port, 
      SUMB_3_13_port, SUMB_3_12_port, SUMB_3_11_port, SUMB_3_10_port, 
      SUMB_3_9_port, SUMB_3_8_port, SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port
      , SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, SUMB_3_1_port, 
      SUMB_2_30_port, SUMB_2_29_port, SUMB_2_28_port, SUMB_2_27_port, 
      SUMB_2_26_port, SUMB_2_25_port, SUMB_2_24_port, SUMB_2_23_port, 
      SUMB_2_22_port, SUMB_2_21_port, SUMB_2_20_port, SUMB_2_19_port, 
      SUMB_2_18_port, SUMB_2_17_port, SUMB_2_16_port, SUMB_2_15_port, 
      SUMB_2_14_port, SUMB_2_13_port, SUMB_2_12_port, SUMB_2_11_port, 
      SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, SUMB_2_7_port, 
      SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port, SUMB_2_2_port
      , SUMB_2_1_port, CARRYB_31_30_port, CARRYB_31_29_port, CARRYB_31_28_port,
      CARRYB_31_27_port, CARRYB_31_26_port, CARRYB_31_25_port, 
      CARRYB_31_24_port, CARRYB_31_23_port, CARRYB_31_22_port, 
      CARRYB_31_21_port, CARRYB_31_20_port, CARRYB_31_19_port, 
      CARRYB_31_18_port, CARRYB_31_17_port, CARRYB_31_16_port, 
      CARRYB_31_15_port, CARRYB_31_14_port, CARRYB_31_13_port, 
      CARRYB_31_12_port, CARRYB_31_11_port, CARRYB_31_10_port, CARRYB_31_9_port
      , CARRYB_31_8_port, CARRYB_31_7_port, CARRYB_31_6_port, CARRYB_31_5_port,
      CARRYB_31_4_port, CARRYB_31_3_port, CARRYB_31_2_port, CARRYB_31_1_port, 
      CARRYB_31_0_port, CARRYB_30_30_port, CARRYB_30_29_port, CARRYB_30_28_port
      , CARRYB_30_27_port, CARRYB_30_26_port, CARRYB_30_25_port, 
      CARRYB_30_24_port, CARRYB_30_23_port, CARRYB_30_22_port, 
      CARRYB_30_21_port, CARRYB_30_20_port, CARRYB_30_19_port, 
      CARRYB_30_18_port, CARRYB_30_17_port, CARRYB_30_16_port, 
      CARRYB_30_15_port, CARRYB_30_14_port, CARRYB_30_13_port, 
      CARRYB_30_12_port, CARRYB_30_11_port, CARRYB_30_10_port, CARRYB_30_9_port
      , CARRYB_30_8_port, CARRYB_30_7_port, CARRYB_30_6_port, CARRYB_30_5_port,
      CARRYB_30_4_port, CARRYB_30_3_port, CARRYB_30_2_port, CARRYB_30_1_port, 
      CARRYB_30_0_port, CARRYB_29_30_port, CARRYB_29_29_port, CARRYB_29_28_port
      , CARRYB_29_27_port, CARRYB_29_26_port, CARRYB_29_25_port, 
      CARRYB_29_24_port, CARRYB_29_23_port, CARRYB_29_22_port, 
      CARRYB_29_21_port, CARRYB_29_20_port, CARRYB_29_19_port, 
      CARRYB_29_18_port, CARRYB_29_17_port, CARRYB_29_16_port, 
      CARRYB_29_15_port, CARRYB_29_14_port, CARRYB_29_13_port, 
      CARRYB_29_12_port, CARRYB_29_11_port, CARRYB_29_10_port, CARRYB_29_9_port
      , CARRYB_29_8_port, CARRYB_29_7_port, CARRYB_29_6_port, CARRYB_29_5_port,
      CARRYB_29_4_port, CARRYB_29_3_port, CARRYB_29_2_port, CARRYB_29_1_port, 
      CARRYB_29_0_port, CARRYB_28_30_port, CARRYB_28_29_port, CARRYB_28_28_port
      , CARRYB_28_27_port, CARRYB_28_26_port, CARRYB_28_25_port, 
      CARRYB_28_24_port, CARRYB_28_23_port, CARRYB_28_22_port, 
      CARRYB_28_21_port, CARRYB_28_20_port, CARRYB_28_19_port, 
      CARRYB_28_18_port, CARRYB_28_17_port, CARRYB_28_16_port, 
      CARRYB_28_15_port, CARRYB_28_14_port, CARRYB_28_13_port, 
      CARRYB_28_12_port, CARRYB_28_11_port, CARRYB_28_10_port, CARRYB_28_9_port
      , CARRYB_28_8_port, CARRYB_28_7_port, CARRYB_28_6_port, CARRYB_28_5_port,
      CARRYB_28_4_port, CARRYB_28_3_port, CARRYB_28_2_port, CARRYB_28_1_port, 
      CARRYB_28_0_port, CARRYB_27_30_port, CARRYB_27_29_port, CARRYB_27_28_port
      , CARRYB_27_27_port, CARRYB_27_26_port, CARRYB_27_25_port, 
      CARRYB_27_24_port, CARRYB_27_23_port, CARRYB_27_22_port, 
      CARRYB_27_21_port, CARRYB_27_20_port, CARRYB_27_19_port, 
      CARRYB_27_18_port, CARRYB_27_17_port, CARRYB_27_16_port, 
      CARRYB_27_15_port, CARRYB_27_14_port, CARRYB_27_13_port, 
      CARRYB_27_12_port, CARRYB_27_11_port, CARRYB_27_10_port, CARRYB_27_9_port
      , CARRYB_27_8_port, CARRYB_27_7_port, CARRYB_27_6_port, CARRYB_27_5_port,
      CARRYB_27_4_port, CARRYB_27_3_port, CARRYB_27_2_port, CARRYB_27_1_port, 
      CARRYB_27_0_port, CARRYB_26_30_port, CARRYB_26_29_port, CARRYB_26_28_port
      , CARRYB_26_27_port, CARRYB_26_26_port, CARRYB_26_25_port, 
      CARRYB_26_24_port, CARRYB_26_23_port, CARRYB_26_22_port, 
      CARRYB_26_21_port, CARRYB_26_20_port, CARRYB_26_19_port, 
      CARRYB_26_18_port, CARRYB_26_17_port, CARRYB_26_16_port, 
      CARRYB_26_15_port, CARRYB_26_14_port, CARRYB_26_13_port, 
      CARRYB_26_12_port, CARRYB_26_11_port, CARRYB_26_10_port, CARRYB_26_9_port
      , CARRYB_26_8_port, CARRYB_26_7_port, CARRYB_26_6_port, CARRYB_26_5_port,
      CARRYB_26_4_port, CARRYB_26_3_port, CARRYB_26_2_port, CARRYB_26_1_port, 
      CARRYB_26_0_port, CARRYB_25_30_port, CARRYB_25_29_port, CARRYB_25_28_port
      , CARRYB_25_27_port, CARRYB_25_26_port, CARRYB_25_25_port, 
      CARRYB_25_24_port, CARRYB_25_23_port, CARRYB_25_22_port, 
      CARRYB_25_21_port, CARRYB_25_20_port, CARRYB_25_19_port, 
      CARRYB_25_18_port, CARRYB_25_17_port, CARRYB_25_16_port, 
      CARRYB_25_15_port, CARRYB_25_14_port, CARRYB_25_13_port, 
      CARRYB_25_12_port, CARRYB_25_11_port, CARRYB_25_10_port, CARRYB_25_9_port
      , CARRYB_25_8_port, CARRYB_25_7_port, CARRYB_25_6_port, CARRYB_25_5_port,
      CARRYB_25_4_port, CARRYB_25_3_port, CARRYB_25_2_port, CARRYB_25_1_port, 
      CARRYB_25_0_port, CARRYB_24_30_port, CARRYB_24_29_port, CARRYB_24_28_port
      , CARRYB_24_27_port, CARRYB_24_26_port, CARRYB_24_25_port, 
      CARRYB_24_24_port, CARRYB_24_23_port, CARRYB_24_22_port, 
      CARRYB_24_21_port, CARRYB_24_20_port, CARRYB_24_19_port, 
      CARRYB_24_18_port, CARRYB_24_17_port, CARRYB_24_16_port, 
      CARRYB_24_15_port, CARRYB_24_14_port, CARRYB_24_13_port, 
      CARRYB_24_12_port, CARRYB_24_11_port, CARRYB_24_10_port, CARRYB_24_9_port
      , CARRYB_24_8_port, CARRYB_24_7_port, CARRYB_24_6_port, CARRYB_24_5_port,
      CARRYB_24_4_port, CARRYB_24_3_port, CARRYB_24_2_port, CARRYB_24_1_port, 
      CARRYB_24_0_port, CARRYB_23_30_port, CARRYB_23_29_port, CARRYB_23_28_port
      , CARRYB_23_27_port, CARRYB_23_26_port, CARRYB_23_25_port, 
      CARRYB_23_24_port, CARRYB_23_23_port, CARRYB_23_22_port, 
      CARRYB_23_21_port, CARRYB_23_20_port, CARRYB_23_19_port, 
      CARRYB_23_18_port, CARRYB_23_17_port, CARRYB_23_16_port, 
      CARRYB_23_15_port, CARRYB_23_14_port, CARRYB_23_13_port, 
      CARRYB_23_12_port, CARRYB_23_11_port, CARRYB_23_10_port, CARRYB_23_9_port
      , CARRYB_23_8_port, CARRYB_23_7_port, CARRYB_23_6_port, CARRYB_23_5_port,
      CARRYB_23_4_port, CARRYB_23_3_port, CARRYB_23_2_port, CARRYB_23_1_port, 
      CARRYB_23_0_port, CARRYB_22_30_port, CARRYB_22_29_port, CARRYB_22_28_port
      , CARRYB_22_27_port, CARRYB_22_26_port, CARRYB_22_25_port, 
      CARRYB_22_24_port, CARRYB_22_23_port, CARRYB_22_22_port, 
      CARRYB_22_21_port, CARRYB_22_20_port, CARRYB_22_19_port, 
      CARRYB_22_18_port, CARRYB_22_17_port, CARRYB_22_16_port, 
      CARRYB_22_15_port, CARRYB_22_14_port, CARRYB_22_13_port, 
      CARRYB_22_12_port, CARRYB_22_11_port, CARRYB_22_10_port, CARRYB_22_9_port
      , CARRYB_22_8_port, CARRYB_22_7_port, CARRYB_22_6_port, CARRYB_22_5_port,
      CARRYB_22_4_port, CARRYB_22_3_port, CARRYB_22_2_port, CARRYB_22_1_port, 
      CARRYB_22_0_port, CARRYB_21_30_port, CARRYB_21_29_port, CARRYB_21_28_port
      , CARRYB_21_27_port, CARRYB_21_26_port, CARRYB_21_25_port, 
      CARRYB_21_24_port, CARRYB_21_23_port, CARRYB_21_22_port, 
      CARRYB_21_21_port, CARRYB_21_20_port, CARRYB_21_19_port, 
      CARRYB_21_18_port, CARRYB_21_17_port, CARRYB_21_16_port, 
      CARRYB_21_15_port, CARRYB_21_14_port, CARRYB_21_13_port, 
      CARRYB_21_12_port, CARRYB_21_11_port, CARRYB_21_10_port, CARRYB_21_9_port
      , CARRYB_21_8_port, CARRYB_21_7_port, CARRYB_21_6_port, CARRYB_21_5_port,
      CARRYB_21_4_port, CARRYB_21_3_port, CARRYB_21_2_port, CARRYB_21_1_port, 
      CARRYB_21_0_port, CARRYB_20_30_port, CARRYB_20_29_port, CARRYB_20_28_port
      , CARRYB_20_27_port, CARRYB_20_26_port, CARRYB_20_25_port, 
      CARRYB_20_24_port, CARRYB_20_23_port, CARRYB_20_22_port, 
      CARRYB_20_21_port, CARRYB_20_20_port, CARRYB_20_19_port, 
      CARRYB_20_18_port, CARRYB_20_17_port, CARRYB_20_16_port, 
      CARRYB_20_15_port, CARRYB_20_14_port, CARRYB_20_13_port, 
      CARRYB_20_12_port, CARRYB_20_11_port, CARRYB_20_10_port, CARRYB_20_9_port
      , CARRYB_20_8_port, CARRYB_20_7_port, CARRYB_20_6_port, CARRYB_20_5_port,
      CARRYB_20_4_port, CARRYB_20_3_port, CARRYB_20_2_port, CARRYB_20_1_port, 
      CARRYB_20_0_port, CARRYB_19_30_port, CARRYB_19_29_port, CARRYB_19_28_port
      , CARRYB_19_27_port, CARRYB_19_26_port, CARRYB_19_25_port, 
      CARRYB_19_24_port, CARRYB_19_23_port, CARRYB_19_22_port, 
      CARRYB_19_21_port, CARRYB_19_20_port, CARRYB_19_19_port, 
      CARRYB_19_18_port, CARRYB_19_17_port, CARRYB_19_16_port, 
      CARRYB_19_15_port, CARRYB_19_14_port, CARRYB_19_13_port, 
      CARRYB_19_12_port, CARRYB_19_11_port, CARRYB_19_10_port, CARRYB_19_9_port
      , CARRYB_19_8_port, CARRYB_19_7_port, CARRYB_19_6_port, CARRYB_19_5_port,
      CARRYB_19_4_port, CARRYB_19_3_port, CARRYB_19_2_port, CARRYB_19_1_port, 
      CARRYB_19_0_port, CARRYB_18_30_port, CARRYB_18_29_port, CARRYB_18_28_port
      , CARRYB_18_27_port, CARRYB_18_26_port, CARRYB_18_25_port, 
      CARRYB_18_24_port, CARRYB_18_23_port, CARRYB_18_22_port, 
      CARRYB_18_21_port, CARRYB_18_20_port, CARRYB_18_19_port, 
      CARRYB_18_18_port, CARRYB_18_17_port, CARRYB_18_16_port, 
      CARRYB_18_15_port, CARRYB_18_14_port, CARRYB_18_13_port, 
      CARRYB_18_12_port, CARRYB_18_11_port, CARRYB_18_10_port, CARRYB_18_9_port
      , CARRYB_18_8_port, CARRYB_18_7_port, CARRYB_18_6_port, CARRYB_18_5_port,
      CARRYB_18_4_port, CARRYB_18_3_port, CARRYB_18_2_port, CARRYB_18_1_port, 
      CARRYB_18_0_port, CARRYB_17_30_port, CARRYB_17_29_port, CARRYB_17_28_port
      , CARRYB_17_27_port, CARRYB_17_26_port, CARRYB_17_25_port, 
      CARRYB_17_24_port, CARRYB_17_23_port, CARRYB_17_22_port, 
      CARRYB_17_21_port, CARRYB_17_20_port, CARRYB_17_19_port, 
      CARRYB_17_18_port, CARRYB_17_17_port, CARRYB_17_16_port, 
      CARRYB_17_15_port, CARRYB_17_14_port, CARRYB_17_13_port, 
      CARRYB_17_12_port, CARRYB_17_11_port, CARRYB_17_10_port, CARRYB_17_9_port
      , CARRYB_17_8_port, CARRYB_17_7_port, CARRYB_17_6_port, CARRYB_17_5_port,
      CARRYB_17_4_port, CARRYB_17_3_port, CARRYB_17_2_port, CARRYB_17_1_port, 
      CARRYB_17_0_port, CARRYB_16_30_port, CARRYB_16_29_port, CARRYB_16_28_port
      , CARRYB_16_27_port, CARRYB_16_26_port, CARRYB_16_25_port, 
      CARRYB_16_24_port, CARRYB_16_23_port, CARRYB_16_22_port, 
      CARRYB_16_21_port, CARRYB_16_20_port, CARRYB_16_19_port, 
      CARRYB_16_18_port, CARRYB_16_17_port, CARRYB_16_16_port, 
      CARRYB_16_15_port, CARRYB_16_14_port, CARRYB_16_13_port, 
      CARRYB_16_12_port, CARRYB_16_11_port, CARRYB_16_10_port, CARRYB_16_9_port
      , CARRYB_16_8_port, CARRYB_16_7_port, CARRYB_16_6_port, CARRYB_16_5_port,
      CARRYB_16_4_port, CARRYB_16_3_port, CARRYB_16_2_port, CARRYB_16_1_port, 
      CARRYB_16_0_port, SUMB_31_30_port, SUMB_31_29_port, SUMB_31_28_port, 
      SUMB_31_27_port, SUMB_31_26_port, SUMB_31_25_port, SUMB_31_24_port, 
      SUMB_31_23_port, SUMB_31_22_port, SUMB_31_21_port, SUMB_31_20_port, 
      SUMB_31_19_port, SUMB_31_18_port, SUMB_31_17_port, SUMB_31_16_port, 
      SUMB_31_15_port, SUMB_31_14_port, SUMB_31_13_port, SUMB_31_12_port, 
      SUMB_31_11_port, SUMB_31_10_port, SUMB_31_9_port, SUMB_31_8_port, 
      SUMB_31_7_port, SUMB_31_6_port, SUMB_31_5_port, SUMB_31_4_port, 
      SUMB_31_3_port, SUMB_31_2_port, SUMB_31_1_port, SUMB_31_0_port, 
      SUMB_30_30_port, SUMB_30_29_port, SUMB_30_28_port, SUMB_30_27_port, 
      SUMB_30_26_port, SUMB_30_25_port, SUMB_30_24_port, SUMB_30_23_port, 
      SUMB_30_22_port, SUMB_30_21_port, SUMB_30_20_port, SUMB_30_19_port, 
      SUMB_30_18_port, SUMB_30_17_port, SUMB_30_16_port, SUMB_30_15_port, 
      SUMB_30_14_port, SUMB_30_13_port, SUMB_30_12_port, SUMB_30_11_port, 
      SUMB_30_10_port, SUMB_30_9_port, SUMB_30_8_port, SUMB_30_7_port, 
      SUMB_30_6_port, SUMB_30_5_port, SUMB_30_4_port, SUMB_30_3_port, 
      SUMB_30_2_port, SUMB_30_1_port, SUMB_29_30_port, SUMB_29_29_port, 
      SUMB_29_28_port, SUMB_29_27_port, SUMB_29_26_port, SUMB_29_25_port, 
      SUMB_29_24_port, SUMB_29_23_port, SUMB_29_22_port, SUMB_29_21_port, 
      SUMB_29_20_port, SUMB_29_19_port, SUMB_29_18_port, SUMB_29_17_port, 
      SUMB_29_16_port, SUMB_29_15_port, SUMB_29_14_port, SUMB_29_13_port, 
      SUMB_29_12_port, SUMB_29_11_port, SUMB_29_10_port, SUMB_29_9_port, 
      SUMB_29_8_port, SUMB_29_7_port, SUMB_29_6_port, SUMB_29_5_port, 
      SUMB_29_4_port, SUMB_29_3_port, SUMB_29_2_port, SUMB_29_1_port, 
      SUMB_28_30_port, SUMB_28_29_port, SUMB_28_28_port, SUMB_28_27_port, 
      SUMB_28_26_port, SUMB_28_25_port, SUMB_28_24_port, SUMB_28_23_port, 
      SUMB_28_22_port, SUMB_28_21_port, SUMB_28_20_port, SUMB_28_19_port, 
      SUMB_28_18_port, SUMB_28_17_port, SUMB_28_16_port, SUMB_28_15_port, 
      SUMB_28_14_port, SUMB_28_13_port, SUMB_28_12_port, SUMB_28_11_port, 
      SUMB_28_10_port, SUMB_28_9_port, SUMB_28_8_port, SUMB_28_7_port, 
      SUMB_28_6_port, SUMB_28_5_port, SUMB_28_4_port, SUMB_28_3_port, 
      SUMB_28_2_port, SUMB_28_1_port, SUMB_27_30_port, SUMB_27_29_port, 
      SUMB_27_28_port, SUMB_27_27_port, SUMB_27_26_port, SUMB_27_25_port, 
      SUMB_27_24_port, SUMB_27_23_port, SUMB_27_22_port, SUMB_27_21_port, 
      SUMB_27_20_port, SUMB_27_19_port, SUMB_27_18_port, SUMB_27_17_port, 
      SUMB_27_16_port, SUMB_27_15_port, SUMB_27_14_port, SUMB_27_13_port, 
      SUMB_27_12_port, SUMB_27_11_port, SUMB_27_10_port, SUMB_27_9_port, 
      SUMB_27_8_port, SUMB_27_7_port, SUMB_27_6_port, SUMB_27_5_port, 
      SUMB_27_4_port, SUMB_27_3_port, SUMB_27_2_port, SUMB_27_1_port, 
      SUMB_26_30_port, SUMB_26_29_port, SUMB_26_28_port, SUMB_26_27_port, 
      SUMB_26_26_port, SUMB_26_25_port, SUMB_26_24_port, SUMB_26_23_port, 
      SUMB_26_22_port, SUMB_26_21_port, SUMB_26_20_port, SUMB_26_19_port, 
      SUMB_26_18_port, SUMB_26_17_port, SUMB_26_16_port, SUMB_26_15_port, 
      SUMB_26_14_port, SUMB_26_13_port, SUMB_26_12_port, SUMB_26_11_port, 
      SUMB_26_10_port, SUMB_26_9_port, SUMB_26_8_port, SUMB_26_7_port, 
      SUMB_26_6_port, SUMB_26_5_port, SUMB_26_4_port, SUMB_26_3_port, 
      SUMB_26_2_port, SUMB_26_1_port, SUMB_25_30_port, SUMB_25_29_port, 
      SUMB_25_28_port, SUMB_25_27_port, SUMB_25_26_port, SUMB_25_25_port, 
      SUMB_25_24_port, SUMB_25_23_port, SUMB_25_22_port, SUMB_25_21_port, 
      SUMB_25_20_port, SUMB_25_19_port, SUMB_25_18_port, SUMB_25_17_port, 
      SUMB_25_16_port, SUMB_25_15_port, SUMB_25_14_port, SUMB_25_13_port, 
      SUMB_25_12_port, SUMB_25_11_port, SUMB_25_10_port, SUMB_25_9_port, 
      SUMB_25_8_port, SUMB_25_7_port, SUMB_25_6_port, SUMB_25_5_port, 
      SUMB_25_4_port, SUMB_25_3_port, SUMB_25_2_port, SUMB_25_1_port, 
      SUMB_24_30_port, SUMB_24_29_port, SUMB_24_28_port, SUMB_24_27_port, 
      SUMB_24_26_port, SUMB_24_25_port, SUMB_24_24_port, SUMB_24_23_port, 
      SUMB_24_22_port, SUMB_24_21_port, SUMB_24_20_port, SUMB_24_19_port, 
      SUMB_24_18_port, SUMB_24_17_port, SUMB_24_16_port, SUMB_24_15_port, 
      SUMB_24_14_port, SUMB_24_13_port, SUMB_24_12_port, SUMB_24_11_port, 
      SUMB_24_10_port, SUMB_24_9_port, SUMB_24_8_port, SUMB_24_7_port, 
      SUMB_24_6_port, SUMB_24_5_port, SUMB_24_4_port, SUMB_24_3_port, 
      SUMB_24_2_port, SUMB_24_1_port, SUMB_23_30_port, SUMB_23_29_port, 
      SUMB_23_28_port, SUMB_23_27_port, SUMB_23_26_port, SUMB_23_25_port, 
      SUMB_23_24_port, SUMB_23_23_port, SUMB_23_22_port, SUMB_23_21_port, 
      SUMB_23_20_port, SUMB_23_19_port, SUMB_23_18_port, SUMB_23_17_port, 
      SUMB_23_16_port, SUMB_23_15_port, SUMB_23_14_port, SUMB_23_13_port, 
      SUMB_23_12_port, SUMB_23_11_port, SUMB_23_10_port, SUMB_23_9_port, 
      SUMB_23_8_port, SUMB_23_7_port, SUMB_23_6_port, SUMB_23_5_port, 
      SUMB_23_4_port, SUMB_23_3_port, SUMB_23_2_port, SUMB_23_1_port, 
      SUMB_22_30_port, SUMB_22_29_port, SUMB_22_28_port, SUMB_22_27_port, 
      SUMB_22_26_port, SUMB_22_25_port, SUMB_22_24_port, SUMB_22_23_port, 
      SUMB_22_22_port, SUMB_22_21_port, SUMB_22_20_port, SUMB_22_19_port, 
      SUMB_22_18_port, SUMB_22_17_port, SUMB_22_16_port, SUMB_22_15_port, 
      SUMB_22_14_port, SUMB_22_13_port, SUMB_22_12_port, SUMB_22_11_port, 
      SUMB_22_10_port, SUMB_22_9_port, SUMB_22_8_port, SUMB_22_7_port, 
      SUMB_22_6_port, SUMB_22_5_port, SUMB_22_4_port, SUMB_22_3_port, 
      SUMB_22_2_port, SUMB_22_1_port, SUMB_21_30_port, SUMB_21_29_port, 
      SUMB_21_28_port, SUMB_21_27_port, SUMB_21_26_port, SUMB_21_25_port, 
      SUMB_21_24_port, SUMB_21_23_port, SUMB_21_22_port, SUMB_21_21_port, 
      SUMB_21_20_port, SUMB_21_19_port, SUMB_21_18_port, SUMB_21_17_port, 
      SUMB_21_16_port, SUMB_21_15_port, SUMB_21_14_port, SUMB_21_13_port, 
      SUMB_21_12_port, SUMB_21_11_port, SUMB_21_10_port, SUMB_21_9_port, 
      SUMB_21_8_port, SUMB_21_7_port, SUMB_21_6_port, SUMB_21_5_port, 
      SUMB_21_4_port, SUMB_21_3_port, SUMB_21_2_port, SUMB_21_1_port, 
      SUMB_20_30_port, SUMB_20_29_port, SUMB_20_28_port, SUMB_20_27_port, 
      SUMB_20_26_port, SUMB_20_25_port, SUMB_20_24_port, SUMB_20_23_port, 
      SUMB_20_22_port, SUMB_20_21_port, SUMB_20_20_port, SUMB_20_19_port, 
      SUMB_20_18_port, SUMB_20_17_port, SUMB_20_16_port, SUMB_20_15_port, 
      SUMB_20_14_port, SUMB_20_13_port, SUMB_20_12_port, SUMB_20_11_port, 
      SUMB_20_10_port, SUMB_20_9_port, SUMB_20_8_port, SUMB_20_7_port, 
      SUMB_20_6_port, SUMB_20_5_port, SUMB_20_4_port, SUMB_20_3_port, 
      SUMB_20_2_port, SUMB_20_1_port, SUMB_19_30_port, SUMB_19_29_port, 
      SUMB_19_28_port, SUMB_19_27_port, SUMB_19_26_port, SUMB_19_25_port, 
      SUMB_19_24_port, SUMB_19_23_port, SUMB_19_22_port, SUMB_19_21_port, 
      SUMB_19_20_port, SUMB_19_19_port, SUMB_19_18_port, SUMB_19_17_port, 
      SUMB_19_16_port, SUMB_19_15_port, SUMB_19_14_port, SUMB_19_13_port, 
      SUMB_19_12_port, SUMB_19_11_port, SUMB_19_10_port, SUMB_19_9_port, 
      SUMB_19_8_port, SUMB_19_7_port, SUMB_19_6_port, SUMB_19_5_port, 
      SUMB_19_4_port, SUMB_19_3_port, SUMB_19_2_port, SUMB_19_1_port, 
      SUMB_18_30_port, SUMB_18_29_port, SUMB_18_28_port, SUMB_18_27_port, 
      SUMB_18_26_port, SUMB_18_25_port, SUMB_18_24_port, SUMB_18_23_port, 
      SUMB_18_22_port, SUMB_18_21_port, SUMB_18_20_port, SUMB_18_19_port, 
      SUMB_18_18_port, SUMB_18_17_port, SUMB_18_16_port, SUMB_18_15_port, 
      SUMB_18_14_port, SUMB_18_13_port, SUMB_18_12_port, SUMB_18_11_port, 
      SUMB_18_10_port, SUMB_18_9_port, SUMB_18_8_port, SUMB_18_7_port, 
      SUMB_18_6_port, SUMB_18_5_port, SUMB_18_4_port, SUMB_18_3_port, 
      SUMB_18_2_port, SUMB_18_1_port, SUMB_17_30_port, SUMB_17_29_port, 
      SUMB_17_28_port, SUMB_17_27_port, SUMB_17_26_port, SUMB_17_25_port, 
      SUMB_17_24_port, SUMB_17_23_port, SUMB_17_22_port, SUMB_17_21_port, 
      SUMB_17_20_port, SUMB_17_19_port, SUMB_17_18_port, SUMB_17_17_port, 
      SUMB_17_16_port, SUMB_17_15_port, SUMB_17_14_port, SUMB_17_13_port, 
      SUMB_17_12_port, SUMB_17_11_port, SUMB_17_10_port, SUMB_17_9_port, 
      SUMB_17_8_port, SUMB_17_7_port, SUMB_17_6_port, SUMB_17_5_port, 
      SUMB_17_4_port, SUMB_17_3_port, SUMB_17_2_port, SUMB_17_1_port, 
      SUMB_16_30_port, SUMB_16_29_port, SUMB_16_28_port, SUMB_16_27_port, 
      SUMB_16_26_port, SUMB_16_25_port, SUMB_16_24_port, SUMB_16_23_port, 
      SUMB_16_22_port, SUMB_16_21_port, SUMB_16_20_port, SUMB_16_19_port, 
      SUMB_16_18_port, SUMB_16_17_port, SUMB_16_16_port, SUMB_16_15_port, 
      SUMB_16_14_port, SUMB_16_13_port, SUMB_16_12_port, SUMB_16_11_port, 
      SUMB_16_10_port, SUMB_16_9_port, SUMB_16_8_port, SUMB_16_7_port, 
      SUMB_16_6_port, SUMB_16_5_port, SUMB_16_4_port, SUMB_16_3_port, 
      SUMB_16_2_port, SUMB_16_1_port, A1_28_port, A1_27_port, A1_26_port, 
      A1_25_port, A1_24_port, A1_23_port, A1_22_port, A1_21_port, A1_20_port, 
      A1_19_port, A1_18_port, A1_17_port, A1_16_port, A1_15_port, A1_14_port, 
      A1_13_port, A1_12_port, A1_11_port, A1_10_port, A1_9_port, A1_8_port, 
      A1_7_port, A1_6_port, A1_5_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n_1038 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_31_0_port, B => CARRYB_30_0_port, CI => 
                           SUMB_30_1_port, CO => CARRYB_31_0_port, S => 
                           SUMB_31_0_port);
   S4_1 : FA_X1 port map( A => ab_31_1_port, B => CARRYB_30_1_port, CI => 
                           SUMB_30_2_port, CO => CARRYB_31_1_port, S => 
                           SUMB_31_1_port);
   S4_2 : FA_X1 port map( A => ab_31_2_port, B => CARRYB_30_2_port, CI => 
                           SUMB_30_3_port, CO => CARRYB_31_2_port, S => 
                           SUMB_31_2_port);
   S4_3 : FA_X1 port map( A => ab_31_3_port, B => CARRYB_30_3_port, CI => 
                           SUMB_30_4_port, CO => CARRYB_31_3_port, S => 
                           SUMB_31_3_port);
   S4_4 : FA_X1 port map( A => ab_31_4_port, B => CARRYB_30_4_port, CI => 
                           SUMB_30_5_port, CO => CARRYB_31_4_port, S => 
                           SUMB_31_4_port);
   S4_5 : FA_X1 port map( A => ab_31_5_port, B => CARRYB_30_5_port, CI => 
                           SUMB_30_6_port, CO => CARRYB_31_5_port, S => 
                           SUMB_31_5_port);
   S4_6 : FA_X1 port map( A => ab_31_6_port, B => CARRYB_30_6_port, CI => 
                           SUMB_30_7_port, CO => CARRYB_31_6_port, S => 
                           SUMB_31_6_port);
   S4_7 : FA_X1 port map( A => ab_31_7_port, B => CARRYB_30_7_port, CI => 
                           SUMB_30_8_port, CO => CARRYB_31_7_port, S => 
                           SUMB_31_7_port);
   S4_8 : FA_X1 port map( A => ab_31_8_port, B => CARRYB_30_8_port, CI => 
                           SUMB_30_9_port, CO => CARRYB_31_8_port, S => 
                           SUMB_31_8_port);
   S4_9 : FA_X1 port map( A => ab_31_9_port, B => CARRYB_30_9_port, CI => 
                           SUMB_30_10_port, CO => CARRYB_31_9_port, S => 
                           SUMB_31_9_port);
   S4_10 : FA_X1 port map( A => ab_31_10_port, B => CARRYB_30_10_port, CI => 
                           SUMB_30_11_port, CO => CARRYB_31_10_port, S => 
                           SUMB_31_10_port);
   S4_11 : FA_X1 port map( A => ab_31_11_port, B => CARRYB_30_11_port, CI => 
                           SUMB_30_12_port, CO => CARRYB_31_11_port, S => 
                           SUMB_31_11_port);
   S4_12 : FA_X1 port map( A => ab_31_12_port, B => CARRYB_30_12_port, CI => 
                           SUMB_30_13_port, CO => CARRYB_31_12_port, S => 
                           SUMB_31_12_port);
   S4_13 : FA_X1 port map( A => ab_31_13_port, B => CARRYB_30_13_port, CI => 
                           SUMB_30_14_port, CO => CARRYB_31_13_port, S => 
                           SUMB_31_13_port);
   S4_14 : FA_X1 port map( A => ab_31_14_port, B => CARRYB_30_14_port, CI => 
                           SUMB_30_15_port, CO => CARRYB_31_14_port, S => 
                           SUMB_31_14_port);
   S4_15 : FA_X1 port map( A => ab_31_15_port, B => CARRYB_30_15_port, CI => 
                           SUMB_30_16_port, CO => CARRYB_31_15_port, S => 
                           SUMB_31_15_port);
   S4_16 : FA_X1 port map( A => ab_31_16_port, B => CARRYB_30_16_port, CI => 
                           SUMB_30_17_port, CO => CARRYB_31_16_port, S => 
                           SUMB_31_16_port);
   S4_17 : FA_X1 port map( A => ab_31_17_port, B => CARRYB_30_17_port, CI => 
                           SUMB_30_18_port, CO => CARRYB_31_17_port, S => 
                           SUMB_31_17_port);
   S4_18 : FA_X1 port map( A => ab_31_18_port, B => CARRYB_30_18_port, CI => 
                           SUMB_30_19_port, CO => CARRYB_31_18_port, S => 
                           SUMB_31_18_port);
   S4_19 : FA_X1 port map( A => ab_31_19_port, B => CARRYB_30_19_port, CI => 
                           SUMB_30_20_port, CO => CARRYB_31_19_port, S => 
                           SUMB_31_19_port);
   S4_20 : FA_X1 port map( A => ab_31_20_port, B => CARRYB_30_20_port, CI => 
                           SUMB_30_21_port, CO => CARRYB_31_20_port, S => 
                           SUMB_31_20_port);
   S4_21 : FA_X1 port map( A => ab_31_21_port, B => CARRYB_30_21_port, CI => 
                           SUMB_30_22_port, CO => CARRYB_31_21_port, S => 
                           SUMB_31_21_port);
   S4_22 : FA_X1 port map( A => ab_31_22_port, B => CARRYB_30_22_port, CI => 
                           SUMB_30_23_port, CO => CARRYB_31_22_port, S => 
                           SUMB_31_22_port);
   S4_23 : FA_X1 port map( A => ab_31_23_port, B => CARRYB_30_23_port, CI => 
                           SUMB_30_24_port, CO => CARRYB_31_23_port, S => 
                           SUMB_31_23_port);
   S4_24 : FA_X1 port map( A => ab_31_24_port, B => CARRYB_30_24_port, CI => 
                           SUMB_30_25_port, CO => CARRYB_31_24_port, S => 
                           SUMB_31_24_port);
   S4_25 : FA_X1 port map( A => ab_31_25_port, B => CARRYB_30_25_port, CI => 
                           SUMB_30_26_port, CO => CARRYB_31_25_port, S => 
                           SUMB_31_25_port);
   S4_26 : FA_X1 port map( A => ab_31_26_port, B => CARRYB_30_26_port, CI => 
                           SUMB_30_27_port, CO => CARRYB_31_26_port, S => 
                           SUMB_31_26_port);
   S4_27 : FA_X1 port map( A => ab_31_27_port, B => CARRYB_30_27_port, CI => 
                           SUMB_30_28_port, CO => CARRYB_31_27_port, S => 
                           SUMB_31_27_port);
   S4_28 : FA_X1 port map( A => ab_31_28_port, B => CARRYB_30_28_port, CI => 
                           SUMB_30_29_port, CO => CARRYB_31_28_port, S => 
                           SUMB_31_28_port);
   S4_29 : FA_X1 port map( A => ab_31_29_port, B => CARRYB_30_29_port, CI => 
                           SUMB_30_30_port, CO => CARRYB_31_29_port, S => 
                           SUMB_31_29_port);
   S5_30 : FA_X1 port map( A => ab_31_30_port, B => CARRYB_30_30_port, CI => 
                           ab_30_31_port, CO => CARRYB_31_30_port, S => 
                           SUMB_31_30_port);
   S1_30_0 : FA_X1 port map( A => ab_30_0_port, B => CARRYB_29_0_port, CI => 
                           SUMB_29_1_port, CO => CARRYB_30_0_port, S => 
                           A1_28_port);
   S2_30_1 : FA_X1 port map( A => ab_30_1_port, B => CARRYB_29_1_port, CI => 
                           SUMB_29_2_port, CO => CARRYB_30_1_port, S => 
                           SUMB_30_1_port);
   S2_30_2 : FA_X1 port map( A => ab_30_2_port, B => CARRYB_29_2_port, CI => 
                           SUMB_29_3_port, CO => CARRYB_30_2_port, S => 
                           SUMB_30_2_port);
   S2_30_3 : FA_X1 port map( A => ab_30_3_port, B => CARRYB_29_3_port, CI => 
                           SUMB_29_4_port, CO => CARRYB_30_3_port, S => 
                           SUMB_30_3_port);
   S2_30_4 : FA_X1 port map( A => ab_30_4_port, B => CARRYB_29_4_port, CI => 
                           SUMB_29_5_port, CO => CARRYB_30_4_port, S => 
                           SUMB_30_4_port);
   S2_30_5 : FA_X1 port map( A => ab_30_5_port, B => CARRYB_29_5_port, CI => 
                           SUMB_29_6_port, CO => CARRYB_30_5_port, S => 
                           SUMB_30_5_port);
   S2_30_6 : FA_X1 port map( A => ab_30_6_port, B => CARRYB_29_6_port, CI => 
                           SUMB_29_7_port, CO => CARRYB_30_6_port, S => 
                           SUMB_30_6_port);
   S2_30_7 : FA_X1 port map( A => ab_30_7_port, B => CARRYB_29_7_port, CI => 
                           SUMB_29_8_port, CO => CARRYB_30_7_port, S => 
                           SUMB_30_7_port);
   S2_30_8 : FA_X1 port map( A => ab_30_8_port, B => CARRYB_29_8_port, CI => 
                           SUMB_29_9_port, CO => CARRYB_30_8_port, S => 
                           SUMB_30_8_port);
   S2_30_9 : FA_X1 port map( A => ab_30_9_port, B => CARRYB_29_9_port, CI => 
                           SUMB_29_10_port, CO => CARRYB_30_9_port, S => 
                           SUMB_30_9_port);
   S2_30_10 : FA_X1 port map( A => ab_30_10_port, B => CARRYB_29_10_port, CI =>
                           SUMB_29_11_port, CO => CARRYB_30_10_port, S => 
                           SUMB_30_10_port);
   S2_30_11 : FA_X1 port map( A => ab_30_11_port, B => CARRYB_29_11_port, CI =>
                           SUMB_29_12_port, CO => CARRYB_30_11_port, S => 
                           SUMB_30_11_port);
   S2_30_12 : FA_X1 port map( A => ab_30_12_port, B => CARRYB_29_12_port, CI =>
                           SUMB_29_13_port, CO => CARRYB_30_12_port, S => 
                           SUMB_30_12_port);
   S2_30_13 : FA_X1 port map( A => ab_30_13_port, B => CARRYB_29_13_port, CI =>
                           SUMB_29_14_port, CO => CARRYB_30_13_port, S => 
                           SUMB_30_13_port);
   S2_30_14 : FA_X1 port map( A => ab_30_14_port, B => CARRYB_29_14_port, CI =>
                           SUMB_29_15_port, CO => CARRYB_30_14_port, S => 
                           SUMB_30_14_port);
   S2_30_15 : FA_X1 port map( A => ab_30_15_port, B => CARRYB_29_15_port, CI =>
                           SUMB_29_16_port, CO => CARRYB_30_15_port, S => 
                           SUMB_30_15_port);
   S2_30_16 : FA_X1 port map( A => ab_30_16_port, B => CARRYB_29_16_port, CI =>
                           SUMB_29_17_port, CO => CARRYB_30_16_port, S => 
                           SUMB_30_16_port);
   S2_30_17 : FA_X1 port map( A => ab_30_17_port, B => CARRYB_29_17_port, CI =>
                           SUMB_29_18_port, CO => CARRYB_30_17_port, S => 
                           SUMB_30_17_port);
   S2_30_18 : FA_X1 port map( A => ab_30_18_port, B => CARRYB_29_18_port, CI =>
                           SUMB_29_19_port, CO => CARRYB_30_18_port, S => 
                           SUMB_30_18_port);
   S2_30_19 : FA_X1 port map( A => ab_30_19_port, B => CARRYB_29_19_port, CI =>
                           SUMB_29_20_port, CO => CARRYB_30_19_port, S => 
                           SUMB_30_19_port);
   S2_30_20 : FA_X1 port map( A => ab_30_20_port, B => CARRYB_29_20_port, CI =>
                           SUMB_29_21_port, CO => CARRYB_30_20_port, S => 
                           SUMB_30_20_port);
   S2_30_21 : FA_X1 port map( A => ab_30_21_port, B => CARRYB_29_21_port, CI =>
                           SUMB_29_22_port, CO => CARRYB_30_21_port, S => 
                           SUMB_30_21_port);
   S2_30_22 : FA_X1 port map( A => ab_30_22_port, B => CARRYB_29_22_port, CI =>
                           SUMB_29_23_port, CO => CARRYB_30_22_port, S => 
                           SUMB_30_22_port);
   S2_30_23 : FA_X1 port map( A => ab_30_23_port, B => CARRYB_29_23_port, CI =>
                           SUMB_29_24_port, CO => CARRYB_30_23_port, S => 
                           SUMB_30_23_port);
   S2_30_24 : FA_X1 port map( A => ab_30_24_port, B => CARRYB_29_24_port, CI =>
                           SUMB_29_25_port, CO => CARRYB_30_24_port, S => 
                           SUMB_30_24_port);
   S2_30_25 : FA_X1 port map( A => ab_30_25_port, B => CARRYB_29_25_port, CI =>
                           SUMB_29_26_port, CO => CARRYB_30_25_port, S => 
                           SUMB_30_25_port);
   S2_30_26 : FA_X1 port map( A => ab_30_26_port, B => CARRYB_29_26_port, CI =>
                           SUMB_29_27_port, CO => CARRYB_30_26_port, S => 
                           SUMB_30_26_port);
   S2_30_27 : FA_X1 port map( A => ab_30_27_port, B => CARRYB_29_27_port, CI =>
                           SUMB_29_28_port, CO => CARRYB_30_27_port, S => 
                           SUMB_30_27_port);
   S2_30_28 : FA_X1 port map( A => ab_30_28_port, B => CARRYB_29_28_port, CI =>
                           SUMB_29_29_port, CO => CARRYB_30_28_port, S => 
                           SUMB_30_28_port);
   S2_30_29 : FA_X1 port map( A => ab_30_29_port, B => CARRYB_29_29_port, CI =>
                           SUMB_29_30_port, CO => CARRYB_30_29_port, S => 
                           SUMB_30_29_port);
   S3_30_30 : FA_X1 port map( A => ab_30_30_port, B => CARRYB_29_30_port, CI =>
                           ab_29_31_port, CO => CARRYB_30_30_port, S => 
                           SUMB_30_30_port);
   S1_29_0 : FA_X1 port map( A => ab_29_0_port, B => CARRYB_28_0_port, CI => 
                           SUMB_28_1_port, CO => CARRYB_29_0_port, S => 
                           A1_27_port);
   S2_29_1 : FA_X1 port map( A => ab_29_1_port, B => CARRYB_28_1_port, CI => 
                           SUMB_28_2_port, CO => CARRYB_29_1_port, S => 
                           SUMB_29_1_port);
   S2_29_2 : FA_X1 port map( A => ab_29_2_port, B => CARRYB_28_2_port, CI => 
                           SUMB_28_3_port, CO => CARRYB_29_2_port, S => 
                           SUMB_29_2_port);
   S2_29_3 : FA_X1 port map( A => ab_29_3_port, B => CARRYB_28_3_port, CI => 
                           SUMB_28_4_port, CO => CARRYB_29_3_port, S => 
                           SUMB_29_3_port);
   S2_29_4 : FA_X1 port map( A => ab_29_4_port, B => CARRYB_28_4_port, CI => 
                           SUMB_28_5_port, CO => CARRYB_29_4_port, S => 
                           SUMB_29_4_port);
   S2_29_5 : FA_X1 port map( A => ab_29_5_port, B => CARRYB_28_5_port, CI => 
                           SUMB_28_6_port, CO => CARRYB_29_5_port, S => 
                           SUMB_29_5_port);
   S2_29_6 : FA_X1 port map( A => ab_29_6_port, B => CARRYB_28_6_port, CI => 
                           SUMB_28_7_port, CO => CARRYB_29_6_port, S => 
                           SUMB_29_6_port);
   S2_29_7 : FA_X1 port map( A => ab_29_7_port, B => CARRYB_28_7_port, CI => 
                           SUMB_28_8_port, CO => CARRYB_29_7_port, S => 
                           SUMB_29_7_port);
   S2_29_8 : FA_X1 port map( A => ab_29_8_port, B => CARRYB_28_8_port, CI => 
                           SUMB_28_9_port, CO => CARRYB_29_8_port, S => 
                           SUMB_29_8_port);
   S2_29_9 : FA_X1 port map( A => ab_29_9_port, B => CARRYB_28_9_port, CI => 
                           SUMB_28_10_port, CO => CARRYB_29_9_port, S => 
                           SUMB_29_9_port);
   S2_29_10 : FA_X1 port map( A => ab_29_10_port, B => CARRYB_28_10_port, CI =>
                           SUMB_28_11_port, CO => CARRYB_29_10_port, S => 
                           SUMB_29_10_port);
   S2_29_11 : FA_X1 port map( A => ab_29_11_port, B => CARRYB_28_11_port, CI =>
                           SUMB_28_12_port, CO => CARRYB_29_11_port, S => 
                           SUMB_29_11_port);
   S2_29_12 : FA_X1 port map( A => ab_29_12_port, B => CARRYB_28_12_port, CI =>
                           SUMB_28_13_port, CO => CARRYB_29_12_port, S => 
                           SUMB_29_12_port);
   S2_29_13 : FA_X1 port map( A => ab_29_13_port, B => CARRYB_28_13_port, CI =>
                           SUMB_28_14_port, CO => CARRYB_29_13_port, S => 
                           SUMB_29_13_port);
   S2_29_14 : FA_X1 port map( A => ab_29_14_port, B => CARRYB_28_14_port, CI =>
                           SUMB_28_15_port, CO => CARRYB_29_14_port, S => 
                           SUMB_29_14_port);
   S2_29_15 : FA_X1 port map( A => ab_29_15_port, B => CARRYB_28_15_port, CI =>
                           SUMB_28_16_port, CO => CARRYB_29_15_port, S => 
                           SUMB_29_15_port);
   S2_29_16 : FA_X1 port map( A => ab_29_16_port, B => CARRYB_28_16_port, CI =>
                           SUMB_28_17_port, CO => CARRYB_29_16_port, S => 
                           SUMB_29_16_port);
   S2_29_17 : FA_X1 port map( A => ab_29_17_port, B => CARRYB_28_17_port, CI =>
                           SUMB_28_18_port, CO => CARRYB_29_17_port, S => 
                           SUMB_29_17_port);
   S2_29_18 : FA_X1 port map( A => ab_29_18_port, B => CARRYB_28_18_port, CI =>
                           SUMB_28_19_port, CO => CARRYB_29_18_port, S => 
                           SUMB_29_18_port);
   S2_29_19 : FA_X1 port map( A => ab_29_19_port, B => CARRYB_28_19_port, CI =>
                           SUMB_28_20_port, CO => CARRYB_29_19_port, S => 
                           SUMB_29_19_port);
   S2_29_20 : FA_X1 port map( A => ab_29_20_port, B => CARRYB_28_20_port, CI =>
                           SUMB_28_21_port, CO => CARRYB_29_20_port, S => 
                           SUMB_29_20_port);
   S2_29_21 : FA_X1 port map( A => ab_29_21_port, B => CARRYB_28_21_port, CI =>
                           SUMB_28_22_port, CO => CARRYB_29_21_port, S => 
                           SUMB_29_21_port);
   S2_29_22 : FA_X1 port map( A => ab_29_22_port, B => CARRYB_28_22_port, CI =>
                           SUMB_28_23_port, CO => CARRYB_29_22_port, S => 
                           SUMB_29_22_port);
   S2_29_23 : FA_X1 port map( A => ab_29_23_port, B => CARRYB_28_23_port, CI =>
                           SUMB_28_24_port, CO => CARRYB_29_23_port, S => 
                           SUMB_29_23_port);
   S2_29_24 : FA_X1 port map( A => ab_29_24_port, B => CARRYB_28_24_port, CI =>
                           SUMB_28_25_port, CO => CARRYB_29_24_port, S => 
                           SUMB_29_24_port);
   S2_29_25 : FA_X1 port map( A => ab_29_25_port, B => CARRYB_28_25_port, CI =>
                           SUMB_28_26_port, CO => CARRYB_29_25_port, S => 
                           SUMB_29_25_port);
   S2_29_26 : FA_X1 port map( A => ab_29_26_port, B => CARRYB_28_26_port, CI =>
                           SUMB_28_27_port, CO => CARRYB_29_26_port, S => 
                           SUMB_29_26_port);
   S2_29_27 : FA_X1 port map( A => ab_29_27_port, B => CARRYB_28_27_port, CI =>
                           SUMB_28_28_port, CO => CARRYB_29_27_port, S => 
                           SUMB_29_27_port);
   S2_29_28 : FA_X1 port map( A => ab_29_28_port, B => CARRYB_28_28_port, CI =>
                           SUMB_28_29_port, CO => CARRYB_29_28_port, S => 
                           SUMB_29_28_port);
   S2_29_29 : FA_X1 port map( A => ab_29_29_port, B => CARRYB_28_29_port, CI =>
                           SUMB_28_30_port, CO => CARRYB_29_29_port, S => 
                           SUMB_29_29_port);
   S3_29_30 : FA_X1 port map( A => ab_29_30_port, B => CARRYB_28_30_port, CI =>
                           ab_28_31_port, CO => CARRYB_29_30_port, S => 
                           SUMB_29_30_port);
   S1_28_0 : FA_X1 port map( A => ab_28_0_port, B => CARRYB_27_0_port, CI => 
                           SUMB_27_1_port, CO => CARRYB_28_0_port, S => 
                           A1_26_port);
   S2_28_1 : FA_X1 port map( A => ab_28_1_port, B => CARRYB_27_1_port, CI => 
                           SUMB_27_2_port, CO => CARRYB_28_1_port, S => 
                           SUMB_28_1_port);
   S2_28_2 : FA_X1 port map( A => ab_28_2_port, B => CARRYB_27_2_port, CI => 
                           SUMB_27_3_port, CO => CARRYB_28_2_port, S => 
                           SUMB_28_2_port);
   S2_28_3 : FA_X1 port map( A => ab_28_3_port, B => CARRYB_27_3_port, CI => 
                           SUMB_27_4_port, CO => CARRYB_28_3_port, S => 
                           SUMB_28_3_port);
   S2_28_4 : FA_X1 port map( A => ab_28_4_port, B => CARRYB_27_4_port, CI => 
                           SUMB_27_5_port, CO => CARRYB_28_4_port, S => 
                           SUMB_28_4_port);
   S2_28_5 : FA_X1 port map( A => ab_28_5_port, B => CARRYB_27_5_port, CI => 
                           SUMB_27_6_port, CO => CARRYB_28_5_port, S => 
                           SUMB_28_5_port);
   S2_28_6 : FA_X1 port map( A => ab_28_6_port, B => CARRYB_27_6_port, CI => 
                           SUMB_27_7_port, CO => CARRYB_28_6_port, S => 
                           SUMB_28_6_port);
   S2_28_7 : FA_X1 port map( A => ab_28_7_port, B => CARRYB_27_7_port, CI => 
                           SUMB_27_8_port, CO => CARRYB_28_7_port, S => 
                           SUMB_28_7_port);
   S2_28_8 : FA_X1 port map( A => ab_28_8_port, B => CARRYB_27_8_port, CI => 
                           SUMB_27_9_port, CO => CARRYB_28_8_port, S => 
                           SUMB_28_8_port);
   S2_28_9 : FA_X1 port map( A => ab_28_9_port, B => CARRYB_27_9_port, CI => 
                           SUMB_27_10_port, CO => CARRYB_28_9_port, S => 
                           SUMB_28_9_port);
   S2_28_10 : FA_X1 port map( A => ab_28_10_port, B => CARRYB_27_10_port, CI =>
                           SUMB_27_11_port, CO => CARRYB_28_10_port, S => 
                           SUMB_28_10_port);
   S2_28_11 : FA_X1 port map( A => ab_28_11_port, B => CARRYB_27_11_port, CI =>
                           SUMB_27_12_port, CO => CARRYB_28_11_port, S => 
                           SUMB_28_11_port);
   S2_28_12 : FA_X1 port map( A => ab_28_12_port, B => CARRYB_27_12_port, CI =>
                           SUMB_27_13_port, CO => CARRYB_28_12_port, S => 
                           SUMB_28_12_port);
   S2_28_13 : FA_X1 port map( A => ab_28_13_port, B => CARRYB_27_13_port, CI =>
                           SUMB_27_14_port, CO => CARRYB_28_13_port, S => 
                           SUMB_28_13_port);
   S2_28_14 : FA_X1 port map( A => ab_28_14_port, B => CARRYB_27_14_port, CI =>
                           SUMB_27_15_port, CO => CARRYB_28_14_port, S => 
                           SUMB_28_14_port);
   S2_28_15 : FA_X1 port map( A => ab_28_15_port, B => CARRYB_27_15_port, CI =>
                           SUMB_27_16_port, CO => CARRYB_28_15_port, S => 
                           SUMB_28_15_port);
   S2_28_16 : FA_X1 port map( A => ab_28_16_port, B => CARRYB_27_16_port, CI =>
                           SUMB_27_17_port, CO => CARRYB_28_16_port, S => 
                           SUMB_28_16_port);
   S2_28_17 : FA_X1 port map( A => ab_28_17_port, B => CARRYB_27_17_port, CI =>
                           SUMB_27_18_port, CO => CARRYB_28_17_port, S => 
                           SUMB_28_17_port);
   S2_28_18 : FA_X1 port map( A => ab_28_18_port, B => CARRYB_27_18_port, CI =>
                           SUMB_27_19_port, CO => CARRYB_28_18_port, S => 
                           SUMB_28_18_port);
   S2_28_19 : FA_X1 port map( A => ab_28_19_port, B => CARRYB_27_19_port, CI =>
                           SUMB_27_20_port, CO => CARRYB_28_19_port, S => 
                           SUMB_28_19_port);
   S2_28_20 : FA_X1 port map( A => ab_28_20_port, B => CARRYB_27_20_port, CI =>
                           SUMB_27_21_port, CO => CARRYB_28_20_port, S => 
                           SUMB_28_20_port);
   S2_28_21 : FA_X1 port map( A => ab_28_21_port, B => CARRYB_27_21_port, CI =>
                           SUMB_27_22_port, CO => CARRYB_28_21_port, S => 
                           SUMB_28_21_port);
   S2_28_22 : FA_X1 port map( A => ab_28_22_port, B => CARRYB_27_22_port, CI =>
                           SUMB_27_23_port, CO => CARRYB_28_22_port, S => 
                           SUMB_28_22_port);
   S2_28_23 : FA_X1 port map( A => ab_28_23_port, B => CARRYB_27_23_port, CI =>
                           SUMB_27_24_port, CO => CARRYB_28_23_port, S => 
                           SUMB_28_23_port);
   S2_28_24 : FA_X1 port map( A => ab_28_24_port, B => CARRYB_27_24_port, CI =>
                           SUMB_27_25_port, CO => CARRYB_28_24_port, S => 
                           SUMB_28_24_port);
   S2_28_25 : FA_X1 port map( A => ab_28_25_port, B => CARRYB_27_25_port, CI =>
                           SUMB_27_26_port, CO => CARRYB_28_25_port, S => 
                           SUMB_28_25_port);
   S2_28_26 : FA_X1 port map( A => ab_28_26_port, B => CARRYB_27_26_port, CI =>
                           SUMB_27_27_port, CO => CARRYB_28_26_port, S => 
                           SUMB_28_26_port);
   S2_28_27 : FA_X1 port map( A => ab_28_27_port, B => CARRYB_27_27_port, CI =>
                           SUMB_27_28_port, CO => CARRYB_28_27_port, S => 
                           SUMB_28_27_port);
   S2_28_28 : FA_X1 port map( A => ab_28_28_port, B => CARRYB_27_28_port, CI =>
                           SUMB_27_29_port, CO => CARRYB_28_28_port, S => 
                           SUMB_28_28_port);
   S2_28_29 : FA_X1 port map( A => ab_28_29_port, B => CARRYB_27_29_port, CI =>
                           SUMB_27_30_port, CO => CARRYB_28_29_port, S => 
                           SUMB_28_29_port);
   S3_28_30 : FA_X1 port map( A => ab_28_30_port, B => CARRYB_27_30_port, CI =>
                           ab_27_31_port, CO => CARRYB_28_30_port, S => 
                           SUMB_28_30_port);
   S1_27_0 : FA_X1 port map( A => ab_27_0_port, B => CARRYB_26_0_port, CI => 
                           SUMB_26_1_port, CO => CARRYB_27_0_port, S => 
                           A1_25_port);
   S2_27_1 : FA_X1 port map( A => ab_27_1_port, B => CARRYB_26_1_port, CI => 
                           SUMB_26_2_port, CO => CARRYB_27_1_port, S => 
                           SUMB_27_1_port);
   S2_27_2 : FA_X1 port map( A => ab_27_2_port, B => CARRYB_26_2_port, CI => 
                           SUMB_26_3_port, CO => CARRYB_27_2_port, S => 
                           SUMB_27_2_port);
   S2_27_3 : FA_X1 port map( A => ab_27_3_port, B => CARRYB_26_3_port, CI => 
                           SUMB_26_4_port, CO => CARRYB_27_3_port, S => 
                           SUMB_27_3_port);
   S2_27_4 : FA_X1 port map( A => ab_27_4_port, B => CARRYB_26_4_port, CI => 
                           SUMB_26_5_port, CO => CARRYB_27_4_port, S => 
                           SUMB_27_4_port);
   S2_27_5 : FA_X1 port map( A => ab_27_5_port, B => CARRYB_26_5_port, CI => 
                           SUMB_26_6_port, CO => CARRYB_27_5_port, S => 
                           SUMB_27_5_port);
   S2_27_6 : FA_X1 port map( A => ab_27_6_port, B => CARRYB_26_6_port, CI => 
                           SUMB_26_7_port, CO => CARRYB_27_6_port, S => 
                           SUMB_27_6_port);
   S2_27_7 : FA_X1 port map( A => ab_27_7_port, B => CARRYB_26_7_port, CI => 
                           SUMB_26_8_port, CO => CARRYB_27_7_port, S => 
                           SUMB_27_7_port);
   S2_27_8 : FA_X1 port map( A => ab_27_8_port, B => CARRYB_26_8_port, CI => 
                           SUMB_26_9_port, CO => CARRYB_27_8_port, S => 
                           SUMB_27_8_port);
   S2_27_9 : FA_X1 port map( A => ab_27_9_port, B => CARRYB_26_9_port, CI => 
                           SUMB_26_10_port, CO => CARRYB_27_9_port, S => 
                           SUMB_27_9_port);
   S2_27_10 : FA_X1 port map( A => ab_27_10_port, B => CARRYB_26_10_port, CI =>
                           SUMB_26_11_port, CO => CARRYB_27_10_port, S => 
                           SUMB_27_10_port);
   S2_27_11 : FA_X1 port map( A => ab_27_11_port, B => CARRYB_26_11_port, CI =>
                           SUMB_26_12_port, CO => CARRYB_27_11_port, S => 
                           SUMB_27_11_port);
   S2_27_12 : FA_X1 port map( A => ab_27_12_port, B => CARRYB_26_12_port, CI =>
                           SUMB_26_13_port, CO => CARRYB_27_12_port, S => 
                           SUMB_27_12_port);
   S2_27_13 : FA_X1 port map( A => ab_27_13_port, B => CARRYB_26_13_port, CI =>
                           SUMB_26_14_port, CO => CARRYB_27_13_port, S => 
                           SUMB_27_13_port);
   S2_27_14 : FA_X1 port map( A => ab_27_14_port, B => CARRYB_26_14_port, CI =>
                           SUMB_26_15_port, CO => CARRYB_27_14_port, S => 
                           SUMB_27_14_port);
   S2_27_15 : FA_X1 port map( A => ab_27_15_port, B => CARRYB_26_15_port, CI =>
                           SUMB_26_16_port, CO => CARRYB_27_15_port, S => 
                           SUMB_27_15_port);
   S2_27_16 : FA_X1 port map( A => ab_27_16_port, B => CARRYB_26_16_port, CI =>
                           SUMB_26_17_port, CO => CARRYB_27_16_port, S => 
                           SUMB_27_16_port);
   S2_27_17 : FA_X1 port map( A => ab_27_17_port, B => CARRYB_26_17_port, CI =>
                           SUMB_26_18_port, CO => CARRYB_27_17_port, S => 
                           SUMB_27_17_port);
   S2_27_18 : FA_X1 port map( A => ab_27_18_port, B => CARRYB_26_18_port, CI =>
                           SUMB_26_19_port, CO => CARRYB_27_18_port, S => 
                           SUMB_27_18_port);
   S2_27_19 : FA_X1 port map( A => ab_27_19_port, B => CARRYB_26_19_port, CI =>
                           SUMB_26_20_port, CO => CARRYB_27_19_port, S => 
                           SUMB_27_19_port);
   S2_27_20 : FA_X1 port map( A => ab_27_20_port, B => CARRYB_26_20_port, CI =>
                           SUMB_26_21_port, CO => CARRYB_27_20_port, S => 
                           SUMB_27_20_port);
   S2_27_21 : FA_X1 port map( A => ab_27_21_port, B => CARRYB_26_21_port, CI =>
                           SUMB_26_22_port, CO => CARRYB_27_21_port, S => 
                           SUMB_27_21_port);
   S2_27_22 : FA_X1 port map( A => ab_27_22_port, B => CARRYB_26_22_port, CI =>
                           SUMB_26_23_port, CO => CARRYB_27_22_port, S => 
                           SUMB_27_22_port);
   S2_27_23 : FA_X1 port map( A => ab_27_23_port, B => CARRYB_26_23_port, CI =>
                           SUMB_26_24_port, CO => CARRYB_27_23_port, S => 
                           SUMB_27_23_port);
   S2_27_24 : FA_X1 port map( A => ab_27_24_port, B => CARRYB_26_24_port, CI =>
                           SUMB_26_25_port, CO => CARRYB_27_24_port, S => 
                           SUMB_27_24_port);
   S2_27_25 : FA_X1 port map( A => ab_27_25_port, B => CARRYB_26_25_port, CI =>
                           SUMB_26_26_port, CO => CARRYB_27_25_port, S => 
                           SUMB_27_25_port);
   S2_27_26 : FA_X1 port map( A => ab_27_26_port, B => CARRYB_26_26_port, CI =>
                           SUMB_26_27_port, CO => CARRYB_27_26_port, S => 
                           SUMB_27_26_port);
   S2_27_27 : FA_X1 port map( A => ab_27_27_port, B => CARRYB_26_27_port, CI =>
                           SUMB_26_28_port, CO => CARRYB_27_27_port, S => 
                           SUMB_27_27_port);
   S2_27_28 : FA_X1 port map( A => ab_27_28_port, B => CARRYB_26_28_port, CI =>
                           SUMB_26_29_port, CO => CARRYB_27_28_port, S => 
                           SUMB_27_28_port);
   S2_27_29 : FA_X1 port map( A => ab_27_29_port, B => CARRYB_26_29_port, CI =>
                           SUMB_26_30_port, CO => CARRYB_27_29_port, S => 
                           SUMB_27_29_port);
   S3_27_30 : FA_X1 port map( A => ab_27_30_port, B => CARRYB_26_30_port, CI =>
                           ab_26_31_port, CO => CARRYB_27_30_port, S => 
                           SUMB_27_30_port);
   S1_26_0 : FA_X1 port map( A => ab_26_0_port, B => CARRYB_25_0_port, CI => 
                           SUMB_25_1_port, CO => CARRYB_26_0_port, S => 
                           A1_24_port);
   S2_26_1 : FA_X1 port map( A => ab_26_1_port, B => CARRYB_25_1_port, CI => 
                           SUMB_25_2_port, CO => CARRYB_26_1_port, S => 
                           SUMB_26_1_port);
   S2_26_2 : FA_X1 port map( A => ab_26_2_port, B => CARRYB_25_2_port, CI => 
                           SUMB_25_3_port, CO => CARRYB_26_2_port, S => 
                           SUMB_26_2_port);
   S2_26_3 : FA_X1 port map( A => ab_26_3_port, B => CARRYB_25_3_port, CI => 
                           SUMB_25_4_port, CO => CARRYB_26_3_port, S => 
                           SUMB_26_3_port);
   S2_26_4 : FA_X1 port map( A => ab_26_4_port, B => CARRYB_25_4_port, CI => 
                           SUMB_25_5_port, CO => CARRYB_26_4_port, S => 
                           SUMB_26_4_port);
   S2_26_5 : FA_X1 port map( A => ab_26_5_port, B => CARRYB_25_5_port, CI => 
                           SUMB_25_6_port, CO => CARRYB_26_5_port, S => 
                           SUMB_26_5_port);
   S2_26_6 : FA_X1 port map( A => ab_26_6_port, B => CARRYB_25_6_port, CI => 
                           SUMB_25_7_port, CO => CARRYB_26_6_port, S => 
                           SUMB_26_6_port);
   S2_26_7 : FA_X1 port map( A => ab_26_7_port, B => CARRYB_25_7_port, CI => 
                           SUMB_25_8_port, CO => CARRYB_26_7_port, S => 
                           SUMB_26_7_port);
   S2_26_8 : FA_X1 port map( A => ab_26_8_port, B => CARRYB_25_8_port, CI => 
                           SUMB_25_9_port, CO => CARRYB_26_8_port, S => 
                           SUMB_26_8_port);
   S2_26_9 : FA_X1 port map( A => ab_26_9_port, B => CARRYB_25_9_port, CI => 
                           SUMB_25_10_port, CO => CARRYB_26_9_port, S => 
                           SUMB_26_9_port);
   S2_26_10 : FA_X1 port map( A => ab_26_10_port, B => CARRYB_25_10_port, CI =>
                           SUMB_25_11_port, CO => CARRYB_26_10_port, S => 
                           SUMB_26_10_port);
   S2_26_11 : FA_X1 port map( A => ab_26_11_port, B => CARRYB_25_11_port, CI =>
                           SUMB_25_12_port, CO => CARRYB_26_11_port, S => 
                           SUMB_26_11_port);
   S2_26_12 : FA_X1 port map( A => ab_26_12_port, B => CARRYB_25_12_port, CI =>
                           SUMB_25_13_port, CO => CARRYB_26_12_port, S => 
                           SUMB_26_12_port);
   S2_26_13 : FA_X1 port map( A => ab_26_13_port, B => CARRYB_25_13_port, CI =>
                           SUMB_25_14_port, CO => CARRYB_26_13_port, S => 
                           SUMB_26_13_port);
   S2_26_14 : FA_X1 port map( A => ab_26_14_port, B => CARRYB_25_14_port, CI =>
                           SUMB_25_15_port, CO => CARRYB_26_14_port, S => 
                           SUMB_26_14_port);
   S2_26_15 : FA_X1 port map( A => ab_26_15_port, B => CARRYB_25_15_port, CI =>
                           SUMB_25_16_port, CO => CARRYB_26_15_port, S => 
                           SUMB_26_15_port);
   S2_26_16 : FA_X1 port map( A => ab_26_16_port, B => CARRYB_25_16_port, CI =>
                           SUMB_25_17_port, CO => CARRYB_26_16_port, S => 
                           SUMB_26_16_port);
   S2_26_17 : FA_X1 port map( A => ab_26_17_port, B => CARRYB_25_17_port, CI =>
                           SUMB_25_18_port, CO => CARRYB_26_17_port, S => 
                           SUMB_26_17_port);
   S2_26_18 : FA_X1 port map( A => ab_26_18_port, B => CARRYB_25_18_port, CI =>
                           SUMB_25_19_port, CO => CARRYB_26_18_port, S => 
                           SUMB_26_18_port);
   S2_26_19 : FA_X1 port map( A => ab_26_19_port, B => CARRYB_25_19_port, CI =>
                           SUMB_25_20_port, CO => CARRYB_26_19_port, S => 
                           SUMB_26_19_port);
   S2_26_20 : FA_X1 port map( A => ab_26_20_port, B => CARRYB_25_20_port, CI =>
                           SUMB_25_21_port, CO => CARRYB_26_20_port, S => 
                           SUMB_26_20_port);
   S2_26_21 : FA_X1 port map( A => ab_26_21_port, B => CARRYB_25_21_port, CI =>
                           SUMB_25_22_port, CO => CARRYB_26_21_port, S => 
                           SUMB_26_21_port);
   S2_26_22 : FA_X1 port map( A => ab_26_22_port, B => CARRYB_25_22_port, CI =>
                           SUMB_25_23_port, CO => CARRYB_26_22_port, S => 
                           SUMB_26_22_port);
   S2_26_23 : FA_X1 port map( A => ab_26_23_port, B => CARRYB_25_23_port, CI =>
                           SUMB_25_24_port, CO => CARRYB_26_23_port, S => 
                           SUMB_26_23_port);
   S2_26_24 : FA_X1 port map( A => ab_26_24_port, B => CARRYB_25_24_port, CI =>
                           SUMB_25_25_port, CO => CARRYB_26_24_port, S => 
                           SUMB_26_24_port);
   S2_26_25 : FA_X1 port map( A => ab_26_25_port, B => CARRYB_25_25_port, CI =>
                           SUMB_25_26_port, CO => CARRYB_26_25_port, S => 
                           SUMB_26_25_port);
   S2_26_26 : FA_X1 port map( A => ab_26_26_port, B => CARRYB_25_26_port, CI =>
                           SUMB_25_27_port, CO => CARRYB_26_26_port, S => 
                           SUMB_26_26_port);
   S2_26_27 : FA_X1 port map( A => ab_26_27_port, B => CARRYB_25_27_port, CI =>
                           SUMB_25_28_port, CO => CARRYB_26_27_port, S => 
                           SUMB_26_27_port);
   S2_26_28 : FA_X1 port map( A => ab_26_28_port, B => CARRYB_25_28_port, CI =>
                           SUMB_25_29_port, CO => CARRYB_26_28_port, S => 
                           SUMB_26_28_port);
   S2_26_29 : FA_X1 port map( A => ab_26_29_port, B => CARRYB_25_29_port, CI =>
                           SUMB_25_30_port, CO => CARRYB_26_29_port, S => 
                           SUMB_26_29_port);
   S3_26_30 : FA_X1 port map( A => ab_26_30_port, B => CARRYB_25_30_port, CI =>
                           ab_25_31_port, CO => CARRYB_26_30_port, S => 
                           SUMB_26_30_port);
   S1_25_0 : FA_X1 port map( A => ab_25_0_port, B => CARRYB_24_0_port, CI => 
                           SUMB_24_1_port, CO => CARRYB_25_0_port, S => 
                           A1_23_port);
   S2_25_1 : FA_X1 port map( A => ab_25_1_port, B => CARRYB_24_1_port, CI => 
                           SUMB_24_2_port, CO => CARRYB_25_1_port, S => 
                           SUMB_25_1_port);
   S2_25_2 : FA_X1 port map( A => ab_25_2_port, B => CARRYB_24_2_port, CI => 
                           SUMB_24_3_port, CO => CARRYB_25_2_port, S => 
                           SUMB_25_2_port);
   S2_25_3 : FA_X1 port map( A => ab_25_3_port, B => CARRYB_24_3_port, CI => 
                           SUMB_24_4_port, CO => CARRYB_25_3_port, S => 
                           SUMB_25_3_port);
   S2_25_4 : FA_X1 port map( A => ab_25_4_port, B => CARRYB_24_4_port, CI => 
                           SUMB_24_5_port, CO => CARRYB_25_4_port, S => 
                           SUMB_25_4_port);
   S2_25_5 : FA_X1 port map( A => ab_25_5_port, B => CARRYB_24_5_port, CI => 
                           SUMB_24_6_port, CO => CARRYB_25_5_port, S => 
                           SUMB_25_5_port);
   S2_25_6 : FA_X1 port map( A => ab_25_6_port, B => CARRYB_24_6_port, CI => 
                           SUMB_24_7_port, CO => CARRYB_25_6_port, S => 
                           SUMB_25_6_port);
   S2_25_7 : FA_X1 port map( A => ab_25_7_port, B => CARRYB_24_7_port, CI => 
                           SUMB_24_8_port, CO => CARRYB_25_7_port, S => 
                           SUMB_25_7_port);
   S2_25_8 : FA_X1 port map( A => ab_25_8_port, B => CARRYB_24_8_port, CI => 
                           SUMB_24_9_port, CO => CARRYB_25_8_port, S => 
                           SUMB_25_8_port);
   S2_25_9 : FA_X1 port map( A => ab_25_9_port, B => CARRYB_24_9_port, CI => 
                           SUMB_24_10_port, CO => CARRYB_25_9_port, S => 
                           SUMB_25_9_port);
   S2_25_10 : FA_X1 port map( A => ab_25_10_port, B => CARRYB_24_10_port, CI =>
                           SUMB_24_11_port, CO => CARRYB_25_10_port, S => 
                           SUMB_25_10_port);
   S2_25_11 : FA_X1 port map( A => ab_25_11_port, B => CARRYB_24_11_port, CI =>
                           SUMB_24_12_port, CO => CARRYB_25_11_port, S => 
                           SUMB_25_11_port);
   S2_25_12 : FA_X1 port map( A => ab_25_12_port, B => CARRYB_24_12_port, CI =>
                           SUMB_24_13_port, CO => CARRYB_25_12_port, S => 
                           SUMB_25_12_port);
   S2_25_13 : FA_X1 port map( A => ab_25_13_port, B => CARRYB_24_13_port, CI =>
                           SUMB_24_14_port, CO => CARRYB_25_13_port, S => 
                           SUMB_25_13_port);
   S2_25_14 : FA_X1 port map( A => ab_25_14_port, B => CARRYB_24_14_port, CI =>
                           SUMB_24_15_port, CO => CARRYB_25_14_port, S => 
                           SUMB_25_14_port);
   S2_25_15 : FA_X1 port map( A => ab_25_15_port, B => CARRYB_24_15_port, CI =>
                           SUMB_24_16_port, CO => CARRYB_25_15_port, S => 
                           SUMB_25_15_port);
   S2_25_16 : FA_X1 port map( A => ab_25_16_port, B => CARRYB_24_16_port, CI =>
                           SUMB_24_17_port, CO => CARRYB_25_16_port, S => 
                           SUMB_25_16_port);
   S2_25_17 : FA_X1 port map( A => ab_25_17_port, B => CARRYB_24_17_port, CI =>
                           SUMB_24_18_port, CO => CARRYB_25_17_port, S => 
                           SUMB_25_17_port);
   S2_25_18 : FA_X1 port map( A => ab_25_18_port, B => CARRYB_24_18_port, CI =>
                           SUMB_24_19_port, CO => CARRYB_25_18_port, S => 
                           SUMB_25_18_port);
   S2_25_19 : FA_X1 port map( A => ab_25_19_port, B => CARRYB_24_19_port, CI =>
                           SUMB_24_20_port, CO => CARRYB_25_19_port, S => 
                           SUMB_25_19_port);
   S2_25_20 : FA_X1 port map( A => ab_25_20_port, B => CARRYB_24_20_port, CI =>
                           SUMB_24_21_port, CO => CARRYB_25_20_port, S => 
                           SUMB_25_20_port);
   S2_25_21 : FA_X1 port map( A => ab_25_21_port, B => CARRYB_24_21_port, CI =>
                           SUMB_24_22_port, CO => CARRYB_25_21_port, S => 
                           SUMB_25_21_port);
   S2_25_22 : FA_X1 port map( A => ab_25_22_port, B => CARRYB_24_22_port, CI =>
                           SUMB_24_23_port, CO => CARRYB_25_22_port, S => 
                           SUMB_25_22_port);
   S2_25_23 : FA_X1 port map( A => ab_25_23_port, B => CARRYB_24_23_port, CI =>
                           SUMB_24_24_port, CO => CARRYB_25_23_port, S => 
                           SUMB_25_23_port);
   S2_25_24 : FA_X1 port map( A => ab_25_24_port, B => CARRYB_24_24_port, CI =>
                           SUMB_24_25_port, CO => CARRYB_25_24_port, S => 
                           SUMB_25_24_port);
   S2_25_25 : FA_X1 port map( A => ab_25_25_port, B => CARRYB_24_25_port, CI =>
                           SUMB_24_26_port, CO => CARRYB_25_25_port, S => 
                           SUMB_25_25_port);
   S2_25_26 : FA_X1 port map( A => ab_25_26_port, B => CARRYB_24_26_port, CI =>
                           SUMB_24_27_port, CO => CARRYB_25_26_port, S => 
                           SUMB_25_26_port);
   S2_25_27 : FA_X1 port map( A => ab_25_27_port, B => CARRYB_24_27_port, CI =>
                           SUMB_24_28_port, CO => CARRYB_25_27_port, S => 
                           SUMB_25_27_port);
   S2_25_28 : FA_X1 port map( A => ab_25_28_port, B => CARRYB_24_28_port, CI =>
                           SUMB_24_29_port, CO => CARRYB_25_28_port, S => 
                           SUMB_25_28_port);
   S2_25_29 : FA_X1 port map( A => ab_25_29_port, B => CARRYB_24_29_port, CI =>
                           SUMB_24_30_port, CO => CARRYB_25_29_port, S => 
                           SUMB_25_29_port);
   S3_25_30 : FA_X1 port map( A => ab_25_30_port, B => CARRYB_24_30_port, CI =>
                           ab_24_31_port, CO => CARRYB_25_30_port, S => 
                           SUMB_25_30_port);
   S1_24_0 : FA_X1 port map( A => ab_24_0_port, B => CARRYB_23_0_port, CI => 
                           SUMB_23_1_port, CO => CARRYB_24_0_port, S => 
                           A1_22_port);
   S2_24_1 : FA_X1 port map( A => ab_24_1_port, B => CARRYB_23_1_port, CI => 
                           SUMB_23_2_port, CO => CARRYB_24_1_port, S => 
                           SUMB_24_1_port);
   S2_24_2 : FA_X1 port map( A => ab_24_2_port, B => CARRYB_23_2_port, CI => 
                           SUMB_23_3_port, CO => CARRYB_24_2_port, S => 
                           SUMB_24_2_port);
   S2_24_3 : FA_X1 port map( A => ab_24_3_port, B => CARRYB_23_3_port, CI => 
                           SUMB_23_4_port, CO => CARRYB_24_3_port, S => 
                           SUMB_24_3_port);
   S2_24_4 : FA_X1 port map( A => ab_24_4_port, B => CARRYB_23_4_port, CI => 
                           SUMB_23_5_port, CO => CARRYB_24_4_port, S => 
                           SUMB_24_4_port);
   S2_24_5 : FA_X1 port map( A => ab_24_5_port, B => CARRYB_23_5_port, CI => 
                           SUMB_23_6_port, CO => CARRYB_24_5_port, S => 
                           SUMB_24_5_port);
   S2_24_6 : FA_X1 port map( A => ab_24_6_port, B => CARRYB_23_6_port, CI => 
                           SUMB_23_7_port, CO => CARRYB_24_6_port, S => 
                           SUMB_24_6_port);
   S2_24_7 : FA_X1 port map( A => ab_24_7_port, B => CARRYB_23_7_port, CI => 
                           SUMB_23_8_port, CO => CARRYB_24_7_port, S => 
                           SUMB_24_7_port);
   S2_24_8 : FA_X1 port map( A => ab_24_8_port, B => CARRYB_23_8_port, CI => 
                           SUMB_23_9_port, CO => CARRYB_24_8_port, S => 
                           SUMB_24_8_port);
   S2_24_9 : FA_X1 port map( A => ab_24_9_port, B => CARRYB_23_9_port, CI => 
                           SUMB_23_10_port, CO => CARRYB_24_9_port, S => 
                           SUMB_24_9_port);
   S2_24_10 : FA_X1 port map( A => ab_24_10_port, B => CARRYB_23_10_port, CI =>
                           SUMB_23_11_port, CO => CARRYB_24_10_port, S => 
                           SUMB_24_10_port);
   S2_24_11 : FA_X1 port map( A => ab_24_11_port, B => CARRYB_23_11_port, CI =>
                           SUMB_23_12_port, CO => CARRYB_24_11_port, S => 
                           SUMB_24_11_port);
   S2_24_12 : FA_X1 port map( A => ab_24_12_port, B => CARRYB_23_12_port, CI =>
                           SUMB_23_13_port, CO => CARRYB_24_12_port, S => 
                           SUMB_24_12_port);
   S2_24_13 : FA_X1 port map( A => ab_24_13_port, B => CARRYB_23_13_port, CI =>
                           SUMB_23_14_port, CO => CARRYB_24_13_port, S => 
                           SUMB_24_13_port);
   S2_24_14 : FA_X1 port map( A => ab_24_14_port, B => CARRYB_23_14_port, CI =>
                           SUMB_23_15_port, CO => CARRYB_24_14_port, S => 
                           SUMB_24_14_port);
   S2_24_15 : FA_X1 port map( A => ab_24_15_port, B => CARRYB_23_15_port, CI =>
                           SUMB_23_16_port, CO => CARRYB_24_15_port, S => 
                           SUMB_24_15_port);
   S2_24_16 : FA_X1 port map( A => ab_24_16_port, B => CARRYB_23_16_port, CI =>
                           SUMB_23_17_port, CO => CARRYB_24_16_port, S => 
                           SUMB_24_16_port);
   S2_24_17 : FA_X1 port map( A => ab_24_17_port, B => CARRYB_23_17_port, CI =>
                           SUMB_23_18_port, CO => CARRYB_24_17_port, S => 
                           SUMB_24_17_port);
   S2_24_18 : FA_X1 port map( A => ab_24_18_port, B => CARRYB_23_18_port, CI =>
                           SUMB_23_19_port, CO => CARRYB_24_18_port, S => 
                           SUMB_24_18_port);
   S2_24_19 : FA_X1 port map( A => ab_24_19_port, B => CARRYB_23_19_port, CI =>
                           SUMB_23_20_port, CO => CARRYB_24_19_port, S => 
                           SUMB_24_19_port);
   S2_24_20 : FA_X1 port map( A => ab_24_20_port, B => CARRYB_23_20_port, CI =>
                           SUMB_23_21_port, CO => CARRYB_24_20_port, S => 
                           SUMB_24_20_port);
   S2_24_21 : FA_X1 port map( A => ab_24_21_port, B => CARRYB_23_21_port, CI =>
                           SUMB_23_22_port, CO => CARRYB_24_21_port, S => 
                           SUMB_24_21_port);
   S2_24_22 : FA_X1 port map( A => ab_24_22_port, B => CARRYB_23_22_port, CI =>
                           SUMB_23_23_port, CO => CARRYB_24_22_port, S => 
                           SUMB_24_22_port);
   S2_24_23 : FA_X1 port map( A => ab_24_23_port, B => CARRYB_23_23_port, CI =>
                           SUMB_23_24_port, CO => CARRYB_24_23_port, S => 
                           SUMB_24_23_port);
   S2_24_24 : FA_X1 port map( A => ab_24_24_port, B => CARRYB_23_24_port, CI =>
                           SUMB_23_25_port, CO => CARRYB_24_24_port, S => 
                           SUMB_24_24_port);
   S2_24_25 : FA_X1 port map( A => ab_24_25_port, B => CARRYB_23_25_port, CI =>
                           SUMB_23_26_port, CO => CARRYB_24_25_port, S => 
                           SUMB_24_25_port);
   S2_24_26 : FA_X1 port map( A => ab_24_26_port, B => CARRYB_23_26_port, CI =>
                           SUMB_23_27_port, CO => CARRYB_24_26_port, S => 
                           SUMB_24_26_port);
   S2_24_27 : FA_X1 port map( A => ab_24_27_port, B => CARRYB_23_27_port, CI =>
                           SUMB_23_28_port, CO => CARRYB_24_27_port, S => 
                           SUMB_24_27_port);
   S2_24_28 : FA_X1 port map( A => ab_24_28_port, B => CARRYB_23_28_port, CI =>
                           SUMB_23_29_port, CO => CARRYB_24_28_port, S => 
                           SUMB_24_28_port);
   S2_24_29 : FA_X1 port map( A => ab_24_29_port, B => CARRYB_23_29_port, CI =>
                           SUMB_23_30_port, CO => CARRYB_24_29_port, S => 
                           SUMB_24_29_port);
   S3_24_30 : FA_X1 port map( A => ab_24_30_port, B => CARRYB_23_30_port, CI =>
                           ab_23_31_port, CO => CARRYB_24_30_port, S => 
                           SUMB_24_30_port);
   S1_23_0 : FA_X1 port map( A => ab_23_0_port, B => CARRYB_22_0_port, CI => 
                           SUMB_22_1_port, CO => CARRYB_23_0_port, S => 
                           A1_21_port);
   S2_23_1 : FA_X1 port map( A => ab_23_1_port, B => CARRYB_22_1_port, CI => 
                           SUMB_22_2_port, CO => CARRYB_23_1_port, S => 
                           SUMB_23_1_port);
   S2_23_2 : FA_X1 port map( A => ab_23_2_port, B => CARRYB_22_2_port, CI => 
                           SUMB_22_3_port, CO => CARRYB_23_2_port, S => 
                           SUMB_23_2_port);
   S2_23_3 : FA_X1 port map( A => ab_23_3_port, B => CARRYB_22_3_port, CI => 
                           SUMB_22_4_port, CO => CARRYB_23_3_port, S => 
                           SUMB_23_3_port);
   S2_23_4 : FA_X1 port map( A => ab_23_4_port, B => CARRYB_22_4_port, CI => 
                           SUMB_22_5_port, CO => CARRYB_23_4_port, S => 
                           SUMB_23_4_port);
   S2_23_5 : FA_X1 port map( A => ab_23_5_port, B => CARRYB_22_5_port, CI => 
                           SUMB_22_6_port, CO => CARRYB_23_5_port, S => 
                           SUMB_23_5_port);
   S2_23_6 : FA_X1 port map( A => ab_23_6_port, B => CARRYB_22_6_port, CI => 
                           SUMB_22_7_port, CO => CARRYB_23_6_port, S => 
                           SUMB_23_6_port);
   S2_23_7 : FA_X1 port map( A => ab_23_7_port, B => CARRYB_22_7_port, CI => 
                           SUMB_22_8_port, CO => CARRYB_23_7_port, S => 
                           SUMB_23_7_port);
   S2_23_8 : FA_X1 port map( A => ab_23_8_port, B => CARRYB_22_8_port, CI => 
                           SUMB_22_9_port, CO => CARRYB_23_8_port, S => 
                           SUMB_23_8_port);
   S2_23_9 : FA_X1 port map( A => ab_23_9_port, B => CARRYB_22_9_port, CI => 
                           SUMB_22_10_port, CO => CARRYB_23_9_port, S => 
                           SUMB_23_9_port);
   S2_23_10 : FA_X1 port map( A => ab_23_10_port, B => CARRYB_22_10_port, CI =>
                           SUMB_22_11_port, CO => CARRYB_23_10_port, S => 
                           SUMB_23_10_port);
   S2_23_11 : FA_X1 port map( A => ab_23_11_port, B => CARRYB_22_11_port, CI =>
                           SUMB_22_12_port, CO => CARRYB_23_11_port, S => 
                           SUMB_23_11_port);
   S2_23_12 : FA_X1 port map( A => ab_23_12_port, B => CARRYB_22_12_port, CI =>
                           SUMB_22_13_port, CO => CARRYB_23_12_port, S => 
                           SUMB_23_12_port);
   S2_23_13 : FA_X1 port map( A => ab_23_13_port, B => CARRYB_22_13_port, CI =>
                           SUMB_22_14_port, CO => CARRYB_23_13_port, S => 
                           SUMB_23_13_port);
   S2_23_14 : FA_X1 port map( A => ab_23_14_port, B => CARRYB_22_14_port, CI =>
                           SUMB_22_15_port, CO => CARRYB_23_14_port, S => 
                           SUMB_23_14_port);
   S2_23_15 : FA_X1 port map( A => ab_23_15_port, B => CARRYB_22_15_port, CI =>
                           SUMB_22_16_port, CO => CARRYB_23_15_port, S => 
                           SUMB_23_15_port);
   S2_23_16 : FA_X1 port map( A => ab_23_16_port, B => CARRYB_22_16_port, CI =>
                           SUMB_22_17_port, CO => CARRYB_23_16_port, S => 
                           SUMB_23_16_port);
   S2_23_17 : FA_X1 port map( A => ab_23_17_port, B => CARRYB_22_17_port, CI =>
                           SUMB_22_18_port, CO => CARRYB_23_17_port, S => 
                           SUMB_23_17_port);
   S2_23_18 : FA_X1 port map( A => ab_23_18_port, B => CARRYB_22_18_port, CI =>
                           SUMB_22_19_port, CO => CARRYB_23_18_port, S => 
                           SUMB_23_18_port);
   S2_23_19 : FA_X1 port map( A => ab_23_19_port, B => CARRYB_22_19_port, CI =>
                           SUMB_22_20_port, CO => CARRYB_23_19_port, S => 
                           SUMB_23_19_port);
   S2_23_20 : FA_X1 port map( A => ab_23_20_port, B => CARRYB_22_20_port, CI =>
                           SUMB_22_21_port, CO => CARRYB_23_20_port, S => 
                           SUMB_23_20_port);
   S2_23_21 : FA_X1 port map( A => ab_23_21_port, B => CARRYB_22_21_port, CI =>
                           SUMB_22_22_port, CO => CARRYB_23_21_port, S => 
                           SUMB_23_21_port);
   S2_23_22 : FA_X1 port map( A => ab_23_22_port, B => CARRYB_22_22_port, CI =>
                           SUMB_22_23_port, CO => CARRYB_23_22_port, S => 
                           SUMB_23_22_port);
   S2_23_23 : FA_X1 port map( A => ab_23_23_port, B => CARRYB_22_23_port, CI =>
                           SUMB_22_24_port, CO => CARRYB_23_23_port, S => 
                           SUMB_23_23_port);
   S2_23_24 : FA_X1 port map( A => ab_23_24_port, B => CARRYB_22_24_port, CI =>
                           SUMB_22_25_port, CO => CARRYB_23_24_port, S => 
                           SUMB_23_24_port);
   S2_23_25 : FA_X1 port map( A => ab_23_25_port, B => CARRYB_22_25_port, CI =>
                           SUMB_22_26_port, CO => CARRYB_23_25_port, S => 
                           SUMB_23_25_port);
   S2_23_26 : FA_X1 port map( A => ab_23_26_port, B => CARRYB_22_26_port, CI =>
                           SUMB_22_27_port, CO => CARRYB_23_26_port, S => 
                           SUMB_23_26_port);
   S2_23_27 : FA_X1 port map( A => ab_23_27_port, B => CARRYB_22_27_port, CI =>
                           SUMB_22_28_port, CO => CARRYB_23_27_port, S => 
                           SUMB_23_27_port);
   S2_23_28 : FA_X1 port map( A => ab_23_28_port, B => CARRYB_22_28_port, CI =>
                           SUMB_22_29_port, CO => CARRYB_23_28_port, S => 
                           SUMB_23_28_port);
   S2_23_29 : FA_X1 port map( A => ab_23_29_port, B => CARRYB_22_29_port, CI =>
                           SUMB_22_30_port, CO => CARRYB_23_29_port, S => 
                           SUMB_23_29_port);
   S3_23_30 : FA_X1 port map( A => ab_23_30_port, B => CARRYB_22_30_port, CI =>
                           ab_22_31_port, CO => CARRYB_23_30_port, S => 
                           SUMB_23_30_port);
   S1_22_0 : FA_X1 port map( A => ab_22_0_port, B => CARRYB_21_0_port, CI => 
                           SUMB_21_1_port, CO => CARRYB_22_0_port, S => 
                           A1_20_port);
   S2_22_1 : FA_X1 port map( A => ab_22_1_port, B => CARRYB_21_1_port, CI => 
                           SUMB_21_2_port, CO => CARRYB_22_1_port, S => 
                           SUMB_22_1_port);
   S2_22_2 : FA_X1 port map( A => ab_22_2_port, B => CARRYB_21_2_port, CI => 
                           SUMB_21_3_port, CO => CARRYB_22_2_port, S => 
                           SUMB_22_2_port);
   S2_22_3 : FA_X1 port map( A => ab_22_3_port, B => CARRYB_21_3_port, CI => 
                           SUMB_21_4_port, CO => CARRYB_22_3_port, S => 
                           SUMB_22_3_port);
   S2_22_4 : FA_X1 port map( A => ab_22_4_port, B => CARRYB_21_4_port, CI => 
                           SUMB_21_5_port, CO => CARRYB_22_4_port, S => 
                           SUMB_22_4_port);
   S2_22_5 : FA_X1 port map( A => ab_22_5_port, B => CARRYB_21_5_port, CI => 
                           SUMB_21_6_port, CO => CARRYB_22_5_port, S => 
                           SUMB_22_5_port);
   S2_22_6 : FA_X1 port map( A => ab_22_6_port, B => CARRYB_21_6_port, CI => 
                           SUMB_21_7_port, CO => CARRYB_22_6_port, S => 
                           SUMB_22_6_port);
   S2_22_7 : FA_X1 port map( A => ab_22_7_port, B => CARRYB_21_7_port, CI => 
                           SUMB_21_8_port, CO => CARRYB_22_7_port, S => 
                           SUMB_22_7_port);
   S2_22_8 : FA_X1 port map( A => ab_22_8_port, B => CARRYB_21_8_port, CI => 
                           SUMB_21_9_port, CO => CARRYB_22_8_port, S => 
                           SUMB_22_8_port);
   S2_22_9 : FA_X1 port map( A => ab_22_9_port, B => CARRYB_21_9_port, CI => 
                           SUMB_21_10_port, CO => CARRYB_22_9_port, S => 
                           SUMB_22_9_port);
   S2_22_10 : FA_X1 port map( A => ab_22_10_port, B => CARRYB_21_10_port, CI =>
                           SUMB_21_11_port, CO => CARRYB_22_10_port, S => 
                           SUMB_22_10_port);
   S2_22_11 : FA_X1 port map( A => ab_22_11_port, B => CARRYB_21_11_port, CI =>
                           SUMB_21_12_port, CO => CARRYB_22_11_port, S => 
                           SUMB_22_11_port);
   S2_22_12 : FA_X1 port map( A => ab_22_12_port, B => CARRYB_21_12_port, CI =>
                           SUMB_21_13_port, CO => CARRYB_22_12_port, S => 
                           SUMB_22_12_port);
   S2_22_13 : FA_X1 port map( A => ab_22_13_port, B => CARRYB_21_13_port, CI =>
                           SUMB_21_14_port, CO => CARRYB_22_13_port, S => 
                           SUMB_22_13_port);
   S2_22_14 : FA_X1 port map( A => ab_22_14_port, B => CARRYB_21_14_port, CI =>
                           SUMB_21_15_port, CO => CARRYB_22_14_port, S => 
                           SUMB_22_14_port);
   S2_22_15 : FA_X1 port map( A => ab_22_15_port, B => CARRYB_21_15_port, CI =>
                           SUMB_21_16_port, CO => CARRYB_22_15_port, S => 
                           SUMB_22_15_port);
   S2_22_16 : FA_X1 port map( A => ab_22_16_port, B => CARRYB_21_16_port, CI =>
                           SUMB_21_17_port, CO => CARRYB_22_16_port, S => 
                           SUMB_22_16_port);
   S2_22_17 : FA_X1 port map( A => ab_22_17_port, B => CARRYB_21_17_port, CI =>
                           SUMB_21_18_port, CO => CARRYB_22_17_port, S => 
                           SUMB_22_17_port);
   S2_22_18 : FA_X1 port map( A => ab_22_18_port, B => CARRYB_21_18_port, CI =>
                           SUMB_21_19_port, CO => CARRYB_22_18_port, S => 
                           SUMB_22_18_port);
   S2_22_19 : FA_X1 port map( A => ab_22_19_port, B => CARRYB_21_19_port, CI =>
                           SUMB_21_20_port, CO => CARRYB_22_19_port, S => 
                           SUMB_22_19_port);
   S2_22_20 : FA_X1 port map( A => ab_22_20_port, B => CARRYB_21_20_port, CI =>
                           SUMB_21_21_port, CO => CARRYB_22_20_port, S => 
                           SUMB_22_20_port);
   S2_22_21 : FA_X1 port map( A => ab_22_21_port, B => CARRYB_21_21_port, CI =>
                           SUMB_21_22_port, CO => CARRYB_22_21_port, S => 
                           SUMB_22_21_port);
   S2_22_22 : FA_X1 port map( A => ab_22_22_port, B => CARRYB_21_22_port, CI =>
                           SUMB_21_23_port, CO => CARRYB_22_22_port, S => 
                           SUMB_22_22_port);
   S2_22_23 : FA_X1 port map( A => ab_22_23_port, B => CARRYB_21_23_port, CI =>
                           SUMB_21_24_port, CO => CARRYB_22_23_port, S => 
                           SUMB_22_23_port);
   S2_22_24 : FA_X1 port map( A => ab_22_24_port, B => CARRYB_21_24_port, CI =>
                           SUMB_21_25_port, CO => CARRYB_22_24_port, S => 
                           SUMB_22_24_port);
   S2_22_25 : FA_X1 port map( A => ab_22_25_port, B => CARRYB_21_25_port, CI =>
                           SUMB_21_26_port, CO => CARRYB_22_25_port, S => 
                           SUMB_22_25_port);
   S2_22_26 : FA_X1 port map( A => ab_22_26_port, B => CARRYB_21_26_port, CI =>
                           SUMB_21_27_port, CO => CARRYB_22_26_port, S => 
                           SUMB_22_26_port);
   S2_22_27 : FA_X1 port map( A => ab_22_27_port, B => CARRYB_21_27_port, CI =>
                           SUMB_21_28_port, CO => CARRYB_22_27_port, S => 
                           SUMB_22_27_port);
   S2_22_28 : FA_X1 port map( A => ab_22_28_port, B => CARRYB_21_28_port, CI =>
                           SUMB_21_29_port, CO => CARRYB_22_28_port, S => 
                           SUMB_22_28_port);
   S2_22_29 : FA_X1 port map( A => ab_22_29_port, B => CARRYB_21_29_port, CI =>
                           SUMB_21_30_port, CO => CARRYB_22_29_port, S => 
                           SUMB_22_29_port);
   S3_22_30 : FA_X1 port map( A => ab_22_30_port, B => CARRYB_21_30_port, CI =>
                           ab_21_31_port, CO => CARRYB_22_30_port, S => 
                           SUMB_22_30_port);
   S1_21_0 : FA_X1 port map( A => ab_21_0_port, B => CARRYB_20_0_port, CI => 
                           SUMB_20_1_port, CO => CARRYB_21_0_port, S => 
                           A1_19_port);
   S2_21_1 : FA_X1 port map( A => ab_21_1_port, B => CARRYB_20_1_port, CI => 
                           SUMB_20_2_port, CO => CARRYB_21_1_port, S => 
                           SUMB_21_1_port);
   S2_21_2 : FA_X1 port map( A => ab_21_2_port, B => CARRYB_20_2_port, CI => 
                           SUMB_20_3_port, CO => CARRYB_21_2_port, S => 
                           SUMB_21_2_port);
   S2_21_3 : FA_X1 port map( A => ab_21_3_port, B => CARRYB_20_3_port, CI => 
                           SUMB_20_4_port, CO => CARRYB_21_3_port, S => 
                           SUMB_21_3_port);
   S2_21_4 : FA_X1 port map( A => ab_21_4_port, B => CARRYB_20_4_port, CI => 
                           SUMB_20_5_port, CO => CARRYB_21_4_port, S => 
                           SUMB_21_4_port);
   S2_21_5 : FA_X1 port map( A => ab_21_5_port, B => CARRYB_20_5_port, CI => 
                           SUMB_20_6_port, CO => CARRYB_21_5_port, S => 
                           SUMB_21_5_port);
   S2_21_6 : FA_X1 port map( A => ab_21_6_port, B => CARRYB_20_6_port, CI => 
                           SUMB_20_7_port, CO => CARRYB_21_6_port, S => 
                           SUMB_21_6_port);
   S2_21_7 : FA_X1 port map( A => ab_21_7_port, B => CARRYB_20_7_port, CI => 
                           SUMB_20_8_port, CO => CARRYB_21_7_port, S => 
                           SUMB_21_7_port);
   S2_21_8 : FA_X1 port map( A => ab_21_8_port, B => CARRYB_20_8_port, CI => 
                           SUMB_20_9_port, CO => CARRYB_21_8_port, S => 
                           SUMB_21_8_port);
   S2_21_9 : FA_X1 port map( A => ab_21_9_port, B => CARRYB_20_9_port, CI => 
                           SUMB_20_10_port, CO => CARRYB_21_9_port, S => 
                           SUMB_21_9_port);
   S2_21_10 : FA_X1 port map( A => ab_21_10_port, B => CARRYB_20_10_port, CI =>
                           SUMB_20_11_port, CO => CARRYB_21_10_port, S => 
                           SUMB_21_10_port);
   S2_21_11 : FA_X1 port map( A => ab_21_11_port, B => CARRYB_20_11_port, CI =>
                           SUMB_20_12_port, CO => CARRYB_21_11_port, S => 
                           SUMB_21_11_port);
   S2_21_12 : FA_X1 port map( A => ab_21_12_port, B => CARRYB_20_12_port, CI =>
                           SUMB_20_13_port, CO => CARRYB_21_12_port, S => 
                           SUMB_21_12_port);
   S2_21_13 : FA_X1 port map( A => ab_21_13_port, B => CARRYB_20_13_port, CI =>
                           SUMB_20_14_port, CO => CARRYB_21_13_port, S => 
                           SUMB_21_13_port);
   S2_21_14 : FA_X1 port map( A => ab_21_14_port, B => CARRYB_20_14_port, CI =>
                           SUMB_20_15_port, CO => CARRYB_21_14_port, S => 
                           SUMB_21_14_port);
   S2_21_15 : FA_X1 port map( A => ab_21_15_port, B => CARRYB_20_15_port, CI =>
                           SUMB_20_16_port, CO => CARRYB_21_15_port, S => 
                           SUMB_21_15_port);
   S2_21_16 : FA_X1 port map( A => ab_21_16_port, B => CARRYB_20_16_port, CI =>
                           SUMB_20_17_port, CO => CARRYB_21_16_port, S => 
                           SUMB_21_16_port);
   S2_21_17 : FA_X1 port map( A => ab_21_17_port, B => CARRYB_20_17_port, CI =>
                           SUMB_20_18_port, CO => CARRYB_21_17_port, S => 
                           SUMB_21_17_port);
   S2_21_18 : FA_X1 port map( A => ab_21_18_port, B => CARRYB_20_18_port, CI =>
                           SUMB_20_19_port, CO => CARRYB_21_18_port, S => 
                           SUMB_21_18_port);
   S2_21_19 : FA_X1 port map( A => ab_21_19_port, B => CARRYB_20_19_port, CI =>
                           SUMB_20_20_port, CO => CARRYB_21_19_port, S => 
                           SUMB_21_19_port);
   S2_21_20 : FA_X1 port map( A => ab_21_20_port, B => CARRYB_20_20_port, CI =>
                           SUMB_20_21_port, CO => CARRYB_21_20_port, S => 
                           SUMB_21_20_port);
   S2_21_21 : FA_X1 port map( A => ab_21_21_port, B => CARRYB_20_21_port, CI =>
                           SUMB_20_22_port, CO => CARRYB_21_21_port, S => 
                           SUMB_21_21_port);
   S2_21_22 : FA_X1 port map( A => ab_21_22_port, B => CARRYB_20_22_port, CI =>
                           SUMB_20_23_port, CO => CARRYB_21_22_port, S => 
                           SUMB_21_22_port);
   S2_21_23 : FA_X1 port map( A => ab_21_23_port, B => CARRYB_20_23_port, CI =>
                           SUMB_20_24_port, CO => CARRYB_21_23_port, S => 
                           SUMB_21_23_port);
   S2_21_24 : FA_X1 port map( A => ab_21_24_port, B => CARRYB_20_24_port, CI =>
                           SUMB_20_25_port, CO => CARRYB_21_24_port, S => 
                           SUMB_21_24_port);
   S2_21_25 : FA_X1 port map( A => ab_21_25_port, B => CARRYB_20_25_port, CI =>
                           SUMB_20_26_port, CO => CARRYB_21_25_port, S => 
                           SUMB_21_25_port);
   S2_21_26 : FA_X1 port map( A => ab_21_26_port, B => CARRYB_20_26_port, CI =>
                           SUMB_20_27_port, CO => CARRYB_21_26_port, S => 
                           SUMB_21_26_port);
   S2_21_27 : FA_X1 port map( A => ab_21_27_port, B => CARRYB_20_27_port, CI =>
                           SUMB_20_28_port, CO => CARRYB_21_27_port, S => 
                           SUMB_21_27_port);
   S2_21_28 : FA_X1 port map( A => ab_21_28_port, B => CARRYB_20_28_port, CI =>
                           SUMB_20_29_port, CO => CARRYB_21_28_port, S => 
                           SUMB_21_28_port);
   S2_21_29 : FA_X1 port map( A => ab_21_29_port, B => CARRYB_20_29_port, CI =>
                           SUMB_20_30_port, CO => CARRYB_21_29_port, S => 
                           SUMB_21_29_port);
   S3_21_30 : FA_X1 port map( A => ab_21_30_port, B => CARRYB_20_30_port, CI =>
                           ab_20_31_port, CO => CARRYB_21_30_port, S => 
                           SUMB_21_30_port);
   S1_20_0 : FA_X1 port map( A => ab_20_0_port, B => CARRYB_19_0_port, CI => 
                           SUMB_19_1_port, CO => CARRYB_20_0_port, S => 
                           A1_18_port);
   S2_20_1 : FA_X1 port map( A => ab_20_1_port, B => CARRYB_19_1_port, CI => 
                           SUMB_19_2_port, CO => CARRYB_20_1_port, S => 
                           SUMB_20_1_port);
   S2_20_2 : FA_X1 port map( A => ab_20_2_port, B => CARRYB_19_2_port, CI => 
                           SUMB_19_3_port, CO => CARRYB_20_2_port, S => 
                           SUMB_20_2_port);
   S2_20_3 : FA_X1 port map( A => ab_20_3_port, B => CARRYB_19_3_port, CI => 
                           SUMB_19_4_port, CO => CARRYB_20_3_port, S => 
                           SUMB_20_3_port);
   S2_20_4 : FA_X1 port map( A => ab_20_4_port, B => CARRYB_19_4_port, CI => 
                           SUMB_19_5_port, CO => CARRYB_20_4_port, S => 
                           SUMB_20_4_port);
   S2_20_5 : FA_X1 port map( A => ab_20_5_port, B => CARRYB_19_5_port, CI => 
                           SUMB_19_6_port, CO => CARRYB_20_5_port, S => 
                           SUMB_20_5_port);
   S2_20_6 : FA_X1 port map( A => ab_20_6_port, B => CARRYB_19_6_port, CI => 
                           SUMB_19_7_port, CO => CARRYB_20_6_port, S => 
                           SUMB_20_6_port);
   S2_20_7 : FA_X1 port map( A => ab_20_7_port, B => CARRYB_19_7_port, CI => 
                           SUMB_19_8_port, CO => CARRYB_20_7_port, S => 
                           SUMB_20_7_port);
   S2_20_8 : FA_X1 port map( A => ab_20_8_port, B => CARRYB_19_8_port, CI => 
                           SUMB_19_9_port, CO => CARRYB_20_8_port, S => 
                           SUMB_20_8_port);
   S2_20_9 : FA_X1 port map( A => ab_20_9_port, B => CARRYB_19_9_port, CI => 
                           SUMB_19_10_port, CO => CARRYB_20_9_port, S => 
                           SUMB_20_9_port);
   S2_20_10 : FA_X1 port map( A => ab_20_10_port, B => CARRYB_19_10_port, CI =>
                           SUMB_19_11_port, CO => CARRYB_20_10_port, S => 
                           SUMB_20_10_port);
   S2_20_11 : FA_X1 port map( A => ab_20_11_port, B => CARRYB_19_11_port, CI =>
                           SUMB_19_12_port, CO => CARRYB_20_11_port, S => 
                           SUMB_20_11_port);
   S2_20_12 : FA_X1 port map( A => ab_20_12_port, B => CARRYB_19_12_port, CI =>
                           SUMB_19_13_port, CO => CARRYB_20_12_port, S => 
                           SUMB_20_12_port);
   S2_20_13 : FA_X1 port map( A => ab_20_13_port, B => CARRYB_19_13_port, CI =>
                           SUMB_19_14_port, CO => CARRYB_20_13_port, S => 
                           SUMB_20_13_port);
   S2_20_14 : FA_X1 port map( A => ab_20_14_port, B => CARRYB_19_14_port, CI =>
                           SUMB_19_15_port, CO => CARRYB_20_14_port, S => 
                           SUMB_20_14_port);
   S2_20_15 : FA_X1 port map( A => ab_20_15_port, B => CARRYB_19_15_port, CI =>
                           SUMB_19_16_port, CO => CARRYB_20_15_port, S => 
                           SUMB_20_15_port);
   S2_20_16 : FA_X1 port map( A => ab_20_16_port, B => CARRYB_19_16_port, CI =>
                           SUMB_19_17_port, CO => CARRYB_20_16_port, S => 
                           SUMB_20_16_port);
   S2_20_17 : FA_X1 port map( A => ab_20_17_port, B => CARRYB_19_17_port, CI =>
                           SUMB_19_18_port, CO => CARRYB_20_17_port, S => 
                           SUMB_20_17_port);
   S2_20_18 : FA_X1 port map( A => ab_20_18_port, B => CARRYB_19_18_port, CI =>
                           SUMB_19_19_port, CO => CARRYB_20_18_port, S => 
                           SUMB_20_18_port);
   S2_20_19 : FA_X1 port map( A => ab_20_19_port, B => CARRYB_19_19_port, CI =>
                           SUMB_19_20_port, CO => CARRYB_20_19_port, S => 
                           SUMB_20_19_port);
   S2_20_20 : FA_X1 port map( A => ab_20_20_port, B => CARRYB_19_20_port, CI =>
                           SUMB_19_21_port, CO => CARRYB_20_20_port, S => 
                           SUMB_20_20_port);
   S2_20_21 : FA_X1 port map( A => ab_20_21_port, B => CARRYB_19_21_port, CI =>
                           SUMB_19_22_port, CO => CARRYB_20_21_port, S => 
                           SUMB_20_21_port);
   S2_20_22 : FA_X1 port map( A => ab_20_22_port, B => CARRYB_19_22_port, CI =>
                           SUMB_19_23_port, CO => CARRYB_20_22_port, S => 
                           SUMB_20_22_port);
   S2_20_23 : FA_X1 port map( A => ab_20_23_port, B => CARRYB_19_23_port, CI =>
                           SUMB_19_24_port, CO => CARRYB_20_23_port, S => 
                           SUMB_20_23_port);
   S2_20_24 : FA_X1 port map( A => ab_20_24_port, B => CARRYB_19_24_port, CI =>
                           SUMB_19_25_port, CO => CARRYB_20_24_port, S => 
                           SUMB_20_24_port);
   S2_20_25 : FA_X1 port map( A => ab_20_25_port, B => CARRYB_19_25_port, CI =>
                           SUMB_19_26_port, CO => CARRYB_20_25_port, S => 
                           SUMB_20_25_port);
   S2_20_26 : FA_X1 port map( A => ab_20_26_port, B => CARRYB_19_26_port, CI =>
                           SUMB_19_27_port, CO => CARRYB_20_26_port, S => 
                           SUMB_20_26_port);
   S2_20_27 : FA_X1 port map( A => ab_20_27_port, B => CARRYB_19_27_port, CI =>
                           SUMB_19_28_port, CO => CARRYB_20_27_port, S => 
                           SUMB_20_27_port);
   S2_20_28 : FA_X1 port map( A => ab_20_28_port, B => CARRYB_19_28_port, CI =>
                           SUMB_19_29_port, CO => CARRYB_20_28_port, S => 
                           SUMB_20_28_port);
   S2_20_29 : FA_X1 port map( A => ab_20_29_port, B => CARRYB_19_29_port, CI =>
                           SUMB_19_30_port, CO => CARRYB_20_29_port, S => 
                           SUMB_20_29_port);
   S3_20_30 : FA_X1 port map( A => ab_20_30_port, B => CARRYB_19_30_port, CI =>
                           ab_19_31_port, CO => CARRYB_20_30_port, S => 
                           SUMB_20_30_port);
   S1_19_0 : FA_X1 port map( A => ab_19_0_port, B => CARRYB_18_0_port, CI => 
                           SUMB_18_1_port, CO => CARRYB_19_0_port, S => 
                           A1_17_port);
   S2_19_1 : FA_X1 port map( A => ab_19_1_port, B => CARRYB_18_1_port, CI => 
                           SUMB_18_2_port, CO => CARRYB_19_1_port, S => 
                           SUMB_19_1_port);
   S2_19_2 : FA_X1 port map( A => ab_19_2_port, B => CARRYB_18_2_port, CI => 
                           SUMB_18_3_port, CO => CARRYB_19_2_port, S => 
                           SUMB_19_2_port);
   S2_19_3 : FA_X1 port map( A => ab_19_3_port, B => CARRYB_18_3_port, CI => 
                           SUMB_18_4_port, CO => CARRYB_19_3_port, S => 
                           SUMB_19_3_port);
   S2_19_4 : FA_X1 port map( A => ab_19_4_port, B => CARRYB_18_4_port, CI => 
                           SUMB_18_5_port, CO => CARRYB_19_4_port, S => 
                           SUMB_19_4_port);
   S2_19_5 : FA_X1 port map( A => ab_19_5_port, B => CARRYB_18_5_port, CI => 
                           SUMB_18_6_port, CO => CARRYB_19_5_port, S => 
                           SUMB_19_5_port);
   S2_19_6 : FA_X1 port map( A => ab_19_6_port, B => CARRYB_18_6_port, CI => 
                           SUMB_18_7_port, CO => CARRYB_19_6_port, S => 
                           SUMB_19_6_port);
   S2_19_7 : FA_X1 port map( A => ab_19_7_port, B => CARRYB_18_7_port, CI => 
                           SUMB_18_8_port, CO => CARRYB_19_7_port, S => 
                           SUMB_19_7_port);
   S2_19_8 : FA_X1 port map( A => ab_19_8_port, B => CARRYB_18_8_port, CI => 
                           SUMB_18_9_port, CO => CARRYB_19_8_port, S => 
                           SUMB_19_8_port);
   S2_19_9 : FA_X1 port map( A => ab_19_9_port, B => CARRYB_18_9_port, CI => 
                           SUMB_18_10_port, CO => CARRYB_19_9_port, S => 
                           SUMB_19_9_port);
   S2_19_10 : FA_X1 port map( A => ab_19_10_port, B => CARRYB_18_10_port, CI =>
                           SUMB_18_11_port, CO => CARRYB_19_10_port, S => 
                           SUMB_19_10_port);
   S2_19_11 : FA_X1 port map( A => ab_19_11_port, B => CARRYB_18_11_port, CI =>
                           SUMB_18_12_port, CO => CARRYB_19_11_port, S => 
                           SUMB_19_11_port);
   S2_19_12 : FA_X1 port map( A => ab_19_12_port, B => CARRYB_18_12_port, CI =>
                           SUMB_18_13_port, CO => CARRYB_19_12_port, S => 
                           SUMB_19_12_port);
   S2_19_13 : FA_X1 port map( A => ab_19_13_port, B => CARRYB_18_13_port, CI =>
                           SUMB_18_14_port, CO => CARRYB_19_13_port, S => 
                           SUMB_19_13_port);
   S2_19_14 : FA_X1 port map( A => ab_19_14_port, B => CARRYB_18_14_port, CI =>
                           SUMB_18_15_port, CO => CARRYB_19_14_port, S => 
                           SUMB_19_14_port);
   S2_19_15 : FA_X1 port map( A => ab_19_15_port, B => CARRYB_18_15_port, CI =>
                           SUMB_18_16_port, CO => CARRYB_19_15_port, S => 
                           SUMB_19_15_port);
   S2_19_16 : FA_X1 port map( A => ab_19_16_port, B => CARRYB_18_16_port, CI =>
                           SUMB_18_17_port, CO => CARRYB_19_16_port, S => 
                           SUMB_19_16_port);
   S2_19_17 : FA_X1 port map( A => ab_19_17_port, B => CARRYB_18_17_port, CI =>
                           SUMB_18_18_port, CO => CARRYB_19_17_port, S => 
                           SUMB_19_17_port);
   S2_19_18 : FA_X1 port map( A => ab_19_18_port, B => CARRYB_18_18_port, CI =>
                           SUMB_18_19_port, CO => CARRYB_19_18_port, S => 
                           SUMB_19_18_port);
   S2_19_19 : FA_X1 port map( A => ab_19_19_port, B => CARRYB_18_19_port, CI =>
                           SUMB_18_20_port, CO => CARRYB_19_19_port, S => 
                           SUMB_19_19_port);
   S2_19_20 : FA_X1 port map( A => ab_19_20_port, B => CARRYB_18_20_port, CI =>
                           SUMB_18_21_port, CO => CARRYB_19_20_port, S => 
                           SUMB_19_20_port);
   S2_19_21 : FA_X1 port map( A => ab_19_21_port, B => CARRYB_18_21_port, CI =>
                           SUMB_18_22_port, CO => CARRYB_19_21_port, S => 
                           SUMB_19_21_port);
   S2_19_22 : FA_X1 port map( A => ab_19_22_port, B => CARRYB_18_22_port, CI =>
                           SUMB_18_23_port, CO => CARRYB_19_22_port, S => 
                           SUMB_19_22_port);
   S2_19_23 : FA_X1 port map( A => ab_19_23_port, B => CARRYB_18_23_port, CI =>
                           SUMB_18_24_port, CO => CARRYB_19_23_port, S => 
                           SUMB_19_23_port);
   S2_19_24 : FA_X1 port map( A => ab_19_24_port, B => CARRYB_18_24_port, CI =>
                           SUMB_18_25_port, CO => CARRYB_19_24_port, S => 
                           SUMB_19_24_port);
   S2_19_25 : FA_X1 port map( A => ab_19_25_port, B => CARRYB_18_25_port, CI =>
                           SUMB_18_26_port, CO => CARRYB_19_25_port, S => 
                           SUMB_19_25_port);
   S2_19_26 : FA_X1 port map( A => ab_19_26_port, B => CARRYB_18_26_port, CI =>
                           SUMB_18_27_port, CO => CARRYB_19_26_port, S => 
                           SUMB_19_26_port);
   S2_19_27 : FA_X1 port map( A => ab_19_27_port, B => CARRYB_18_27_port, CI =>
                           SUMB_18_28_port, CO => CARRYB_19_27_port, S => 
                           SUMB_19_27_port);
   S2_19_28 : FA_X1 port map( A => ab_19_28_port, B => CARRYB_18_28_port, CI =>
                           SUMB_18_29_port, CO => CARRYB_19_28_port, S => 
                           SUMB_19_28_port);
   S2_19_29 : FA_X1 port map( A => ab_19_29_port, B => CARRYB_18_29_port, CI =>
                           SUMB_18_30_port, CO => CARRYB_19_29_port, S => 
                           SUMB_19_29_port);
   S3_19_30 : FA_X1 port map( A => ab_19_30_port, B => CARRYB_18_30_port, CI =>
                           ab_18_31_port, CO => CARRYB_19_30_port, S => 
                           SUMB_19_30_port);
   S1_18_0 : FA_X1 port map( A => ab_18_0_port, B => CARRYB_17_0_port, CI => 
                           SUMB_17_1_port, CO => CARRYB_18_0_port, S => 
                           A1_16_port);
   S2_18_1 : FA_X1 port map( A => ab_18_1_port, B => CARRYB_17_1_port, CI => 
                           SUMB_17_2_port, CO => CARRYB_18_1_port, S => 
                           SUMB_18_1_port);
   S2_18_2 : FA_X1 port map( A => ab_18_2_port, B => CARRYB_17_2_port, CI => 
                           SUMB_17_3_port, CO => CARRYB_18_2_port, S => 
                           SUMB_18_2_port);
   S2_18_3 : FA_X1 port map( A => ab_18_3_port, B => CARRYB_17_3_port, CI => 
                           SUMB_17_4_port, CO => CARRYB_18_3_port, S => 
                           SUMB_18_3_port);
   S2_18_4 : FA_X1 port map( A => ab_18_4_port, B => CARRYB_17_4_port, CI => 
                           SUMB_17_5_port, CO => CARRYB_18_4_port, S => 
                           SUMB_18_4_port);
   S2_18_5 : FA_X1 port map( A => ab_18_5_port, B => CARRYB_17_5_port, CI => 
                           SUMB_17_6_port, CO => CARRYB_18_5_port, S => 
                           SUMB_18_5_port);
   S2_18_6 : FA_X1 port map( A => ab_18_6_port, B => CARRYB_17_6_port, CI => 
                           SUMB_17_7_port, CO => CARRYB_18_6_port, S => 
                           SUMB_18_6_port);
   S2_18_7 : FA_X1 port map( A => ab_18_7_port, B => CARRYB_17_7_port, CI => 
                           SUMB_17_8_port, CO => CARRYB_18_7_port, S => 
                           SUMB_18_7_port);
   S2_18_8 : FA_X1 port map( A => ab_18_8_port, B => CARRYB_17_8_port, CI => 
                           SUMB_17_9_port, CO => CARRYB_18_8_port, S => 
                           SUMB_18_8_port);
   S2_18_9 : FA_X1 port map( A => ab_18_9_port, B => CARRYB_17_9_port, CI => 
                           SUMB_17_10_port, CO => CARRYB_18_9_port, S => 
                           SUMB_18_9_port);
   S2_18_10 : FA_X1 port map( A => ab_18_10_port, B => CARRYB_17_10_port, CI =>
                           SUMB_17_11_port, CO => CARRYB_18_10_port, S => 
                           SUMB_18_10_port);
   S2_18_11 : FA_X1 port map( A => ab_18_11_port, B => CARRYB_17_11_port, CI =>
                           SUMB_17_12_port, CO => CARRYB_18_11_port, S => 
                           SUMB_18_11_port);
   S2_18_12 : FA_X1 port map( A => ab_18_12_port, B => CARRYB_17_12_port, CI =>
                           SUMB_17_13_port, CO => CARRYB_18_12_port, S => 
                           SUMB_18_12_port);
   S2_18_13 : FA_X1 port map( A => ab_18_13_port, B => CARRYB_17_13_port, CI =>
                           SUMB_17_14_port, CO => CARRYB_18_13_port, S => 
                           SUMB_18_13_port);
   S2_18_14 : FA_X1 port map( A => ab_18_14_port, B => CARRYB_17_14_port, CI =>
                           SUMB_17_15_port, CO => CARRYB_18_14_port, S => 
                           SUMB_18_14_port);
   S2_18_15 : FA_X1 port map( A => ab_18_15_port, B => CARRYB_17_15_port, CI =>
                           SUMB_17_16_port, CO => CARRYB_18_15_port, S => 
                           SUMB_18_15_port);
   S2_18_16 : FA_X1 port map( A => ab_18_16_port, B => CARRYB_17_16_port, CI =>
                           SUMB_17_17_port, CO => CARRYB_18_16_port, S => 
                           SUMB_18_16_port);
   S2_18_17 : FA_X1 port map( A => ab_18_17_port, B => CARRYB_17_17_port, CI =>
                           SUMB_17_18_port, CO => CARRYB_18_17_port, S => 
                           SUMB_18_17_port);
   S2_18_18 : FA_X1 port map( A => ab_18_18_port, B => CARRYB_17_18_port, CI =>
                           SUMB_17_19_port, CO => CARRYB_18_18_port, S => 
                           SUMB_18_18_port);
   S2_18_19 : FA_X1 port map( A => ab_18_19_port, B => CARRYB_17_19_port, CI =>
                           SUMB_17_20_port, CO => CARRYB_18_19_port, S => 
                           SUMB_18_19_port);
   S2_18_20 : FA_X1 port map( A => ab_18_20_port, B => CARRYB_17_20_port, CI =>
                           SUMB_17_21_port, CO => CARRYB_18_20_port, S => 
                           SUMB_18_20_port);
   S2_18_21 : FA_X1 port map( A => ab_18_21_port, B => CARRYB_17_21_port, CI =>
                           SUMB_17_22_port, CO => CARRYB_18_21_port, S => 
                           SUMB_18_21_port);
   S2_18_22 : FA_X1 port map( A => ab_18_22_port, B => CARRYB_17_22_port, CI =>
                           SUMB_17_23_port, CO => CARRYB_18_22_port, S => 
                           SUMB_18_22_port);
   S2_18_23 : FA_X1 port map( A => ab_18_23_port, B => CARRYB_17_23_port, CI =>
                           SUMB_17_24_port, CO => CARRYB_18_23_port, S => 
                           SUMB_18_23_port);
   S2_18_24 : FA_X1 port map( A => ab_18_24_port, B => CARRYB_17_24_port, CI =>
                           SUMB_17_25_port, CO => CARRYB_18_24_port, S => 
                           SUMB_18_24_port);
   S2_18_25 : FA_X1 port map( A => ab_18_25_port, B => CARRYB_17_25_port, CI =>
                           SUMB_17_26_port, CO => CARRYB_18_25_port, S => 
                           SUMB_18_25_port);
   S2_18_26 : FA_X1 port map( A => ab_18_26_port, B => CARRYB_17_26_port, CI =>
                           SUMB_17_27_port, CO => CARRYB_18_26_port, S => 
                           SUMB_18_26_port);
   S2_18_27 : FA_X1 port map( A => ab_18_27_port, B => CARRYB_17_27_port, CI =>
                           SUMB_17_28_port, CO => CARRYB_18_27_port, S => 
                           SUMB_18_27_port);
   S2_18_28 : FA_X1 port map( A => ab_18_28_port, B => CARRYB_17_28_port, CI =>
                           SUMB_17_29_port, CO => CARRYB_18_28_port, S => 
                           SUMB_18_28_port);
   S2_18_29 : FA_X1 port map( A => ab_18_29_port, B => CARRYB_17_29_port, CI =>
                           SUMB_17_30_port, CO => CARRYB_18_29_port, S => 
                           SUMB_18_29_port);
   S3_18_30 : FA_X1 port map( A => ab_18_30_port, B => CARRYB_17_30_port, CI =>
                           ab_17_31_port, CO => CARRYB_18_30_port, S => 
                           SUMB_18_30_port);
   S1_17_0 : FA_X1 port map( A => ab_17_0_port, B => CARRYB_16_0_port, CI => 
                           SUMB_16_1_port, CO => CARRYB_17_0_port, S => 
                           A1_15_port);
   S2_17_1 : FA_X1 port map( A => ab_17_1_port, B => CARRYB_16_1_port, CI => 
                           SUMB_16_2_port, CO => CARRYB_17_1_port, S => 
                           SUMB_17_1_port);
   S2_17_2 : FA_X1 port map( A => ab_17_2_port, B => CARRYB_16_2_port, CI => 
                           SUMB_16_3_port, CO => CARRYB_17_2_port, S => 
                           SUMB_17_2_port);
   S2_17_3 : FA_X1 port map( A => ab_17_3_port, B => CARRYB_16_3_port, CI => 
                           SUMB_16_4_port, CO => CARRYB_17_3_port, S => 
                           SUMB_17_3_port);
   S2_17_4 : FA_X1 port map( A => ab_17_4_port, B => CARRYB_16_4_port, CI => 
                           SUMB_16_5_port, CO => CARRYB_17_4_port, S => 
                           SUMB_17_4_port);
   S2_17_5 : FA_X1 port map( A => ab_17_5_port, B => CARRYB_16_5_port, CI => 
                           SUMB_16_6_port, CO => CARRYB_17_5_port, S => 
                           SUMB_17_5_port);
   S2_17_6 : FA_X1 port map( A => ab_17_6_port, B => CARRYB_16_6_port, CI => 
                           SUMB_16_7_port, CO => CARRYB_17_6_port, S => 
                           SUMB_17_6_port);
   S2_17_7 : FA_X1 port map( A => ab_17_7_port, B => CARRYB_16_7_port, CI => 
                           SUMB_16_8_port, CO => CARRYB_17_7_port, S => 
                           SUMB_17_7_port);
   S2_17_8 : FA_X1 port map( A => ab_17_8_port, B => CARRYB_16_8_port, CI => 
                           SUMB_16_9_port, CO => CARRYB_17_8_port, S => 
                           SUMB_17_8_port);
   S2_17_9 : FA_X1 port map( A => ab_17_9_port, B => CARRYB_16_9_port, CI => 
                           SUMB_16_10_port, CO => CARRYB_17_9_port, S => 
                           SUMB_17_9_port);
   S2_17_10 : FA_X1 port map( A => ab_17_10_port, B => CARRYB_16_10_port, CI =>
                           SUMB_16_11_port, CO => CARRYB_17_10_port, S => 
                           SUMB_17_10_port);
   S2_17_11 : FA_X1 port map( A => ab_17_11_port, B => CARRYB_16_11_port, CI =>
                           SUMB_16_12_port, CO => CARRYB_17_11_port, S => 
                           SUMB_17_11_port);
   S2_17_12 : FA_X1 port map( A => ab_17_12_port, B => CARRYB_16_12_port, CI =>
                           SUMB_16_13_port, CO => CARRYB_17_12_port, S => 
                           SUMB_17_12_port);
   S2_17_13 : FA_X1 port map( A => ab_17_13_port, B => CARRYB_16_13_port, CI =>
                           SUMB_16_14_port, CO => CARRYB_17_13_port, S => 
                           SUMB_17_13_port);
   S2_17_14 : FA_X1 port map( A => ab_17_14_port, B => CARRYB_16_14_port, CI =>
                           SUMB_16_15_port, CO => CARRYB_17_14_port, S => 
                           SUMB_17_14_port);
   S2_17_15 : FA_X1 port map( A => ab_17_15_port, B => CARRYB_16_15_port, CI =>
                           SUMB_16_16_port, CO => CARRYB_17_15_port, S => 
                           SUMB_17_15_port);
   S2_17_16 : FA_X1 port map( A => ab_17_16_port, B => CARRYB_16_16_port, CI =>
                           SUMB_16_17_port, CO => CARRYB_17_16_port, S => 
                           SUMB_17_16_port);
   S2_17_17 : FA_X1 port map( A => ab_17_17_port, B => CARRYB_16_17_port, CI =>
                           SUMB_16_18_port, CO => CARRYB_17_17_port, S => 
                           SUMB_17_17_port);
   S2_17_18 : FA_X1 port map( A => ab_17_18_port, B => CARRYB_16_18_port, CI =>
                           SUMB_16_19_port, CO => CARRYB_17_18_port, S => 
                           SUMB_17_18_port);
   S2_17_19 : FA_X1 port map( A => ab_17_19_port, B => CARRYB_16_19_port, CI =>
                           SUMB_16_20_port, CO => CARRYB_17_19_port, S => 
                           SUMB_17_19_port);
   S2_17_20 : FA_X1 port map( A => ab_17_20_port, B => CARRYB_16_20_port, CI =>
                           SUMB_16_21_port, CO => CARRYB_17_20_port, S => 
                           SUMB_17_20_port);
   S2_17_21 : FA_X1 port map( A => ab_17_21_port, B => CARRYB_16_21_port, CI =>
                           SUMB_16_22_port, CO => CARRYB_17_21_port, S => 
                           SUMB_17_21_port);
   S2_17_22 : FA_X1 port map( A => ab_17_22_port, B => CARRYB_16_22_port, CI =>
                           SUMB_16_23_port, CO => CARRYB_17_22_port, S => 
                           SUMB_17_22_port);
   S2_17_23 : FA_X1 port map( A => ab_17_23_port, B => CARRYB_16_23_port, CI =>
                           SUMB_16_24_port, CO => CARRYB_17_23_port, S => 
                           SUMB_17_23_port);
   S2_17_24 : FA_X1 port map( A => ab_17_24_port, B => CARRYB_16_24_port, CI =>
                           SUMB_16_25_port, CO => CARRYB_17_24_port, S => 
                           SUMB_17_24_port);
   S2_17_25 : FA_X1 port map( A => ab_17_25_port, B => CARRYB_16_25_port, CI =>
                           SUMB_16_26_port, CO => CARRYB_17_25_port, S => 
                           SUMB_17_25_port);
   S2_17_26 : FA_X1 port map( A => ab_17_26_port, B => CARRYB_16_26_port, CI =>
                           SUMB_16_27_port, CO => CARRYB_17_26_port, S => 
                           SUMB_17_26_port);
   S2_17_27 : FA_X1 port map( A => ab_17_27_port, B => CARRYB_16_27_port, CI =>
                           SUMB_16_28_port, CO => CARRYB_17_27_port, S => 
                           SUMB_17_27_port);
   S2_17_28 : FA_X1 port map( A => ab_17_28_port, B => CARRYB_16_28_port, CI =>
                           SUMB_16_29_port, CO => CARRYB_17_28_port, S => 
                           SUMB_17_28_port);
   S2_17_29 : FA_X1 port map( A => ab_17_29_port, B => CARRYB_16_29_port, CI =>
                           SUMB_16_30_port, CO => CARRYB_17_29_port, S => 
                           SUMB_17_29_port);
   S3_17_30 : FA_X1 port map( A => ab_17_30_port, B => CARRYB_16_30_port, CI =>
                           ab_16_31_port, CO => CARRYB_17_30_port, S => 
                           SUMB_17_30_port);
   S1_16_0 : FA_X1 port map( A => ab_16_0_port, B => CARRYB_15_0_port, CI => 
                           SUMB_15_1_port, CO => CARRYB_16_0_port, S => 
                           A1_14_port);
   S2_16_1 : FA_X1 port map( A => ab_16_1_port, B => CARRYB_15_1_port, CI => 
                           SUMB_15_2_port, CO => CARRYB_16_1_port, S => 
                           SUMB_16_1_port);
   S2_16_2 : FA_X1 port map( A => ab_16_2_port, B => CARRYB_15_2_port, CI => 
                           SUMB_15_3_port, CO => CARRYB_16_2_port, S => 
                           SUMB_16_2_port);
   S2_16_3 : FA_X1 port map( A => ab_16_3_port, B => CARRYB_15_3_port, CI => 
                           SUMB_15_4_port, CO => CARRYB_16_3_port, S => 
                           SUMB_16_3_port);
   S2_16_4 : FA_X1 port map( A => ab_16_4_port, B => CARRYB_15_4_port, CI => 
                           SUMB_15_5_port, CO => CARRYB_16_4_port, S => 
                           SUMB_16_4_port);
   S2_16_5 : FA_X1 port map( A => ab_16_5_port, B => CARRYB_15_5_port, CI => 
                           SUMB_15_6_port, CO => CARRYB_16_5_port, S => 
                           SUMB_16_5_port);
   S2_16_6 : FA_X1 port map( A => ab_16_6_port, B => CARRYB_15_6_port, CI => 
                           SUMB_15_7_port, CO => CARRYB_16_6_port, S => 
                           SUMB_16_6_port);
   S2_16_7 : FA_X1 port map( A => ab_16_7_port, B => CARRYB_15_7_port, CI => 
                           SUMB_15_8_port, CO => CARRYB_16_7_port, S => 
                           SUMB_16_7_port);
   S2_16_8 : FA_X1 port map( A => ab_16_8_port, B => CARRYB_15_8_port, CI => 
                           SUMB_15_9_port, CO => CARRYB_16_8_port, S => 
                           SUMB_16_8_port);
   S2_16_9 : FA_X1 port map( A => ab_16_9_port, B => CARRYB_15_9_port, CI => 
                           SUMB_15_10_port, CO => CARRYB_16_9_port, S => 
                           SUMB_16_9_port);
   S2_16_10 : FA_X1 port map( A => ab_16_10_port, B => CARRYB_15_10_port, CI =>
                           SUMB_15_11_port, CO => CARRYB_16_10_port, S => 
                           SUMB_16_10_port);
   S2_16_11 : FA_X1 port map( A => ab_16_11_port, B => CARRYB_15_11_port, CI =>
                           SUMB_15_12_port, CO => CARRYB_16_11_port, S => 
                           SUMB_16_11_port);
   S2_16_12 : FA_X1 port map( A => ab_16_12_port, B => CARRYB_15_12_port, CI =>
                           SUMB_15_13_port, CO => CARRYB_16_12_port, S => 
                           SUMB_16_12_port);
   S2_16_13 : FA_X1 port map( A => ab_16_13_port, B => CARRYB_15_13_port, CI =>
                           SUMB_15_14_port, CO => CARRYB_16_13_port, S => 
                           SUMB_16_13_port);
   S2_16_14 : FA_X1 port map( A => ab_16_14_port, B => CARRYB_15_14_port, CI =>
                           SUMB_15_15_port, CO => CARRYB_16_14_port, S => 
                           SUMB_16_14_port);
   S2_16_15 : FA_X1 port map( A => ab_16_15_port, B => CARRYB_15_15_port, CI =>
                           SUMB_15_16_port, CO => CARRYB_16_15_port, S => 
                           SUMB_16_15_port);
   S2_16_16 : FA_X1 port map( A => ab_16_16_port, B => CARRYB_15_16_port, CI =>
                           SUMB_15_17_port, CO => CARRYB_16_16_port, S => 
                           SUMB_16_16_port);
   S2_16_17 : FA_X1 port map( A => ab_16_17_port, B => CARRYB_15_17_port, CI =>
                           SUMB_15_18_port, CO => CARRYB_16_17_port, S => 
                           SUMB_16_17_port);
   S2_16_18 : FA_X1 port map( A => ab_16_18_port, B => CARRYB_15_18_port, CI =>
                           SUMB_15_19_port, CO => CARRYB_16_18_port, S => 
                           SUMB_16_18_port);
   S2_16_19 : FA_X1 port map( A => ab_16_19_port, B => CARRYB_15_19_port, CI =>
                           SUMB_15_20_port, CO => CARRYB_16_19_port, S => 
                           SUMB_16_19_port);
   S2_16_20 : FA_X1 port map( A => ab_16_20_port, B => CARRYB_15_20_port, CI =>
                           SUMB_15_21_port, CO => CARRYB_16_20_port, S => 
                           SUMB_16_20_port);
   S2_16_21 : FA_X1 port map( A => ab_16_21_port, B => CARRYB_15_21_port, CI =>
                           SUMB_15_22_port, CO => CARRYB_16_21_port, S => 
                           SUMB_16_21_port);
   S2_16_22 : FA_X1 port map( A => ab_16_22_port, B => CARRYB_15_22_port, CI =>
                           SUMB_15_23_port, CO => CARRYB_16_22_port, S => 
                           SUMB_16_22_port);
   S2_16_23 : FA_X1 port map( A => ab_16_23_port, B => CARRYB_15_23_port, CI =>
                           SUMB_15_24_port, CO => CARRYB_16_23_port, S => 
                           SUMB_16_23_port);
   S2_16_24 : FA_X1 port map( A => ab_16_24_port, B => CARRYB_15_24_port, CI =>
                           SUMB_15_25_port, CO => CARRYB_16_24_port, S => 
                           SUMB_16_24_port);
   S2_16_25 : FA_X1 port map( A => ab_16_25_port, B => CARRYB_15_25_port, CI =>
                           SUMB_15_26_port, CO => CARRYB_16_25_port, S => 
                           SUMB_16_25_port);
   S2_16_26 : FA_X1 port map( A => ab_16_26_port, B => CARRYB_15_26_port, CI =>
                           SUMB_15_27_port, CO => CARRYB_16_26_port, S => 
                           SUMB_16_26_port);
   S2_16_27 : FA_X1 port map( A => ab_16_27_port, B => CARRYB_15_27_port, CI =>
                           SUMB_15_28_port, CO => CARRYB_16_27_port, S => 
                           SUMB_16_27_port);
   S2_16_28 : FA_X1 port map( A => ab_16_28_port, B => CARRYB_15_28_port, CI =>
                           SUMB_15_29_port, CO => CARRYB_16_28_port, S => 
                           SUMB_16_28_port);
   S2_16_29 : FA_X1 port map( A => ab_16_29_port, B => CARRYB_15_29_port, CI =>
                           SUMB_15_30_port, CO => CARRYB_16_29_port, S => 
                           SUMB_16_29_port);
   S3_16_30 : FA_X1 port map( A => ab_16_30_port, B => CARRYB_15_30_port, CI =>
                           ab_15_31_port, CO => CARRYB_16_30_port, S => 
                           SUMB_16_30_port);
   S1_15_0 : FA_X1 port map( A => ab_15_0_port, B => CARRYB_14_0_port, CI => 
                           SUMB_14_1_port, CO => CARRYB_15_0_port, S => 
                           A1_13_port);
   S2_15_1 : FA_X1 port map( A => ab_15_1_port, B => CARRYB_14_1_port, CI => 
                           SUMB_14_2_port, CO => CARRYB_15_1_port, S => 
                           SUMB_15_1_port);
   S2_15_2 : FA_X1 port map( A => ab_15_2_port, B => CARRYB_14_2_port, CI => 
                           SUMB_14_3_port, CO => CARRYB_15_2_port, S => 
                           SUMB_15_2_port);
   S2_15_3 : FA_X1 port map( A => ab_15_3_port, B => CARRYB_14_3_port, CI => 
                           SUMB_14_4_port, CO => CARRYB_15_3_port, S => 
                           SUMB_15_3_port);
   S2_15_4 : FA_X1 port map( A => ab_15_4_port, B => CARRYB_14_4_port, CI => 
                           SUMB_14_5_port, CO => CARRYB_15_4_port, S => 
                           SUMB_15_4_port);
   S2_15_5 : FA_X1 port map( A => ab_15_5_port, B => CARRYB_14_5_port, CI => 
                           SUMB_14_6_port, CO => CARRYB_15_5_port, S => 
                           SUMB_15_5_port);
   S2_15_6 : FA_X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, CI => 
                           SUMB_14_7_port, CO => CARRYB_15_6_port, S => 
                           SUMB_15_6_port);
   S2_15_7 : FA_X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, CI => 
                           SUMB_14_8_port, CO => CARRYB_15_7_port, S => 
                           SUMB_15_7_port);
   S2_15_8 : FA_X1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, CI => 
                           SUMB_14_9_port, CO => CARRYB_15_8_port, S => 
                           SUMB_15_8_port);
   S2_15_9 : FA_X1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, CI => 
                           SUMB_14_10_port, CO => CARRYB_15_9_port, S => 
                           SUMB_15_9_port);
   S2_15_10 : FA_X1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, CI =>
                           SUMB_14_11_port, CO => CARRYB_15_10_port, S => 
                           SUMB_15_10_port);
   S2_15_11 : FA_X1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, CI =>
                           SUMB_14_12_port, CO => CARRYB_15_11_port, S => 
                           SUMB_15_11_port);
   S2_15_12 : FA_X1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, CI =>
                           SUMB_14_13_port, CO => CARRYB_15_12_port, S => 
                           SUMB_15_12_port);
   S2_15_13 : FA_X1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, CI =>
                           SUMB_14_14_port, CO => CARRYB_15_13_port, S => 
                           SUMB_15_13_port);
   S2_15_14 : FA_X1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, CI =>
                           SUMB_14_15_port, CO => CARRYB_15_14_port, S => 
                           SUMB_15_14_port);
   S2_15_15 : FA_X1 port map( A => ab_15_15_port, B => CARRYB_14_15_port, CI =>
                           SUMB_14_16_port, CO => CARRYB_15_15_port, S => 
                           SUMB_15_15_port);
   S2_15_16 : FA_X1 port map( A => ab_15_16_port, B => CARRYB_14_16_port, CI =>
                           SUMB_14_17_port, CO => CARRYB_15_16_port, S => 
                           SUMB_15_16_port);
   S2_15_17 : FA_X1 port map( A => ab_15_17_port, B => CARRYB_14_17_port, CI =>
                           SUMB_14_18_port, CO => CARRYB_15_17_port, S => 
                           SUMB_15_17_port);
   S2_15_18 : FA_X1 port map( A => ab_15_18_port, B => CARRYB_14_18_port, CI =>
                           SUMB_14_19_port, CO => CARRYB_15_18_port, S => 
                           SUMB_15_18_port);
   S2_15_19 : FA_X1 port map( A => ab_15_19_port, B => CARRYB_14_19_port, CI =>
                           SUMB_14_20_port, CO => CARRYB_15_19_port, S => 
                           SUMB_15_19_port);
   S2_15_20 : FA_X1 port map( A => ab_15_20_port, B => CARRYB_14_20_port, CI =>
                           SUMB_14_21_port, CO => CARRYB_15_20_port, S => 
                           SUMB_15_20_port);
   S2_15_21 : FA_X1 port map( A => ab_15_21_port, B => CARRYB_14_21_port, CI =>
                           SUMB_14_22_port, CO => CARRYB_15_21_port, S => 
                           SUMB_15_21_port);
   S2_15_22 : FA_X1 port map( A => ab_15_22_port, B => CARRYB_14_22_port, CI =>
                           SUMB_14_23_port, CO => CARRYB_15_22_port, S => 
                           SUMB_15_22_port);
   S2_15_23 : FA_X1 port map( A => ab_15_23_port, B => CARRYB_14_23_port, CI =>
                           SUMB_14_24_port, CO => CARRYB_15_23_port, S => 
                           SUMB_15_23_port);
   S2_15_24 : FA_X1 port map( A => ab_15_24_port, B => CARRYB_14_24_port, CI =>
                           SUMB_14_25_port, CO => CARRYB_15_24_port, S => 
                           SUMB_15_24_port);
   S2_15_25 : FA_X1 port map( A => ab_15_25_port, B => CARRYB_14_25_port, CI =>
                           SUMB_14_26_port, CO => CARRYB_15_25_port, S => 
                           SUMB_15_25_port);
   S2_15_26 : FA_X1 port map( A => ab_15_26_port, B => CARRYB_14_26_port, CI =>
                           SUMB_14_27_port, CO => CARRYB_15_26_port, S => 
                           SUMB_15_26_port);
   S2_15_27 : FA_X1 port map( A => ab_15_27_port, B => CARRYB_14_27_port, CI =>
                           SUMB_14_28_port, CO => CARRYB_15_27_port, S => 
                           SUMB_15_27_port);
   S2_15_28 : FA_X1 port map( A => ab_15_28_port, B => CARRYB_14_28_port, CI =>
                           SUMB_14_29_port, CO => CARRYB_15_28_port, S => 
                           SUMB_15_28_port);
   S2_15_29 : FA_X1 port map( A => ab_15_29_port, B => CARRYB_14_29_port, CI =>
                           SUMB_14_30_port, CO => CARRYB_15_29_port, S => 
                           SUMB_15_29_port);
   S3_15_30 : FA_X1 port map( A => ab_15_30_port, B => CARRYB_14_30_port, CI =>
                           ab_14_31_port, CO => CARRYB_15_30_port, S => 
                           SUMB_15_30_port);
   S1_14_0 : FA_X1 port map( A => ab_14_0_port, B => CARRYB_13_0_port, CI => 
                           SUMB_13_1_port, CO => CARRYB_14_0_port, S => 
                           A1_12_port);
   S2_14_1 : FA_X1 port map( A => ab_14_1_port, B => CARRYB_13_1_port, CI => 
                           SUMB_13_2_port, CO => CARRYB_14_1_port, S => 
                           SUMB_14_1_port);
   S2_14_2 : FA_X1 port map( A => ab_14_2_port, B => CARRYB_13_2_port, CI => 
                           SUMB_13_3_port, CO => CARRYB_14_2_port, S => 
                           SUMB_14_2_port);
   S2_14_3 : FA_X1 port map( A => ab_14_3_port, B => CARRYB_13_3_port, CI => 
                           SUMB_13_4_port, CO => CARRYB_14_3_port, S => 
                           SUMB_14_3_port);
   S2_14_4 : FA_X1 port map( A => ab_14_4_port, B => CARRYB_13_4_port, CI => 
                           SUMB_13_5_port, CO => CARRYB_14_4_port, S => 
                           SUMB_14_4_port);
   S2_14_5 : FA_X1 port map( A => ab_14_5_port, B => CARRYB_13_5_port, CI => 
                           SUMB_13_6_port, CO => CARRYB_14_5_port, S => 
                           SUMB_14_5_port);
   S2_14_6 : FA_X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, CI => 
                           SUMB_13_7_port, CO => CARRYB_14_6_port, S => 
                           SUMB_14_6_port);
   S2_14_7 : FA_X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, CI => 
                           SUMB_13_8_port, CO => CARRYB_14_7_port, S => 
                           SUMB_14_7_port);
   S2_14_8 : FA_X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, CI => 
                           SUMB_13_9_port, CO => CARRYB_14_8_port, S => 
                           SUMB_14_8_port);
   S2_14_9 : FA_X1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, CI => 
                           SUMB_13_10_port, CO => CARRYB_14_9_port, S => 
                           SUMB_14_9_port);
   S2_14_10 : FA_X1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, CI =>
                           SUMB_13_11_port, CO => CARRYB_14_10_port, S => 
                           SUMB_14_10_port);
   S2_14_11 : FA_X1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, CI =>
                           SUMB_13_12_port, CO => CARRYB_14_11_port, S => 
                           SUMB_14_11_port);
   S2_14_12 : FA_X1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, CI =>
                           SUMB_13_13_port, CO => CARRYB_14_12_port, S => 
                           SUMB_14_12_port);
   S2_14_13 : FA_X1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, CI =>
                           SUMB_13_14_port, CO => CARRYB_14_13_port, S => 
                           SUMB_14_13_port);
   S2_14_14 : FA_X1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, CI =>
                           SUMB_13_15_port, CO => CARRYB_14_14_port, S => 
                           SUMB_14_14_port);
   S2_14_15 : FA_X1 port map( A => ab_14_15_port, B => CARRYB_13_15_port, CI =>
                           SUMB_13_16_port, CO => CARRYB_14_15_port, S => 
                           SUMB_14_15_port);
   S2_14_16 : FA_X1 port map( A => ab_14_16_port, B => CARRYB_13_16_port, CI =>
                           SUMB_13_17_port, CO => CARRYB_14_16_port, S => 
                           SUMB_14_16_port);
   S2_14_17 : FA_X1 port map( A => ab_14_17_port, B => CARRYB_13_17_port, CI =>
                           SUMB_13_18_port, CO => CARRYB_14_17_port, S => 
                           SUMB_14_17_port);
   S2_14_18 : FA_X1 port map( A => ab_14_18_port, B => CARRYB_13_18_port, CI =>
                           SUMB_13_19_port, CO => CARRYB_14_18_port, S => 
                           SUMB_14_18_port);
   S2_14_19 : FA_X1 port map( A => ab_14_19_port, B => CARRYB_13_19_port, CI =>
                           SUMB_13_20_port, CO => CARRYB_14_19_port, S => 
                           SUMB_14_19_port);
   S2_14_20 : FA_X1 port map( A => ab_14_20_port, B => CARRYB_13_20_port, CI =>
                           SUMB_13_21_port, CO => CARRYB_14_20_port, S => 
                           SUMB_14_20_port);
   S2_14_21 : FA_X1 port map( A => ab_14_21_port, B => CARRYB_13_21_port, CI =>
                           SUMB_13_22_port, CO => CARRYB_14_21_port, S => 
                           SUMB_14_21_port);
   S2_14_22 : FA_X1 port map( A => ab_14_22_port, B => CARRYB_13_22_port, CI =>
                           SUMB_13_23_port, CO => CARRYB_14_22_port, S => 
                           SUMB_14_22_port);
   S2_14_23 : FA_X1 port map( A => ab_14_23_port, B => CARRYB_13_23_port, CI =>
                           SUMB_13_24_port, CO => CARRYB_14_23_port, S => 
                           SUMB_14_23_port);
   S2_14_24 : FA_X1 port map( A => ab_14_24_port, B => CARRYB_13_24_port, CI =>
                           SUMB_13_25_port, CO => CARRYB_14_24_port, S => 
                           SUMB_14_24_port);
   S2_14_25 : FA_X1 port map( A => ab_14_25_port, B => CARRYB_13_25_port, CI =>
                           SUMB_13_26_port, CO => CARRYB_14_25_port, S => 
                           SUMB_14_25_port);
   S2_14_26 : FA_X1 port map( A => ab_14_26_port, B => CARRYB_13_26_port, CI =>
                           SUMB_13_27_port, CO => CARRYB_14_26_port, S => 
                           SUMB_14_26_port);
   S2_14_27 : FA_X1 port map( A => ab_14_27_port, B => CARRYB_13_27_port, CI =>
                           SUMB_13_28_port, CO => CARRYB_14_27_port, S => 
                           SUMB_14_27_port);
   S2_14_28 : FA_X1 port map( A => ab_14_28_port, B => CARRYB_13_28_port, CI =>
                           SUMB_13_29_port, CO => CARRYB_14_28_port, S => 
                           SUMB_14_28_port);
   S2_14_29 : FA_X1 port map( A => ab_14_29_port, B => CARRYB_13_29_port, CI =>
                           SUMB_13_30_port, CO => CARRYB_14_29_port, S => 
                           SUMB_14_29_port);
   S3_14_30 : FA_X1 port map( A => ab_14_30_port, B => CARRYB_13_30_port, CI =>
                           ab_13_31_port, CO => CARRYB_14_30_port, S => 
                           SUMB_14_30_port);
   S1_13_0 : FA_X1 port map( A => ab_13_0_port, B => CARRYB_12_0_port, CI => 
                           SUMB_12_1_port, CO => CARRYB_13_0_port, S => 
                           A1_11_port);
   S2_13_1 : FA_X1 port map( A => ab_13_1_port, B => CARRYB_12_1_port, CI => 
                           SUMB_12_2_port, CO => CARRYB_13_1_port, S => 
                           SUMB_13_1_port);
   S2_13_2 : FA_X1 port map( A => ab_13_2_port, B => CARRYB_12_2_port, CI => 
                           SUMB_12_3_port, CO => CARRYB_13_2_port, S => 
                           SUMB_13_2_port);
   S2_13_3 : FA_X1 port map( A => ab_13_3_port, B => CARRYB_12_3_port, CI => 
                           SUMB_12_4_port, CO => CARRYB_13_3_port, S => 
                           SUMB_13_3_port);
   S2_13_4 : FA_X1 port map( A => ab_13_4_port, B => CARRYB_12_4_port, CI => 
                           SUMB_12_5_port, CO => CARRYB_13_4_port, S => 
                           SUMB_13_4_port);
   S2_13_5 : FA_X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, CI => 
                           SUMB_12_6_port, CO => CARRYB_13_5_port, S => 
                           SUMB_13_5_port);
   S2_13_6 : FA_X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, CI => 
                           SUMB_12_7_port, CO => CARRYB_13_6_port, S => 
                           SUMB_13_6_port);
   S2_13_7 : FA_X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, CI => 
                           SUMB_12_8_port, CO => CARRYB_13_7_port, S => 
                           SUMB_13_7_port);
   S2_13_8 : FA_X1 port map( A => ab_13_8_port, B => CARRYB_12_8_port, CI => 
                           SUMB_12_9_port, CO => CARRYB_13_8_port, S => 
                           SUMB_13_8_port);
   S2_13_9 : FA_X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, CI => 
                           SUMB_12_10_port, CO => CARRYB_13_9_port, S => 
                           SUMB_13_9_port);
   S2_13_10 : FA_X1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, CI =>
                           SUMB_12_11_port, CO => CARRYB_13_10_port, S => 
                           SUMB_13_10_port);
   S2_13_11 : FA_X1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, CI =>
                           SUMB_12_12_port, CO => CARRYB_13_11_port, S => 
                           SUMB_13_11_port);
   S2_13_12 : FA_X1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, CI =>
                           SUMB_12_13_port, CO => CARRYB_13_12_port, S => 
                           SUMB_13_12_port);
   S2_13_13 : FA_X1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, CI =>
                           SUMB_12_14_port, CO => CARRYB_13_13_port, S => 
                           SUMB_13_13_port);
   S2_13_14 : FA_X1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, CI =>
                           SUMB_12_15_port, CO => CARRYB_13_14_port, S => 
                           SUMB_13_14_port);
   S2_13_15 : FA_X1 port map( A => ab_13_15_port, B => CARRYB_12_15_port, CI =>
                           SUMB_12_16_port, CO => CARRYB_13_15_port, S => 
                           SUMB_13_15_port);
   S2_13_16 : FA_X1 port map( A => ab_13_16_port, B => CARRYB_12_16_port, CI =>
                           SUMB_12_17_port, CO => CARRYB_13_16_port, S => 
                           SUMB_13_16_port);
   S2_13_17 : FA_X1 port map( A => ab_13_17_port, B => CARRYB_12_17_port, CI =>
                           SUMB_12_18_port, CO => CARRYB_13_17_port, S => 
                           SUMB_13_17_port);
   S2_13_18 : FA_X1 port map( A => ab_13_18_port, B => CARRYB_12_18_port, CI =>
                           SUMB_12_19_port, CO => CARRYB_13_18_port, S => 
                           SUMB_13_18_port);
   S2_13_19 : FA_X1 port map( A => ab_13_19_port, B => CARRYB_12_19_port, CI =>
                           SUMB_12_20_port, CO => CARRYB_13_19_port, S => 
                           SUMB_13_19_port);
   S2_13_20 : FA_X1 port map( A => ab_13_20_port, B => CARRYB_12_20_port, CI =>
                           SUMB_12_21_port, CO => CARRYB_13_20_port, S => 
                           SUMB_13_20_port);
   S2_13_21 : FA_X1 port map( A => ab_13_21_port, B => CARRYB_12_21_port, CI =>
                           SUMB_12_22_port, CO => CARRYB_13_21_port, S => 
                           SUMB_13_21_port);
   S2_13_22 : FA_X1 port map( A => ab_13_22_port, B => CARRYB_12_22_port, CI =>
                           SUMB_12_23_port, CO => CARRYB_13_22_port, S => 
                           SUMB_13_22_port);
   S2_13_23 : FA_X1 port map( A => ab_13_23_port, B => CARRYB_12_23_port, CI =>
                           SUMB_12_24_port, CO => CARRYB_13_23_port, S => 
                           SUMB_13_23_port);
   S2_13_24 : FA_X1 port map( A => ab_13_24_port, B => CARRYB_12_24_port, CI =>
                           SUMB_12_25_port, CO => CARRYB_13_24_port, S => 
                           SUMB_13_24_port);
   S2_13_25 : FA_X1 port map( A => ab_13_25_port, B => CARRYB_12_25_port, CI =>
                           SUMB_12_26_port, CO => CARRYB_13_25_port, S => 
                           SUMB_13_25_port);
   S2_13_26 : FA_X1 port map( A => ab_13_26_port, B => CARRYB_12_26_port, CI =>
                           SUMB_12_27_port, CO => CARRYB_13_26_port, S => 
                           SUMB_13_26_port);
   S2_13_27 : FA_X1 port map( A => ab_13_27_port, B => CARRYB_12_27_port, CI =>
                           SUMB_12_28_port, CO => CARRYB_13_27_port, S => 
                           SUMB_13_27_port);
   S2_13_28 : FA_X1 port map( A => ab_13_28_port, B => CARRYB_12_28_port, CI =>
                           SUMB_12_29_port, CO => CARRYB_13_28_port, S => 
                           SUMB_13_28_port);
   S2_13_29 : FA_X1 port map( A => ab_13_29_port, B => CARRYB_12_29_port, CI =>
                           SUMB_12_30_port, CO => CARRYB_13_29_port, S => 
                           SUMB_13_29_port);
   S3_13_30 : FA_X1 port map( A => ab_13_30_port, B => CARRYB_12_30_port, CI =>
                           ab_12_31_port, CO => CARRYB_13_30_port, S => 
                           SUMB_13_30_port);
   S1_12_0 : FA_X1 port map( A => ab_12_0_port, B => CARRYB_11_0_port, CI => 
                           SUMB_11_1_port, CO => CARRYB_12_0_port, S => 
                           A1_10_port);
   S2_12_1 : FA_X1 port map( A => ab_12_1_port, B => CARRYB_11_1_port, CI => 
                           SUMB_11_2_port, CO => CARRYB_12_1_port, S => 
                           SUMB_12_1_port);
   S2_12_2 : FA_X1 port map( A => ab_12_2_port, B => CARRYB_11_2_port, CI => 
                           SUMB_11_3_port, CO => CARRYB_12_2_port, S => 
                           SUMB_12_2_port);
   S2_12_3 : FA_X1 port map( A => ab_12_3_port, B => CARRYB_11_3_port, CI => 
                           SUMB_11_4_port, CO => CARRYB_12_3_port, S => 
                           SUMB_12_3_port);
   S2_12_4 : FA_X1 port map( A => ab_12_4_port, B => CARRYB_11_4_port, CI => 
                           SUMB_11_5_port, CO => CARRYB_12_4_port, S => 
                           SUMB_12_4_port);
   S2_12_5 : FA_X1 port map( A => ab_12_5_port, B => CARRYB_11_5_port, CI => 
                           SUMB_11_6_port, CO => CARRYB_12_5_port, S => 
                           SUMB_12_5_port);
   S2_12_6 : FA_X1 port map( A => ab_12_6_port, B => CARRYB_11_6_port, CI => 
                           SUMB_11_7_port, CO => CARRYB_12_6_port, S => 
                           SUMB_12_6_port);
   S2_12_7 : FA_X1 port map( A => ab_12_7_port, B => CARRYB_11_7_port, CI => 
                           SUMB_11_8_port, CO => CARRYB_12_7_port, S => 
                           SUMB_12_7_port);
   S2_12_8 : FA_X1 port map( A => ab_12_8_port, B => CARRYB_11_8_port, CI => 
                           SUMB_11_9_port, CO => CARRYB_12_8_port, S => 
                           SUMB_12_8_port);
   S2_12_9 : FA_X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, CI => 
                           SUMB_11_10_port, CO => CARRYB_12_9_port, S => 
                           SUMB_12_9_port);
   S2_12_10 : FA_X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, CI =>
                           SUMB_11_11_port, CO => CARRYB_12_10_port, S => 
                           SUMB_12_10_port);
   S2_12_11 : FA_X1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, CI =>
                           SUMB_11_12_port, CO => CARRYB_12_11_port, S => 
                           SUMB_12_11_port);
   S2_12_12 : FA_X1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, CI =>
                           SUMB_11_13_port, CO => CARRYB_12_12_port, S => 
                           SUMB_12_12_port);
   S2_12_13 : FA_X1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, CI =>
                           SUMB_11_14_port, CO => CARRYB_12_13_port, S => 
                           SUMB_12_13_port);
   S2_12_14 : FA_X1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, CI =>
                           SUMB_11_15_port, CO => CARRYB_12_14_port, S => 
                           SUMB_12_14_port);
   S2_12_15 : FA_X1 port map( A => ab_12_15_port, B => CARRYB_11_15_port, CI =>
                           SUMB_11_16_port, CO => CARRYB_12_15_port, S => 
                           SUMB_12_15_port);
   S2_12_16 : FA_X1 port map( A => ab_12_16_port, B => CARRYB_11_16_port, CI =>
                           SUMB_11_17_port, CO => CARRYB_12_16_port, S => 
                           SUMB_12_16_port);
   S2_12_17 : FA_X1 port map( A => ab_12_17_port, B => CARRYB_11_17_port, CI =>
                           SUMB_11_18_port, CO => CARRYB_12_17_port, S => 
                           SUMB_12_17_port);
   S2_12_18 : FA_X1 port map( A => ab_12_18_port, B => CARRYB_11_18_port, CI =>
                           SUMB_11_19_port, CO => CARRYB_12_18_port, S => 
                           SUMB_12_18_port);
   S2_12_19 : FA_X1 port map( A => ab_12_19_port, B => CARRYB_11_19_port, CI =>
                           SUMB_11_20_port, CO => CARRYB_12_19_port, S => 
                           SUMB_12_19_port);
   S2_12_20 : FA_X1 port map( A => ab_12_20_port, B => CARRYB_11_20_port, CI =>
                           SUMB_11_21_port, CO => CARRYB_12_20_port, S => 
                           SUMB_12_20_port);
   S2_12_21 : FA_X1 port map( A => ab_12_21_port, B => CARRYB_11_21_port, CI =>
                           SUMB_11_22_port, CO => CARRYB_12_21_port, S => 
                           SUMB_12_21_port);
   S2_12_22 : FA_X1 port map( A => ab_12_22_port, B => CARRYB_11_22_port, CI =>
                           SUMB_11_23_port, CO => CARRYB_12_22_port, S => 
                           SUMB_12_22_port);
   S2_12_23 : FA_X1 port map( A => ab_12_23_port, B => CARRYB_11_23_port, CI =>
                           SUMB_11_24_port, CO => CARRYB_12_23_port, S => 
                           SUMB_12_23_port);
   S2_12_24 : FA_X1 port map( A => ab_12_24_port, B => CARRYB_11_24_port, CI =>
                           SUMB_11_25_port, CO => CARRYB_12_24_port, S => 
                           SUMB_12_24_port);
   S2_12_25 : FA_X1 port map( A => ab_12_25_port, B => CARRYB_11_25_port, CI =>
                           SUMB_11_26_port, CO => CARRYB_12_25_port, S => 
                           SUMB_12_25_port);
   S2_12_26 : FA_X1 port map( A => ab_12_26_port, B => CARRYB_11_26_port, CI =>
                           SUMB_11_27_port, CO => CARRYB_12_26_port, S => 
                           SUMB_12_26_port);
   S2_12_27 : FA_X1 port map( A => ab_12_27_port, B => CARRYB_11_27_port, CI =>
                           SUMB_11_28_port, CO => CARRYB_12_27_port, S => 
                           SUMB_12_27_port);
   S2_12_28 : FA_X1 port map( A => ab_12_28_port, B => CARRYB_11_28_port, CI =>
                           SUMB_11_29_port, CO => CARRYB_12_28_port, S => 
                           SUMB_12_28_port);
   S2_12_29 : FA_X1 port map( A => ab_12_29_port, B => CARRYB_11_29_port, CI =>
                           SUMB_11_30_port, CO => CARRYB_12_29_port, S => 
                           SUMB_12_29_port);
   S3_12_30 : FA_X1 port map( A => ab_12_30_port, B => CARRYB_11_30_port, CI =>
                           ab_11_31_port, CO => CARRYB_12_30_port, S => 
                           SUMB_12_30_port);
   S1_11_0 : FA_X1 port map( A => ab_11_0_port, B => CARRYB_10_0_port, CI => 
                           SUMB_10_1_port, CO => CARRYB_11_0_port, S => 
                           A1_9_port);
   S2_11_1 : FA_X1 port map( A => ab_11_1_port, B => CARRYB_10_1_port, CI => 
                           SUMB_10_2_port, CO => CARRYB_11_1_port, S => 
                           SUMB_11_1_port);
   S2_11_2 : FA_X1 port map( A => ab_11_2_port, B => CARRYB_10_2_port, CI => 
                           SUMB_10_3_port, CO => CARRYB_11_2_port, S => 
                           SUMB_11_2_port);
   S2_11_3 : FA_X1 port map( A => ab_11_3_port, B => CARRYB_10_3_port, CI => 
                           SUMB_10_4_port, CO => CARRYB_11_3_port, S => 
                           SUMB_11_3_port);
   S2_11_4 : FA_X1 port map( A => ab_11_4_port, B => CARRYB_10_4_port, CI => 
                           SUMB_10_5_port, CO => CARRYB_11_4_port, S => 
                           SUMB_11_4_port);
   S2_11_5 : FA_X1 port map( A => ab_11_5_port, B => CARRYB_10_5_port, CI => 
                           SUMB_10_6_port, CO => CARRYB_11_5_port, S => 
                           SUMB_11_5_port);
   S2_11_6 : FA_X1 port map( A => ab_11_6_port, B => CARRYB_10_6_port, CI => 
                           SUMB_10_7_port, CO => CARRYB_11_6_port, S => 
                           SUMB_11_6_port);
   S2_11_7 : FA_X1 port map( A => ab_11_7_port, B => CARRYB_10_7_port, CI => 
                           SUMB_10_8_port, CO => CARRYB_11_7_port, S => 
                           SUMB_11_7_port);
   S2_11_8 : FA_X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, CI => 
                           SUMB_10_9_port, CO => CARRYB_11_8_port, S => 
                           SUMB_11_8_port);
   S2_11_9 : FA_X1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, CI => 
                           SUMB_10_10_port, CO => CARRYB_11_9_port, S => 
                           SUMB_11_9_port);
   S2_11_10 : FA_X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, CI =>
                           SUMB_10_11_port, CO => CARRYB_11_10_port, S => 
                           SUMB_11_10_port);
   S2_11_11 : FA_X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, CI =>
                           SUMB_10_12_port, CO => CARRYB_11_11_port, S => 
                           SUMB_11_11_port);
   S2_11_12 : FA_X1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, CI =>
                           SUMB_10_13_port, CO => CARRYB_11_12_port, S => 
                           SUMB_11_12_port);
   S2_11_13 : FA_X1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, CI =>
                           SUMB_10_14_port, CO => CARRYB_11_13_port, S => 
                           SUMB_11_13_port);
   S2_11_14 : FA_X1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, CI =>
                           SUMB_10_15_port, CO => CARRYB_11_14_port, S => 
                           SUMB_11_14_port);
   S2_11_15 : FA_X1 port map( A => ab_11_15_port, B => CARRYB_10_15_port, CI =>
                           SUMB_10_16_port, CO => CARRYB_11_15_port, S => 
                           SUMB_11_15_port);
   S2_11_16 : FA_X1 port map( A => ab_11_16_port, B => CARRYB_10_16_port, CI =>
                           SUMB_10_17_port, CO => CARRYB_11_16_port, S => 
                           SUMB_11_16_port);
   S2_11_17 : FA_X1 port map( A => ab_11_17_port, B => CARRYB_10_17_port, CI =>
                           SUMB_10_18_port, CO => CARRYB_11_17_port, S => 
                           SUMB_11_17_port);
   S2_11_18 : FA_X1 port map( A => ab_11_18_port, B => CARRYB_10_18_port, CI =>
                           SUMB_10_19_port, CO => CARRYB_11_18_port, S => 
                           SUMB_11_18_port);
   S2_11_19 : FA_X1 port map( A => ab_11_19_port, B => CARRYB_10_19_port, CI =>
                           SUMB_10_20_port, CO => CARRYB_11_19_port, S => 
                           SUMB_11_19_port);
   S2_11_20 : FA_X1 port map( A => ab_11_20_port, B => CARRYB_10_20_port, CI =>
                           SUMB_10_21_port, CO => CARRYB_11_20_port, S => 
                           SUMB_11_20_port);
   S2_11_21 : FA_X1 port map( A => ab_11_21_port, B => CARRYB_10_21_port, CI =>
                           SUMB_10_22_port, CO => CARRYB_11_21_port, S => 
                           SUMB_11_21_port);
   S2_11_22 : FA_X1 port map( A => ab_11_22_port, B => CARRYB_10_22_port, CI =>
                           SUMB_10_23_port, CO => CARRYB_11_22_port, S => 
                           SUMB_11_22_port);
   S2_11_23 : FA_X1 port map( A => ab_11_23_port, B => CARRYB_10_23_port, CI =>
                           SUMB_10_24_port, CO => CARRYB_11_23_port, S => 
                           SUMB_11_23_port);
   S2_11_24 : FA_X1 port map( A => ab_11_24_port, B => CARRYB_10_24_port, CI =>
                           SUMB_10_25_port, CO => CARRYB_11_24_port, S => 
                           SUMB_11_24_port);
   S2_11_25 : FA_X1 port map( A => ab_11_25_port, B => CARRYB_10_25_port, CI =>
                           SUMB_10_26_port, CO => CARRYB_11_25_port, S => 
                           SUMB_11_25_port);
   S2_11_26 : FA_X1 port map( A => ab_11_26_port, B => CARRYB_10_26_port, CI =>
                           SUMB_10_27_port, CO => CARRYB_11_26_port, S => 
                           SUMB_11_26_port);
   S2_11_27 : FA_X1 port map( A => ab_11_27_port, B => CARRYB_10_27_port, CI =>
                           SUMB_10_28_port, CO => CARRYB_11_27_port, S => 
                           SUMB_11_27_port);
   S2_11_28 : FA_X1 port map( A => ab_11_28_port, B => CARRYB_10_28_port, CI =>
                           SUMB_10_29_port, CO => CARRYB_11_28_port, S => 
                           SUMB_11_28_port);
   S2_11_29 : FA_X1 port map( A => ab_11_29_port, B => CARRYB_10_29_port, CI =>
                           SUMB_10_30_port, CO => CARRYB_11_29_port, S => 
                           SUMB_11_29_port);
   S3_11_30 : FA_X1 port map( A => ab_11_30_port, B => CARRYB_10_30_port, CI =>
                           ab_10_31_port, CO => CARRYB_11_30_port, S => 
                           SUMB_11_30_port);
   S1_10_0 : FA_X1 port map( A => ab_10_0_port, B => CARRYB_9_0_port, CI => 
                           SUMB_9_1_port, CO => CARRYB_10_0_port, S => 
                           A1_8_port);
   S2_10_1 : FA_X1 port map( A => ab_10_1_port, B => CARRYB_9_1_port, CI => 
                           SUMB_9_2_port, CO => CARRYB_10_1_port, S => 
                           SUMB_10_1_port);
   S2_10_2 : FA_X1 port map( A => ab_10_2_port, B => CARRYB_9_2_port, CI => 
                           SUMB_9_3_port, CO => CARRYB_10_2_port, S => 
                           SUMB_10_2_port);
   S2_10_3 : FA_X1 port map( A => ab_10_3_port, B => CARRYB_9_3_port, CI => 
                           SUMB_9_4_port, CO => CARRYB_10_3_port, S => 
                           SUMB_10_3_port);
   S2_10_4 : FA_X1 port map( A => ab_10_4_port, B => CARRYB_9_4_port, CI => 
                           SUMB_9_5_port, CO => CARRYB_10_4_port, S => 
                           SUMB_10_4_port);
   S2_10_5 : FA_X1 port map( A => ab_10_5_port, B => CARRYB_9_5_port, CI => 
                           SUMB_9_6_port, CO => CARRYB_10_5_port, S => 
                           SUMB_10_5_port);
   S2_10_6 : FA_X1 port map( A => ab_10_6_port, B => CARRYB_9_6_port, CI => 
                           SUMB_9_7_port, CO => CARRYB_10_6_port, S => 
                           SUMB_10_6_port);
   S2_10_7 : FA_X1 port map( A => ab_10_7_port, B => CARRYB_9_7_port, CI => 
                           SUMB_9_8_port, CO => CARRYB_10_7_port, S => 
                           SUMB_10_7_port);
   S2_10_8 : FA_X1 port map( A => ab_10_8_port, B => CARRYB_9_8_port, CI => 
                           SUMB_9_9_port, CO => CARRYB_10_8_port, S => 
                           SUMB_10_8_port);
   S2_10_9 : FA_X1 port map( A => ab_10_9_port, B => CARRYB_9_9_port, CI => 
                           SUMB_9_10_port, CO => CARRYB_10_9_port, S => 
                           SUMB_10_9_port);
   S2_10_10 : FA_X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, CI => 
                           SUMB_9_11_port, CO => CARRYB_10_10_port, S => 
                           SUMB_10_10_port);
   S2_10_11 : FA_X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, CI => 
                           SUMB_9_12_port, CO => CARRYB_10_11_port, S => 
                           SUMB_10_11_port);
   S2_10_12 : FA_X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, CI => 
                           SUMB_9_13_port, CO => CARRYB_10_12_port, S => 
                           SUMB_10_12_port);
   S2_10_13 : FA_X1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, CI => 
                           SUMB_9_14_port, CO => CARRYB_10_13_port, S => 
                           SUMB_10_13_port);
   S2_10_14 : FA_X1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, CI => 
                           SUMB_9_15_port, CO => CARRYB_10_14_port, S => 
                           SUMB_10_14_port);
   S2_10_15 : FA_X1 port map( A => ab_10_15_port, B => CARRYB_9_15_port, CI => 
                           SUMB_9_16_port, CO => CARRYB_10_15_port, S => 
                           SUMB_10_15_port);
   S2_10_16 : FA_X1 port map( A => ab_10_16_port, B => CARRYB_9_16_port, CI => 
                           SUMB_9_17_port, CO => CARRYB_10_16_port, S => 
                           SUMB_10_16_port);
   S2_10_17 : FA_X1 port map( A => ab_10_17_port, B => CARRYB_9_17_port, CI => 
                           SUMB_9_18_port, CO => CARRYB_10_17_port, S => 
                           SUMB_10_17_port);
   S2_10_18 : FA_X1 port map( A => ab_10_18_port, B => CARRYB_9_18_port, CI => 
                           SUMB_9_19_port, CO => CARRYB_10_18_port, S => 
                           SUMB_10_18_port);
   S2_10_19 : FA_X1 port map( A => ab_10_19_port, B => CARRYB_9_19_port, CI => 
                           SUMB_9_20_port, CO => CARRYB_10_19_port, S => 
                           SUMB_10_19_port);
   S2_10_20 : FA_X1 port map( A => ab_10_20_port, B => CARRYB_9_20_port, CI => 
                           SUMB_9_21_port, CO => CARRYB_10_20_port, S => 
                           SUMB_10_20_port);
   S2_10_21 : FA_X1 port map( A => ab_10_21_port, B => CARRYB_9_21_port, CI => 
                           SUMB_9_22_port, CO => CARRYB_10_21_port, S => 
                           SUMB_10_21_port);
   S2_10_22 : FA_X1 port map( A => ab_10_22_port, B => CARRYB_9_22_port, CI => 
                           SUMB_9_23_port, CO => CARRYB_10_22_port, S => 
                           SUMB_10_22_port);
   S2_10_23 : FA_X1 port map( A => ab_10_23_port, B => CARRYB_9_23_port, CI => 
                           SUMB_9_24_port, CO => CARRYB_10_23_port, S => 
                           SUMB_10_23_port);
   S2_10_24 : FA_X1 port map( A => ab_10_24_port, B => CARRYB_9_24_port, CI => 
                           SUMB_9_25_port, CO => CARRYB_10_24_port, S => 
                           SUMB_10_24_port);
   S2_10_25 : FA_X1 port map( A => ab_10_25_port, B => CARRYB_9_25_port, CI => 
                           SUMB_9_26_port, CO => CARRYB_10_25_port, S => 
                           SUMB_10_25_port);
   S2_10_26 : FA_X1 port map( A => ab_10_26_port, B => CARRYB_9_26_port, CI => 
                           SUMB_9_27_port, CO => CARRYB_10_26_port, S => 
                           SUMB_10_26_port);
   S2_10_27 : FA_X1 port map( A => ab_10_27_port, B => CARRYB_9_27_port, CI => 
                           SUMB_9_28_port, CO => CARRYB_10_27_port, S => 
                           SUMB_10_27_port);
   S2_10_28 : FA_X1 port map( A => ab_10_28_port, B => CARRYB_9_28_port, CI => 
                           SUMB_9_29_port, CO => CARRYB_10_28_port, S => 
                           SUMB_10_28_port);
   S2_10_29 : FA_X1 port map( A => ab_10_29_port, B => CARRYB_9_29_port, CI => 
                           SUMB_9_30_port, CO => CARRYB_10_29_port, S => 
                           SUMB_10_29_port);
   S3_10_30 : FA_X1 port map( A => ab_10_30_port, B => CARRYB_9_30_port, CI => 
                           ab_9_31_port, CO => CARRYB_10_30_port, S => 
                           SUMB_10_30_port);
   S1_9_0 : FA_X1 port map( A => ab_9_0_port, B => CARRYB_8_0_port, CI => 
                           SUMB_8_1_port, CO => CARRYB_9_0_port, S => A1_7_port
                           );
   S2_9_1 : FA_X1 port map( A => ab_9_1_port, B => CARRYB_8_1_port, CI => 
                           SUMB_8_2_port, CO => CARRYB_9_1_port, S => 
                           SUMB_9_1_port);
   S2_9_2 : FA_X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, CI => 
                           SUMB_8_3_port, CO => CARRYB_9_2_port, S => 
                           SUMB_9_2_port);
   S2_9_3 : FA_X1 port map( A => ab_9_3_port, B => CARRYB_8_3_port, CI => 
                           SUMB_8_4_port, CO => CARRYB_9_3_port, S => 
                           SUMB_9_3_port);
   S2_9_4 : FA_X1 port map( A => ab_9_4_port, B => CARRYB_8_4_port, CI => 
                           SUMB_8_5_port, CO => CARRYB_9_4_port, S => 
                           SUMB_9_4_port);
   S2_9_5 : FA_X1 port map( A => ab_9_5_port, B => CARRYB_8_5_port, CI => 
                           SUMB_8_6_port, CO => CARRYB_9_5_port, S => 
                           SUMB_9_5_port);
   S2_9_6 : FA_X1 port map( A => ab_9_6_port, B => CARRYB_8_6_port, CI => 
                           SUMB_8_7_port, CO => CARRYB_9_6_port, S => 
                           SUMB_9_6_port);
   S2_9_7 : FA_X1 port map( A => ab_9_7_port, B => CARRYB_8_7_port, CI => 
                           SUMB_8_8_port, CO => CARRYB_9_7_port, S => 
                           SUMB_9_7_port);
   S2_9_8 : FA_X1 port map( A => ab_9_8_port, B => CARRYB_8_8_port, CI => 
                           SUMB_8_9_port, CO => CARRYB_9_8_port, S => 
                           SUMB_9_8_port);
   S2_9_9 : FA_X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, CI => 
                           SUMB_8_10_port, CO => CARRYB_9_9_port, S => 
                           SUMB_9_9_port);
   S2_9_10 : FA_X1 port map( A => ab_9_10_port, B => CARRYB_8_10_port, CI => 
                           SUMB_8_11_port, CO => CARRYB_9_10_port, S => 
                           SUMB_9_10_port);
   S2_9_11 : FA_X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, CI => 
                           SUMB_8_12_port, CO => CARRYB_9_11_port, S => 
                           SUMB_9_11_port);
   S2_9_12 : FA_X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, CI => 
                           SUMB_8_13_port, CO => CARRYB_9_12_port, S => 
                           SUMB_9_12_port);
   S2_9_13 : FA_X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, CI => 
                           SUMB_8_14_port, CO => CARRYB_9_13_port, S => 
                           SUMB_9_13_port);
   S2_9_14 : FA_X1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, CI => 
                           SUMB_8_15_port, CO => CARRYB_9_14_port, S => 
                           SUMB_9_14_port);
   S2_9_15 : FA_X1 port map( A => ab_9_15_port, B => CARRYB_8_15_port, CI => 
                           SUMB_8_16_port, CO => CARRYB_9_15_port, S => 
                           SUMB_9_15_port);
   S2_9_16 : FA_X1 port map( A => ab_9_16_port, B => CARRYB_8_16_port, CI => 
                           SUMB_8_17_port, CO => CARRYB_9_16_port, S => 
                           SUMB_9_16_port);
   S2_9_17 : FA_X1 port map( A => ab_9_17_port, B => CARRYB_8_17_port, CI => 
                           SUMB_8_18_port, CO => CARRYB_9_17_port, S => 
                           SUMB_9_17_port);
   S2_9_18 : FA_X1 port map( A => ab_9_18_port, B => CARRYB_8_18_port, CI => 
                           SUMB_8_19_port, CO => CARRYB_9_18_port, S => 
                           SUMB_9_18_port);
   S2_9_19 : FA_X1 port map( A => ab_9_19_port, B => CARRYB_8_19_port, CI => 
                           SUMB_8_20_port, CO => CARRYB_9_19_port, S => 
                           SUMB_9_19_port);
   S2_9_20 : FA_X1 port map( A => ab_9_20_port, B => CARRYB_8_20_port, CI => 
                           SUMB_8_21_port, CO => CARRYB_9_20_port, S => 
                           SUMB_9_20_port);
   S2_9_21 : FA_X1 port map( A => ab_9_21_port, B => CARRYB_8_21_port, CI => 
                           SUMB_8_22_port, CO => CARRYB_9_21_port, S => 
                           SUMB_9_21_port);
   S2_9_22 : FA_X1 port map( A => ab_9_22_port, B => CARRYB_8_22_port, CI => 
                           SUMB_8_23_port, CO => CARRYB_9_22_port, S => 
                           SUMB_9_22_port);
   S2_9_23 : FA_X1 port map( A => ab_9_23_port, B => CARRYB_8_23_port, CI => 
                           SUMB_8_24_port, CO => CARRYB_9_23_port, S => 
                           SUMB_9_23_port);
   S2_9_24 : FA_X1 port map( A => ab_9_24_port, B => CARRYB_8_24_port, CI => 
                           SUMB_8_25_port, CO => CARRYB_9_24_port, S => 
                           SUMB_9_24_port);
   S2_9_25 : FA_X1 port map( A => ab_9_25_port, B => CARRYB_8_25_port, CI => 
                           SUMB_8_26_port, CO => CARRYB_9_25_port, S => 
                           SUMB_9_25_port);
   S2_9_26 : FA_X1 port map( A => ab_9_26_port, B => CARRYB_8_26_port, CI => 
                           SUMB_8_27_port, CO => CARRYB_9_26_port, S => 
                           SUMB_9_26_port);
   S2_9_27 : FA_X1 port map( A => ab_9_27_port, B => CARRYB_8_27_port, CI => 
                           SUMB_8_28_port, CO => CARRYB_9_27_port, S => 
                           SUMB_9_27_port);
   S2_9_28 : FA_X1 port map( A => ab_9_28_port, B => CARRYB_8_28_port, CI => 
                           SUMB_8_29_port, CO => CARRYB_9_28_port, S => 
                           SUMB_9_28_port);
   S2_9_29 : FA_X1 port map( A => ab_9_29_port, B => CARRYB_8_29_port, CI => 
                           SUMB_8_30_port, CO => CARRYB_9_29_port, S => 
                           SUMB_9_29_port);
   S3_9_30 : FA_X1 port map( A => ab_9_30_port, B => CARRYB_8_30_port, CI => 
                           ab_8_31_port, CO => CARRYB_9_30_port, S => 
                           SUMB_9_30_port);
   S1_8_0 : FA_X1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, CI => 
                           SUMB_7_1_port, CO => CARRYB_8_0_port, S => A1_6_port
                           );
   S2_8_1 : FA_X1 port map( A => ab_8_1_port, B => CARRYB_7_1_port, CI => 
                           SUMB_7_2_port, CO => CARRYB_8_1_port, S => 
                           SUMB_8_1_port);
   S2_8_2 : FA_X1 port map( A => ab_8_2_port, B => CARRYB_7_2_port, CI => 
                           SUMB_7_3_port, CO => CARRYB_8_2_port, S => 
                           SUMB_8_2_port);
   S2_8_3 : FA_X1 port map( A => ab_8_3_port, B => CARRYB_7_3_port, CI => 
                           SUMB_7_4_port, CO => CARRYB_8_3_port, S => 
                           SUMB_8_3_port);
   S2_8_4 : FA_X1 port map( A => ab_8_4_port, B => CARRYB_7_4_port, CI => 
                           SUMB_7_5_port, CO => CARRYB_8_4_port, S => 
                           SUMB_8_4_port);
   S2_8_5 : FA_X1 port map( A => ab_8_5_port, B => CARRYB_7_5_port, CI => 
                           SUMB_7_6_port, CO => CARRYB_8_5_port, S => 
                           SUMB_8_5_port);
   S2_8_6 : FA_X1 port map( A => ab_8_6_port, B => CARRYB_7_6_port, CI => 
                           SUMB_7_7_port, CO => CARRYB_8_6_port, S => 
                           SUMB_8_6_port);
   S2_8_7 : FA_X1 port map( A => ab_8_7_port, B => CARRYB_7_7_port, CI => 
                           SUMB_7_8_port, CO => CARRYB_8_7_port, S => 
                           SUMB_8_7_port);
   S2_8_8 : FA_X1 port map( A => ab_8_8_port, B => CARRYB_7_8_port, CI => 
                           SUMB_7_9_port, CO => CARRYB_8_8_port, S => 
                           SUMB_8_8_port);
   S2_8_9 : FA_X1 port map( A => ab_8_9_port, B => CARRYB_7_9_port, CI => 
                           SUMB_7_10_port, CO => CARRYB_8_9_port, S => 
                           SUMB_8_9_port);
   S2_8_10 : FA_X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, CI => 
                           SUMB_7_11_port, CO => CARRYB_8_10_port, S => 
                           SUMB_8_10_port);
   S2_8_11 : FA_X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, CI => 
                           SUMB_7_12_port, CO => CARRYB_8_11_port, S => 
                           SUMB_8_11_port);
   S2_8_12 : FA_X1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, CI => 
                           SUMB_7_13_port, CO => CARRYB_8_12_port, S => 
                           SUMB_8_12_port);
   S2_8_13 : FA_X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, CI => 
                           SUMB_7_14_port, CO => CARRYB_8_13_port, S => 
                           SUMB_8_13_port);
   S2_8_14 : FA_X1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, CI => 
                           SUMB_7_15_port, CO => CARRYB_8_14_port, S => 
                           SUMB_8_14_port);
   S2_8_15 : FA_X1 port map( A => ab_8_15_port, B => CARRYB_7_15_port, CI => 
                           SUMB_7_16_port, CO => CARRYB_8_15_port, S => 
                           SUMB_8_15_port);
   S2_8_16 : FA_X1 port map( A => ab_8_16_port, B => CARRYB_7_16_port, CI => 
                           SUMB_7_17_port, CO => CARRYB_8_16_port, S => 
                           SUMB_8_16_port);
   S2_8_17 : FA_X1 port map( A => ab_8_17_port, B => CARRYB_7_17_port, CI => 
                           SUMB_7_18_port, CO => CARRYB_8_17_port, S => 
                           SUMB_8_17_port);
   S2_8_18 : FA_X1 port map( A => ab_8_18_port, B => CARRYB_7_18_port, CI => 
                           SUMB_7_19_port, CO => CARRYB_8_18_port, S => 
                           SUMB_8_18_port);
   S2_8_19 : FA_X1 port map( A => ab_8_19_port, B => CARRYB_7_19_port, CI => 
                           SUMB_7_20_port, CO => CARRYB_8_19_port, S => 
                           SUMB_8_19_port);
   S2_8_20 : FA_X1 port map( A => ab_8_20_port, B => CARRYB_7_20_port, CI => 
                           SUMB_7_21_port, CO => CARRYB_8_20_port, S => 
                           SUMB_8_20_port);
   S2_8_21 : FA_X1 port map( A => ab_8_21_port, B => CARRYB_7_21_port, CI => 
                           SUMB_7_22_port, CO => CARRYB_8_21_port, S => 
                           SUMB_8_21_port);
   S2_8_22 : FA_X1 port map( A => ab_8_22_port, B => CARRYB_7_22_port, CI => 
                           SUMB_7_23_port, CO => CARRYB_8_22_port, S => 
                           SUMB_8_22_port);
   S2_8_23 : FA_X1 port map( A => ab_8_23_port, B => CARRYB_7_23_port, CI => 
                           SUMB_7_24_port, CO => CARRYB_8_23_port, S => 
                           SUMB_8_23_port);
   S2_8_24 : FA_X1 port map( A => ab_8_24_port, B => CARRYB_7_24_port, CI => 
                           SUMB_7_25_port, CO => CARRYB_8_24_port, S => 
                           SUMB_8_24_port);
   S2_8_25 : FA_X1 port map( A => ab_8_25_port, B => CARRYB_7_25_port, CI => 
                           SUMB_7_26_port, CO => CARRYB_8_25_port, S => 
                           SUMB_8_25_port);
   S2_8_26 : FA_X1 port map( A => ab_8_26_port, B => CARRYB_7_26_port, CI => 
                           SUMB_7_27_port, CO => CARRYB_8_26_port, S => 
                           SUMB_8_26_port);
   S2_8_27 : FA_X1 port map( A => ab_8_27_port, B => CARRYB_7_27_port, CI => 
                           SUMB_7_28_port, CO => CARRYB_8_27_port, S => 
                           SUMB_8_27_port);
   S2_8_28 : FA_X1 port map( A => ab_8_28_port, B => CARRYB_7_28_port, CI => 
                           SUMB_7_29_port, CO => CARRYB_8_28_port, S => 
                           SUMB_8_28_port);
   S2_8_29 : FA_X1 port map( A => ab_8_29_port, B => CARRYB_7_29_port, CI => 
                           SUMB_7_30_port, CO => CARRYB_8_29_port, S => 
                           SUMB_8_29_port);
   S3_8_30 : FA_X1 port map( A => ab_8_30_port, B => CARRYB_7_30_port, CI => 
                           ab_7_31_port, CO => CARRYB_8_30_port, S => 
                           SUMB_8_30_port);
   S1_7_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => A1_5_port
                           );
   S2_7_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S2_7_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S2_7_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S2_7_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S2_7_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S2_7_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           SUMB_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S2_7_7 : FA_X1 port map( A => ab_7_7_port, B => CARRYB_6_7_port, CI => 
                           SUMB_6_8_port, CO => CARRYB_7_7_port, S => 
                           SUMB_7_7_port);
   S2_7_8 : FA_X1 port map( A => ab_7_8_port, B => CARRYB_6_8_port, CI => 
                           SUMB_6_9_port, CO => CARRYB_7_8_port, S => 
                           SUMB_7_8_port);
   S2_7_9 : FA_X1 port map( A => ab_7_9_port, B => CARRYB_6_9_port, CI => 
                           SUMB_6_10_port, CO => CARRYB_7_9_port, S => 
                           SUMB_7_9_port);
   S2_7_10 : FA_X1 port map( A => ab_7_10_port, B => CARRYB_6_10_port, CI => 
                           SUMB_6_11_port, CO => CARRYB_7_10_port, S => 
                           SUMB_7_10_port);
   S2_7_11 : FA_X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, CI => 
                           SUMB_6_12_port, CO => CARRYB_7_11_port, S => 
                           SUMB_7_11_port);
   S2_7_12 : FA_X1 port map( A => ab_7_12_port, B => CARRYB_6_12_port, CI => 
                           SUMB_6_13_port, CO => CARRYB_7_12_port, S => 
                           SUMB_7_12_port);
   S2_7_13 : FA_X1 port map( A => ab_7_13_port, B => CARRYB_6_13_port, CI => 
                           SUMB_6_14_port, CO => CARRYB_7_13_port, S => 
                           SUMB_7_13_port);
   S2_7_14 : FA_X1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, CI => 
                           SUMB_6_15_port, CO => CARRYB_7_14_port, S => 
                           SUMB_7_14_port);
   S2_7_15 : FA_X1 port map( A => ab_7_15_port, B => CARRYB_6_15_port, CI => 
                           SUMB_6_16_port, CO => CARRYB_7_15_port, S => 
                           SUMB_7_15_port);
   S2_7_16 : FA_X1 port map( A => ab_7_16_port, B => CARRYB_6_16_port, CI => 
                           SUMB_6_17_port, CO => CARRYB_7_16_port, S => 
                           SUMB_7_16_port);
   S2_7_17 : FA_X1 port map( A => ab_7_17_port, B => CARRYB_6_17_port, CI => 
                           SUMB_6_18_port, CO => CARRYB_7_17_port, S => 
                           SUMB_7_17_port);
   S2_7_18 : FA_X1 port map( A => ab_7_18_port, B => CARRYB_6_18_port, CI => 
                           SUMB_6_19_port, CO => CARRYB_7_18_port, S => 
                           SUMB_7_18_port);
   S2_7_19 : FA_X1 port map( A => ab_7_19_port, B => CARRYB_6_19_port, CI => 
                           SUMB_6_20_port, CO => CARRYB_7_19_port, S => 
                           SUMB_7_19_port);
   S2_7_20 : FA_X1 port map( A => ab_7_20_port, B => CARRYB_6_20_port, CI => 
                           SUMB_6_21_port, CO => CARRYB_7_20_port, S => 
                           SUMB_7_20_port);
   S2_7_21 : FA_X1 port map( A => ab_7_21_port, B => CARRYB_6_21_port, CI => 
                           SUMB_6_22_port, CO => CARRYB_7_21_port, S => 
                           SUMB_7_21_port);
   S2_7_22 : FA_X1 port map( A => ab_7_22_port, B => CARRYB_6_22_port, CI => 
                           SUMB_6_23_port, CO => CARRYB_7_22_port, S => 
                           SUMB_7_22_port);
   S2_7_23 : FA_X1 port map( A => ab_7_23_port, B => CARRYB_6_23_port, CI => 
                           SUMB_6_24_port, CO => CARRYB_7_23_port, S => 
                           SUMB_7_23_port);
   S2_7_24 : FA_X1 port map( A => ab_7_24_port, B => CARRYB_6_24_port, CI => 
                           SUMB_6_25_port, CO => CARRYB_7_24_port, S => 
                           SUMB_7_24_port);
   S2_7_25 : FA_X1 port map( A => ab_7_25_port, B => CARRYB_6_25_port, CI => 
                           SUMB_6_26_port, CO => CARRYB_7_25_port, S => 
                           SUMB_7_25_port);
   S2_7_26 : FA_X1 port map( A => ab_7_26_port, B => CARRYB_6_26_port, CI => 
                           SUMB_6_27_port, CO => CARRYB_7_26_port, S => 
                           SUMB_7_26_port);
   S2_7_27 : FA_X1 port map( A => ab_7_27_port, B => CARRYB_6_27_port, CI => 
                           SUMB_6_28_port, CO => CARRYB_7_27_port, S => 
                           SUMB_7_27_port);
   S2_7_28 : FA_X1 port map( A => ab_7_28_port, B => CARRYB_6_28_port, CI => 
                           SUMB_6_29_port, CO => CARRYB_7_28_port, S => 
                           SUMB_7_28_port);
   S2_7_29 : FA_X1 port map( A => ab_7_29_port, B => CARRYB_6_29_port, CI => 
                           SUMB_6_30_port, CO => CARRYB_7_29_port, S => 
                           SUMB_7_29_port);
   S3_7_30 : FA_X1 port map( A => ab_7_30_port, B => CARRYB_6_30_port, CI => 
                           ab_6_31_port, CO => CARRYB_7_30_port, S => 
                           SUMB_7_30_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S2_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           SUMB_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S2_6_7 : FA_X1 port map( A => ab_6_7_port, B => CARRYB_5_7_port, CI => 
                           SUMB_5_8_port, CO => CARRYB_6_7_port, S => 
                           SUMB_6_7_port);
   S2_6_8 : FA_X1 port map( A => ab_6_8_port, B => CARRYB_5_8_port, CI => 
                           SUMB_5_9_port, CO => CARRYB_6_8_port, S => 
                           SUMB_6_8_port);
   S2_6_9 : FA_X1 port map( A => ab_6_9_port, B => CARRYB_5_9_port, CI => 
                           SUMB_5_10_port, CO => CARRYB_6_9_port, S => 
                           SUMB_6_9_port);
   S2_6_10 : FA_X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, CI => 
                           SUMB_5_11_port, CO => CARRYB_6_10_port, S => 
                           SUMB_6_10_port);
   S2_6_11 : FA_X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, CI => 
                           SUMB_5_12_port, CO => CARRYB_6_11_port, S => 
                           SUMB_6_11_port);
   S2_6_12 : FA_X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, CI => 
                           SUMB_5_13_port, CO => CARRYB_6_12_port, S => 
                           SUMB_6_12_port);
   S2_6_13 : FA_X1 port map( A => ab_6_13_port, B => CARRYB_5_13_port, CI => 
                           SUMB_5_14_port, CO => CARRYB_6_13_port, S => 
                           SUMB_6_13_port);
   S2_6_14 : FA_X1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, CI => 
                           SUMB_5_15_port, CO => CARRYB_6_14_port, S => 
                           SUMB_6_14_port);
   S2_6_15 : FA_X1 port map( A => ab_6_15_port, B => CARRYB_5_15_port, CI => 
                           SUMB_5_16_port, CO => CARRYB_6_15_port, S => 
                           SUMB_6_15_port);
   S2_6_16 : FA_X1 port map( A => ab_6_16_port, B => CARRYB_5_16_port, CI => 
                           SUMB_5_17_port, CO => CARRYB_6_16_port, S => 
                           SUMB_6_16_port);
   S2_6_17 : FA_X1 port map( A => ab_6_17_port, B => CARRYB_5_17_port, CI => 
                           SUMB_5_18_port, CO => CARRYB_6_17_port, S => 
                           SUMB_6_17_port);
   S2_6_18 : FA_X1 port map( A => ab_6_18_port, B => CARRYB_5_18_port, CI => 
                           SUMB_5_19_port, CO => CARRYB_6_18_port, S => 
                           SUMB_6_18_port);
   S2_6_19 : FA_X1 port map( A => ab_6_19_port, B => CARRYB_5_19_port, CI => 
                           SUMB_5_20_port, CO => CARRYB_6_19_port, S => 
                           SUMB_6_19_port);
   S2_6_20 : FA_X1 port map( A => ab_6_20_port, B => CARRYB_5_20_port, CI => 
                           SUMB_5_21_port, CO => CARRYB_6_20_port, S => 
                           SUMB_6_20_port);
   S2_6_21 : FA_X1 port map( A => ab_6_21_port, B => CARRYB_5_21_port, CI => 
                           SUMB_5_22_port, CO => CARRYB_6_21_port, S => 
                           SUMB_6_21_port);
   S2_6_22 : FA_X1 port map( A => ab_6_22_port, B => CARRYB_5_22_port, CI => 
                           SUMB_5_23_port, CO => CARRYB_6_22_port, S => 
                           SUMB_6_22_port);
   S2_6_23 : FA_X1 port map( A => ab_6_23_port, B => CARRYB_5_23_port, CI => 
                           SUMB_5_24_port, CO => CARRYB_6_23_port, S => 
                           SUMB_6_23_port);
   S2_6_24 : FA_X1 port map( A => ab_6_24_port, B => CARRYB_5_24_port, CI => 
                           SUMB_5_25_port, CO => CARRYB_6_24_port, S => 
                           SUMB_6_24_port);
   S2_6_25 : FA_X1 port map( A => ab_6_25_port, B => CARRYB_5_25_port, CI => 
                           SUMB_5_26_port, CO => CARRYB_6_25_port, S => 
                           SUMB_6_25_port);
   S2_6_26 : FA_X1 port map( A => ab_6_26_port, B => CARRYB_5_26_port, CI => 
                           SUMB_5_27_port, CO => CARRYB_6_26_port, S => 
                           SUMB_6_26_port);
   S2_6_27 : FA_X1 port map( A => ab_6_27_port, B => CARRYB_5_27_port, CI => 
                           SUMB_5_28_port, CO => CARRYB_6_27_port, S => 
                           SUMB_6_27_port);
   S2_6_28 : FA_X1 port map( A => ab_6_28_port, B => CARRYB_5_28_port, CI => 
                           SUMB_5_29_port, CO => CARRYB_6_28_port, S => 
                           SUMB_6_28_port);
   S2_6_29 : FA_X1 port map( A => ab_6_29_port, B => CARRYB_5_29_port, CI => 
                           SUMB_5_30_port, CO => CARRYB_6_29_port, S => 
                           SUMB_6_29_port);
   S3_6_30 : FA_X1 port map( A => ab_6_30_port, B => CARRYB_5_30_port, CI => 
                           ab_5_31_port, CO => CARRYB_6_30_port, S => 
                           SUMB_6_30_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S2_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           SUMB_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S2_5_7 : FA_X1 port map( A => ab_5_7_port, B => CARRYB_4_7_port, CI => 
                           SUMB_4_8_port, CO => CARRYB_5_7_port, S => 
                           SUMB_5_7_port);
   S2_5_8 : FA_X1 port map( A => ab_5_8_port, B => CARRYB_4_8_port, CI => 
                           SUMB_4_9_port, CO => CARRYB_5_8_port, S => 
                           SUMB_5_8_port);
   S2_5_9 : FA_X1 port map( A => ab_5_9_port, B => CARRYB_4_9_port, CI => 
                           SUMB_4_10_port, CO => CARRYB_5_9_port, S => 
                           SUMB_5_9_port);
   S2_5_10 : FA_X1 port map( A => ab_5_10_port, B => CARRYB_4_10_port, CI => 
                           SUMB_4_11_port, CO => CARRYB_5_10_port, S => 
                           SUMB_5_10_port);
   S2_5_11 : FA_X1 port map( A => ab_5_11_port, B => CARRYB_4_11_port, CI => 
                           SUMB_4_12_port, CO => CARRYB_5_11_port, S => 
                           SUMB_5_11_port);
   S2_5_12 : FA_X1 port map( A => ab_5_12_port, B => CARRYB_4_12_port, CI => 
                           SUMB_4_13_port, CO => CARRYB_5_12_port, S => 
                           SUMB_5_12_port);
   S2_5_13 : FA_X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, CI => 
                           SUMB_4_14_port, CO => CARRYB_5_13_port, S => 
                           SUMB_5_13_port);
   S2_5_14 : FA_X1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, CI => 
                           SUMB_4_15_port, CO => CARRYB_5_14_port, S => 
                           SUMB_5_14_port);
   S2_5_15 : FA_X1 port map( A => ab_5_15_port, B => CARRYB_4_15_port, CI => 
                           SUMB_4_16_port, CO => CARRYB_5_15_port, S => 
                           SUMB_5_15_port);
   S2_5_16 : FA_X1 port map( A => ab_5_16_port, B => CARRYB_4_16_port, CI => 
                           SUMB_4_17_port, CO => CARRYB_5_16_port, S => 
                           SUMB_5_16_port);
   S2_5_17 : FA_X1 port map( A => ab_5_17_port, B => CARRYB_4_17_port, CI => 
                           SUMB_4_18_port, CO => CARRYB_5_17_port, S => 
                           SUMB_5_17_port);
   S2_5_18 : FA_X1 port map( A => ab_5_18_port, B => CARRYB_4_18_port, CI => 
                           SUMB_4_19_port, CO => CARRYB_5_18_port, S => 
                           SUMB_5_18_port);
   S2_5_19 : FA_X1 port map( A => ab_5_19_port, B => CARRYB_4_19_port, CI => 
                           SUMB_4_20_port, CO => CARRYB_5_19_port, S => 
                           SUMB_5_19_port);
   S2_5_20 : FA_X1 port map( A => ab_5_20_port, B => CARRYB_4_20_port, CI => 
                           SUMB_4_21_port, CO => CARRYB_5_20_port, S => 
                           SUMB_5_20_port);
   S2_5_21 : FA_X1 port map( A => ab_5_21_port, B => CARRYB_4_21_port, CI => 
                           SUMB_4_22_port, CO => CARRYB_5_21_port, S => 
                           SUMB_5_21_port);
   S2_5_22 : FA_X1 port map( A => ab_5_22_port, B => CARRYB_4_22_port, CI => 
                           SUMB_4_23_port, CO => CARRYB_5_22_port, S => 
                           SUMB_5_22_port);
   S2_5_23 : FA_X1 port map( A => ab_5_23_port, B => CARRYB_4_23_port, CI => 
                           SUMB_4_24_port, CO => CARRYB_5_23_port, S => 
                           SUMB_5_23_port);
   S2_5_24 : FA_X1 port map( A => ab_5_24_port, B => CARRYB_4_24_port, CI => 
                           SUMB_4_25_port, CO => CARRYB_5_24_port, S => 
                           SUMB_5_24_port);
   S2_5_25 : FA_X1 port map( A => ab_5_25_port, B => CARRYB_4_25_port, CI => 
                           SUMB_4_26_port, CO => CARRYB_5_25_port, S => 
                           SUMB_5_25_port);
   S2_5_26 : FA_X1 port map( A => ab_5_26_port, B => CARRYB_4_26_port, CI => 
                           SUMB_4_27_port, CO => CARRYB_5_26_port, S => 
                           SUMB_5_26_port);
   S2_5_27 : FA_X1 port map( A => ab_5_27_port, B => CARRYB_4_27_port, CI => 
                           SUMB_4_28_port, CO => CARRYB_5_27_port, S => 
                           SUMB_5_27_port);
   S2_5_28 : FA_X1 port map( A => ab_5_28_port, B => CARRYB_4_28_port, CI => 
                           SUMB_4_29_port, CO => CARRYB_5_28_port, S => 
                           SUMB_5_28_port);
   S2_5_29 : FA_X1 port map( A => ab_5_29_port, B => CARRYB_4_29_port, CI => 
                           SUMB_4_30_port, CO => CARRYB_5_29_port, S => 
                           SUMB_5_29_port);
   S3_5_30 : FA_X1 port map( A => ab_5_30_port, B => CARRYB_4_30_port, CI => 
                           ab_4_31_port, CO => CARRYB_5_30_port, S => 
                           SUMB_5_30_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S2_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           SUMB_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S2_4_7 : FA_X1 port map( A => ab_4_7_port, B => CARRYB_3_7_port, CI => 
                           SUMB_3_8_port, CO => CARRYB_4_7_port, S => 
                           SUMB_4_7_port);
   S2_4_8 : FA_X1 port map( A => ab_4_8_port, B => CARRYB_3_8_port, CI => 
                           SUMB_3_9_port, CO => CARRYB_4_8_port, S => 
                           SUMB_4_8_port);
   S2_4_9 : FA_X1 port map( A => ab_4_9_port, B => CARRYB_3_9_port, CI => 
                           SUMB_3_10_port, CO => CARRYB_4_9_port, S => 
                           SUMB_4_9_port);
   S2_4_10 : FA_X1 port map( A => ab_4_10_port, B => CARRYB_3_10_port, CI => 
                           SUMB_3_11_port, CO => CARRYB_4_10_port, S => 
                           SUMB_4_10_port);
   S2_4_11 : FA_X1 port map( A => ab_4_11_port, B => CARRYB_3_11_port, CI => 
                           SUMB_3_12_port, CO => CARRYB_4_11_port, S => 
                           SUMB_4_11_port);
   S2_4_12 : FA_X1 port map( A => ab_4_12_port, B => CARRYB_3_12_port, CI => 
                           SUMB_3_13_port, CO => CARRYB_4_12_port, S => 
                           SUMB_4_12_port);
   S2_4_13 : FA_X1 port map( A => ab_4_13_port, B => CARRYB_3_13_port, CI => 
                           SUMB_3_14_port, CO => CARRYB_4_13_port, S => 
                           SUMB_4_13_port);
   S2_4_14 : FA_X1 port map( A => ab_4_14_port, B => CARRYB_3_14_port, CI => 
                           SUMB_3_15_port, CO => CARRYB_4_14_port, S => 
                           SUMB_4_14_port);
   S2_4_15 : FA_X1 port map( A => ab_4_15_port, B => CARRYB_3_15_port, CI => 
                           SUMB_3_16_port, CO => CARRYB_4_15_port, S => 
                           SUMB_4_15_port);
   S2_4_16 : FA_X1 port map( A => ab_4_16_port, B => CARRYB_3_16_port, CI => 
                           SUMB_3_17_port, CO => CARRYB_4_16_port, S => 
                           SUMB_4_16_port);
   S2_4_17 : FA_X1 port map( A => ab_4_17_port, B => CARRYB_3_17_port, CI => 
                           SUMB_3_18_port, CO => CARRYB_4_17_port, S => 
                           SUMB_4_17_port);
   S2_4_18 : FA_X1 port map( A => ab_4_18_port, B => CARRYB_3_18_port, CI => 
                           SUMB_3_19_port, CO => CARRYB_4_18_port, S => 
                           SUMB_4_18_port);
   S2_4_19 : FA_X1 port map( A => ab_4_19_port, B => CARRYB_3_19_port, CI => 
                           SUMB_3_20_port, CO => CARRYB_4_19_port, S => 
                           SUMB_4_19_port);
   S2_4_20 : FA_X1 port map( A => ab_4_20_port, B => CARRYB_3_20_port, CI => 
                           SUMB_3_21_port, CO => CARRYB_4_20_port, S => 
                           SUMB_4_20_port);
   S2_4_21 : FA_X1 port map( A => ab_4_21_port, B => CARRYB_3_21_port, CI => 
                           SUMB_3_22_port, CO => CARRYB_4_21_port, S => 
                           SUMB_4_21_port);
   S2_4_22 : FA_X1 port map( A => ab_4_22_port, B => CARRYB_3_22_port, CI => 
                           SUMB_3_23_port, CO => CARRYB_4_22_port, S => 
                           SUMB_4_22_port);
   S2_4_23 : FA_X1 port map( A => ab_4_23_port, B => CARRYB_3_23_port, CI => 
                           SUMB_3_24_port, CO => CARRYB_4_23_port, S => 
                           SUMB_4_23_port);
   S2_4_24 : FA_X1 port map( A => ab_4_24_port, B => CARRYB_3_24_port, CI => 
                           SUMB_3_25_port, CO => CARRYB_4_24_port, S => 
                           SUMB_4_24_port);
   S2_4_25 : FA_X1 port map( A => ab_4_25_port, B => CARRYB_3_25_port, CI => 
                           SUMB_3_26_port, CO => CARRYB_4_25_port, S => 
                           SUMB_4_25_port);
   S2_4_26 : FA_X1 port map( A => ab_4_26_port, B => CARRYB_3_26_port, CI => 
                           SUMB_3_27_port, CO => CARRYB_4_26_port, S => 
                           SUMB_4_26_port);
   S2_4_27 : FA_X1 port map( A => ab_4_27_port, B => CARRYB_3_27_port, CI => 
                           SUMB_3_28_port, CO => CARRYB_4_27_port, S => 
                           SUMB_4_27_port);
   S2_4_28 : FA_X1 port map( A => ab_4_28_port, B => CARRYB_3_28_port, CI => 
                           SUMB_3_29_port, CO => CARRYB_4_28_port, S => 
                           SUMB_4_28_port);
   S2_4_29 : FA_X1 port map( A => ab_4_29_port, B => CARRYB_3_29_port, CI => 
                           SUMB_3_30_port, CO => CARRYB_4_29_port, S => 
                           SUMB_4_29_port);
   S3_4_30 : FA_X1 port map( A => ab_4_30_port, B => CARRYB_3_30_port, CI => 
                           ab_3_31_port, CO => CARRYB_4_30_port, S => 
                           SUMB_4_30_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S2_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           SUMB_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S2_3_7 : FA_X1 port map( A => ab_3_7_port, B => CARRYB_2_7_port, CI => 
                           SUMB_2_8_port, CO => CARRYB_3_7_port, S => 
                           SUMB_3_7_port);
   S2_3_8 : FA_X1 port map( A => ab_3_8_port, B => CARRYB_2_8_port, CI => 
                           SUMB_2_9_port, CO => CARRYB_3_8_port, S => 
                           SUMB_3_8_port);
   S2_3_9 : FA_X1 port map( A => ab_3_9_port, B => CARRYB_2_9_port, CI => 
                           SUMB_2_10_port, CO => CARRYB_3_9_port, S => 
                           SUMB_3_9_port);
   S2_3_10 : FA_X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, CI => 
                           SUMB_2_11_port, CO => CARRYB_3_10_port, S => 
                           SUMB_3_10_port);
   S2_3_11 : FA_X1 port map( A => ab_3_11_port, B => CARRYB_2_11_port, CI => 
                           SUMB_2_12_port, CO => CARRYB_3_11_port, S => 
                           SUMB_3_11_port);
   S2_3_12 : FA_X1 port map( A => ab_3_12_port, B => CARRYB_2_12_port, CI => 
                           SUMB_2_13_port, CO => CARRYB_3_12_port, S => 
                           SUMB_3_12_port);
   S2_3_13 : FA_X1 port map( A => ab_3_13_port, B => CARRYB_2_13_port, CI => 
                           SUMB_2_14_port, CO => CARRYB_3_13_port, S => 
                           SUMB_3_13_port);
   S2_3_14 : FA_X1 port map( A => ab_3_14_port, B => CARRYB_2_14_port, CI => 
                           SUMB_2_15_port, CO => CARRYB_3_14_port, S => 
                           SUMB_3_14_port);
   S2_3_15 : FA_X1 port map( A => ab_3_15_port, B => CARRYB_2_15_port, CI => 
                           SUMB_2_16_port, CO => CARRYB_3_15_port, S => 
                           SUMB_3_15_port);
   S2_3_16 : FA_X1 port map( A => ab_3_16_port, B => CARRYB_2_16_port, CI => 
                           SUMB_2_17_port, CO => CARRYB_3_16_port, S => 
                           SUMB_3_16_port);
   S2_3_17 : FA_X1 port map( A => ab_3_17_port, B => CARRYB_2_17_port, CI => 
                           SUMB_2_18_port, CO => CARRYB_3_17_port, S => 
                           SUMB_3_17_port);
   S2_3_18 : FA_X1 port map( A => ab_3_18_port, B => CARRYB_2_18_port, CI => 
                           SUMB_2_19_port, CO => CARRYB_3_18_port, S => 
                           SUMB_3_18_port);
   S2_3_19 : FA_X1 port map( A => ab_3_19_port, B => CARRYB_2_19_port, CI => 
                           SUMB_2_20_port, CO => CARRYB_3_19_port, S => 
                           SUMB_3_19_port);
   S2_3_20 : FA_X1 port map( A => ab_3_20_port, B => CARRYB_2_20_port, CI => 
                           SUMB_2_21_port, CO => CARRYB_3_20_port, S => 
                           SUMB_3_20_port);
   S2_3_21 : FA_X1 port map( A => ab_3_21_port, B => CARRYB_2_21_port, CI => 
                           SUMB_2_22_port, CO => CARRYB_3_21_port, S => 
                           SUMB_3_21_port);
   S2_3_22 : FA_X1 port map( A => ab_3_22_port, B => CARRYB_2_22_port, CI => 
                           SUMB_2_23_port, CO => CARRYB_3_22_port, S => 
                           SUMB_3_22_port);
   S2_3_23 : FA_X1 port map( A => ab_3_23_port, B => CARRYB_2_23_port, CI => 
                           SUMB_2_24_port, CO => CARRYB_3_23_port, S => 
                           SUMB_3_23_port);
   S2_3_24 : FA_X1 port map( A => ab_3_24_port, B => CARRYB_2_24_port, CI => 
                           SUMB_2_25_port, CO => CARRYB_3_24_port, S => 
                           SUMB_3_24_port);
   S2_3_25 : FA_X1 port map( A => ab_3_25_port, B => CARRYB_2_25_port, CI => 
                           SUMB_2_26_port, CO => CARRYB_3_25_port, S => 
                           SUMB_3_25_port);
   S2_3_26 : FA_X1 port map( A => ab_3_26_port, B => CARRYB_2_26_port, CI => 
                           SUMB_2_27_port, CO => CARRYB_3_26_port, S => 
                           SUMB_3_26_port);
   S2_3_27 : FA_X1 port map( A => ab_3_27_port, B => CARRYB_2_27_port, CI => 
                           SUMB_2_28_port, CO => CARRYB_3_27_port, S => 
                           SUMB_3_27_port);
   S2_3_28 : FA_X1 port map( A => ab_3_28_port, B => CARRYB_2_28_port, CI => 
                           SUMB_2_29_port, CO => CARRYB_3_28_port, S => 
                           SUMB_3_28_port);
   S2_3_29 : FA_X1 port map( A => ab_3_29_port, B => CARRYB_2_29_port, CI => 
                           SUMB_2_30_port, CO => CARRYB_3_29_port, S => 
                           SUMB_3_29_port);
   S3_3_30 : FA_X1 port map( A => ab_3_30_port, B => CARRYB_2_30_port, CI => 
                           ab_2_31_port, CO => CARRYB_3_30_port, S => 
                           SUMB_3_30_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n31, CI => n62, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n30, CI => n61, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n29, CI => n60, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n28, CI => n59, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n27, CI => n58, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n26, CI => n57, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S2_2_6 : FA_X1 port map( A => ab_2_6_port, B => n25, CI => n56, CO => 
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   S2_2_7 : FA_X1 port map( A => ab_2_7_port, B => n24, CI => n55, CO => 
                           CARRYB_2_7_port, S => SUMB_2_7_port);
   S2_2_8 : FA_X1 port map( A => ab_2_8_port, B => n23, CI => n54, CO => 
                           CARRYB_2_8_port, S => SUMB_2_8_port);
   S2_2_9 : FA_X1 port map( A => ab_2_9_port, B => n22, CI => n53, CO => 
                           CARRYB_2_9_port, S => SUMB_2_9_port);
   S2_2_10 : FA_X1 port map( A => ab_2_10_port, B => n21, CI => n52, CO => 
                           CARRYB_2_10_port, S => SUMB_2_10_port);
   S2_2_11 : FA_X1 port map( A => ab_2_11_port, B => n20, CI => n51, CO => 
                           CARRYB_2_11_port, S => SUMB_2_11_port);
   S2_2_12 : FA_X1 port map( A => ab_2_12_port, B => n19, CI => n50, CO => 
                           CARRYB_2_12_port, S => SUMB_2_12_port);
   S2_2_13 : FA_X1 port map( A => ab_2_13_port, B => n18, CI => n49, CO => 
                           CARRYB_2_13_port, S => SUMB_2_13_port);
   S2_2_14 : FA_X1 port map( A => ab_2_14_port, B => n17, CI => n48, CO => 
                           CARRYB_2_14_port, S => SUMB_2_14_port);
   S2_2_15 : FA_X1 port map( A => ab_2_15_port, B => n16, CI => n47, CO => 
                           CARRYB_2_15_port, S => SUMB_2_15_port);
   S2_2_16 : FA_X1 port map( A => ab_2_16_port, B => n15, CI => n46, CO => 
                           CARRYB_2_16_port, S => SUMB_2_16_port);
   S2_2_17 : FA_X1 port map( A => ab_2_17_port, B => n14, CI => n45, CO => 
                           CARRYB_2_17_port, S => SUMB_2_17_port);
   S2_2_18 : FA_X1 port map( A => ab_2_18_port, B => n13, CI => n44, CO => 
                           CARRYB_2_18_port, S => SUMB_2_18_port);
   S2_2_19 : FA_X1 port map( A => ab_2_19_port, B => n12, CI => n43, CO => 
                           CARRYB_2_19_port, S => SUMB_2_19_port);
   S2_2_20 : FA_X1 port map( A => ab_2_20_port, B => n11, CI => n42, CO => 
                           CARRYB_2_20_port, S => SUMB_2_20_port);
   S2_2_21 : FA_X1 port map( A => ab_2_21_port, B => n10, CI => n41, CO => 
                           CARRYB_2_21_port, S => SUMB_2_21_port);
   S2_2_22 : FA_X1 port map( A => ab_2_22_port, B => n9, CI => n40, CO => 
                           CARRYB_2_22_port, S => SUMB_2_22_port);
   S2_2_23 : FA_X1 port map( A => ab_2_23_port, B => n8, CI => n39, CO => 
                           CARRYB_2_23_port, S => SUMB_2_23_port);
   S2_2_24 : FA_X1 port map( A => ab_2_24_port, B => n7, CI => n38, CO => 
                           CARRYB_2_24_port, S => SUMB_2_24_port);
   S2_2_25 : FA_X1 port map( A => ab_2_25_port, B => n6, CI => n37, CO => 
                           CARRYB_2_25_port, S => SUMB_2_25_port);
   S2_2_26 : FA_X1 port map( A => ab_2_26_port, B => n5, CI => n36, CO => 
                           CARRYB_2_26_port, S => SUMB_2_26_port);
   S2_2_27 : FA_X1 port map( A => ab_2_27_port, B => n4, CI => n35, CO => 
                           CARRYB_2_27_port, S => SUMB_2_27_port);
   S2_2_28 : FA_X1 port map( A => ab_2_28_port, B => n3, CI => n34, CO => 
                           CARRYB_2_28_port, S => SUMB_2_28_port);
   S2_2_29 : FA_X1 port map( A => ab_2_29_port, B => n2, CI => n33, CO => 
                           CARRYB_2_29_port, S => SUMB_2_29_port);
   S3_2_30 : FA_X1 port map( A => ab_2_30_port, B => n32, CI => ab_1_31_port, 
                           CO => CARRYB_2_30_port, S => SUMB_2_30_port);
   FS_1 : ALU_N64_DW01_add_0 port map( A(61) => n190, A(60) => n63, A(59) => 
                           n109, A(58) => n75, A(57) => n108, A(56) => n74, 
                           A(55) => n107, A(54) => n73, A(53) => n106, A(52) =>
                           n72, A(51) => n105, A(50) => n71, A(49) => n104, 
                           A(48) => n70, A(47) => n81, A(46) => n111, A(45) => 
                           n80, A(44) => n103, A(43) => n69, A(42) => n102, 
                           A(41) => n67, A(40) => n68, A(39) => n79, A(38) => 
                           n110, A(37) => n78, A(36) => n66, A(35) => n64, 
                           A(34) => n101, A(33) => n77, A(32) => n65, A(31) => 
                           n76, A(30) => n125, A(29) => SUMB_31_0_port, A(28) 
                           => A1_28_port, A(27) => A1_27_port, A(26) => 
                           A1_26_port, A(25) => A1_25_port, A(24) => A1_24_port
                           , A(23) => A1_23_port, A(22) => A1_22_port, A(21) =>
                           A1_21_port, A(20) => A1_20_port, A(19) => A1_19_port
                           , A(18) => A1_18_port, A(17) => A1_17_port, A(16) =>
                           A1_16_port, A(15) => A1_15_port, A(14) => A1_14_port
                           , A(13) => A1_13_port, A(12) => A1_12_port, A(11) =>
                           A1_11_port, A(10) => A1_10_port, A(9) => A1_9_port, 
                           A(8) => A1_8_port, A(7) => A1_7_port, A(6) => 
                           A1_6_port, A(5) => A1_5_port, A(4) => A1_4_port, 
                           A(3) => A1_3_port, A(2) => A1_2_port, A(1) => 
                           A1_1_port, A(0) => A1_0_port, B(61) => n124, B(60) 
                           => n100, B(59) => n121, B(58) => n93, B(57) => n120,
                           B(56) => n92, B(55) => n119, B(54) => n91, B(53) => 
                           n118, B(52) => n90, B(51) => n117, B(50) => n89, 
                           B(49) => n116, B(48) => n88, B(47) => n99, B(46) => 
                           n123, B(45) => n98, B(44) => n115, B(43) => n87, 
                           B(42) => n114, B(41) => n85, B(40) => n86, B(39) => 
                           n97, B(38) => n122, B(37) => n96, B(36) => n84, 
                           B(35) => n82, B(34) => n113, B(33) => n95, B(32) => 
                           n83, B(31) => n94, B(30) => n190, B(29) => n191, 
                           B(28) => n191, B(27) => n191, B(26) => n191, B(25) 
                           => n191, B(24) => n191, B(23) => n191, B(22) => n191
                           , B(21) => n191, B(20) => n191, B(19) => n191, B(18)
                           => n191, B(17) => n191, B(16) => n191, B(15) => n191
                           , B(14) => n191, B(13) => n191, B(12) => n191, B(11)
                           => n191, B(10) => n191, B(9) => n191, B(8) => n191, 
                           B(7) => n191, B(6) => n191, B(5) => n191, B(4) => 
                           n191, B(3) => n191, B(2) => n191, B(1) => n191, B(0)
                           => X_Logic0_port, CI => X_Logic0_port, SUM(61) => 
                           PRODUCT(63), SUM(60) => PRODUCT(62), SUM(59) => 
                           PRODUCT(61), SUM(58) => PRODUCT(60), SUM(57) => 
                           PRODUCT(59), SUM(56) => PRODUCT(58), SUM(55) => 
                           PRODUCT(57), SUM(54) => PRODUCT(56), SUM(53) => 
                           PRODUCT(55), SUM(52) => PRODUCT(54), SUM(51) => 
                           PRODUCT(53), SUM(50) => PRODUCT(52), SUM(49) => 
                           PRODUCT(51), SUM(48) => PRODUCT(50), SUM(47) => 
                           PRODUCT(49), SUM(46) => PRODUCT(48), SUM(45) => 
                           PRODUCT(47), SUM(44) => PRODUCT(46), SUM(43) => 
                           PRODUCT(45), SUM(42) => PRODUCT(44), SUM(41) => 
                           PRODUCT(43), SUM(40) => PRODUCT(42), SUM(39) => 
                           PRODUCT(41), SUM(38) => PRODUCT(40), SUM(37) => 
                           PRODUCT(39), SUM(36) => PRODUCT(38), SUM(35) => 
                           PRODUCT(37), SUM(34) => PRODUCT(36), SUM(33) => 
                           PRODUCT(35), SUM(32) => PRODUCT(34), SUM(31) => 
                           PRODUCT(33), SUM(30) => PRODUCT(32), SUM(29) => 
                           PRODUCT(31), SUM(28) => PRODUCT(30), SUM(27) => 
                           PRODUCT(29), SUM(26) => PRODUCT(28), SUM(25) => 
                           PRODUCT(27), SUM(24) => PRODUCT(26), SUM(23) => 
                           PRODUCT(25), SUM(22) => PRODUCT(24), SUM(21) => 
                           PRODUCT(23), SUM(20) => PRODUCT(22), SUM(19) => 
                           PRODUCT(21), SUM(18) => PRODUCT(20), SUM(17) => 
                           PRODUCT(19), SUM(16) => PRODUCT(18), SUM(15) => 
                           PRODUCT(17), SUM(14) => PRODUCT(16), SUM(13) => 
                           PRODUCT(15), SUM(12) => PRODUCT(14), SUM(11) => 
                           PRODUCT(13), SUM(10) => PRODUCT(12), SUM(9) => 
                           PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7) => 
                           PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1038);
   U2 : AND2_X1 port map( A1 => ab_0_30_port, A2 => ab_1_29_port, ZN => n2);
   U3 : AND2_X1 port map( A1 => ab_0_29_port, A2 => ab_1_28_port, ZN => n3);
   U4 : AND2_X1 port map( A1 => ab_0_28_port, A2 => ab_1_27_port, ZN => n4);
   U5 : AND2_X1 port map( A1 => ab_0_27_port, A2 => ab_1_26_port, ZN => n5);
   U6 : AND2_X1 port map( A1 => ab_0_26_port, A2 => ab_1_25_port, ZN => n6);
   U7 : AND2_X1 port map( A1 => ab_0_25_port, A2 => ab_1_24_port, ZN => n7);
   U8 : AND2_X1 port map( A1 => ab_0_24_port, A2 => ab_1_23_port, ZN => n8);
   U9 : AND2_X1 port map( A1 => ab_0_23_port, A2 => ab_1_22_port, ZN => n9);
   U10 : AND2_X1 port map( A1 => ab_0_22_port, A2 => ab_1_21_port, ZN => n10);
   U11 : AND2_X1 port map( A1 => ab_0_21_port, A2 => ab_1_20_port, ZN => n11);
   U12 : AND2_X1 port map( A1 => ab_0_20_port, A2 => ab_1_19_port, ZN => n12);
   U13 : AND2_X1 port map( A1 => ab_0_19_port, A2 => ab_1_18_port, ZN => n13);
   U14 : AND2_X1 port map( A1 => ab_0_18_port, A2 => ab_1_17_port, ZN => n14);
   U15 : AND2_X1 port map( A1 => ab_0_17_port, A2 => ab_1_16_port, ZN => n15);
   U16 : AND2_X1 port map( A1 => ab_0_16_port, A2 => ab_1_15_port, ZN => n16);
   U17 : AND2_X1 port map( A1 => ab_0_15_port, A2 => ab_1_14_port, ZN => n17);
   U18 : AND2_X1 port map( A1 => ab_0_14_port, A2 => ab_1_13_port, ZN => n18);
   U19 : AND2_X1 port map( A1 => ab_0_13_port, A2 => ab_1_12_port, ZN => n19);
   U20 : AND2_X1 port map( A1 => ab_0_12_port, A2 => ab_1_11_port, ZN => n20);
   U21 : AND2_X1 port map( A1 => ab_0_11_port, A2 => ab_1_10_port, ZN => n21);
   U22 : AND2_X1 port map( A1 => ab_0_10_port, A2 => ab_1_9_port, ZN => n22);
   U23 : AND2_X1 port map( A1 => ab_0_9_port, A2 => ab_1_8_port, ZN => n23);
   U24 : AND2_X1 port map( A1 => ab_0_8_port, A2 => ab_1_7_port, ZN => n24);
   U25 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n25);
   U26 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n26);
   U27 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n27);
   U28 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n28);
   U29 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n29);
   U30 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n30);
   U31 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n31);
   U32 : AND2_X1 port map( A1 => ab_0_31_port, A2 => ab_1_30_port, ZN => n32);
   U33 : XOR2_X1 port map( A => ab_1_30_port, B => ab_0_31_port, Z => n33);
   U34 : XOR2_X1 port map( A => ab_1_29_port, B => ab_0_30_port, Z => n34);
   U35 : XOR2_X1 port map( A => ab_1_28_port, B => ab_0_29_port, Z => n35);
   U36 : XOR2_X1 port map( A => ab_1_27_port, B => ab_0_28_port, Z => n36);
   U37 : XOR2_X1 port map( A => ab_1_26_port, B => ab_0_27_port, Z => n37);
   U38 : XOR2_X1 port map( A => ab_1_25_port, B => ab_0_26_port, Z => n38);
   U39 : XOR2_X1 port map( A => ab_1_24_port, B => ab_0_25_port, Z => n39);
   U40 : XOR2_X1 port map( A => ab_1_23_port, B => ab_0_24_port, Z => n40);
   U41 : XOR2_X1 port map( A => ab_1_22_port, B => ab_0_23_port, Z => n41);
   U42 : XOR2_X1 port map( A => ab_1_21_port, B => ab_0_22_port, Z => n42);
   U43 : XOR2_X1 port map( A => ab_1_20_port, B => ab_0_21_port, Z => n43);
   U44 : XOR2_X1 port map( A => ab_1_19_port, B => ab_0_20_port, Z => n44);
   U45 : XOR2_X1 port map( A => ab_1_18_port, B => ab_0_19_port, Z => n45);
   U46 : XOR2_X1 port map( A => ab_1_17_port, B => ab_0_18_port, Z => n46);
   U47 : XOR2_X1 port map( A => ab_1_16_port, B => ab_0_17_port, Z => n47);
   U48 : XOR2_X1 port map( A => ab_1_15_port, B => ab_0_16_port, Z => n48);
   U49 : XOR2_X1 port map( A => ab_1_14_port, B => ab_0_15_port, Z => n49);
   U50 : XOR2_X1 port map( A => ab_1_13_port, B => ab_0_14_port, Z => n50);
   U51 : XOR2_X1 port map( A => ab_1_12_port, B => ab_0_13_port, Z => n51);
   U52 : XOR2_X1 port map( A => ab_1_11_port, B => ab_0_12_port, Z => n52);
   U53 : XOR2_X1 port map( A => ab_1_10_port, B => ab_0_11_port, Z => n53);
   U54 : XOR2_X1 port map( A => ab_1_9_port, B => ab_0_10_port, Z => n54);
   U55 : XOR2_X1 port map( A => ab_1_8_port, B => ab_0_9_port, Z => n55);
   U56 : XOR2_X1 port map( A => ab_1_7_port, B => ab_0_8_port, Z => n56);
   U57 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n57);
   U58 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n58);
   U59 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n59);
   U60 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n60);
   U61 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n61);
   U62 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n62);
   U63 : XOR2_X1 port map( A => CARRYB_31_30_port, B => ab_31_31_port, Z => n63
                           );
   U64 : XOR2_X1 port map( A => CARRYB_31_5_port, B => SUMB_31_6_port, Z => n64
                           );
   U65 : XOR2_X1 port map( A => CARRYB_31_2_port, B => SUMB_31_3_port, Z => n65
                           );
   U66 : XOR2_X1 port map( A => CARRYB_31_6_port, B => SUMB_31_7_port, Z => n66
                           );
   U67 : XOR2_X1 port map( A => CARRYB_31_11_port, B => SUMB_31_12_port, Z => 
                           n67);
   U68 : XOR2_X1 port map( A => CARRYB_31_10_port, B => SUMB_31_11_port, Z => 
                           n68);
   U69 : XOR2_X1 port map( A => CARRYB_31_13_port, B => SUMB_31_14_port, Z => 
                           n69);
   U70 : XOR2_X1 port map( A => CARRYB_31_18_port, B => SUMB_31_19_port, Z => 
                           n70);
   U71 : XOR2_X1 port map( A => CARRYB_31_20_port, B => SUMB_31_21_port, Z => 
                           n71);
   U72 : XOR2_X1 port map( A => CARRYB_31_22_port, B => SUMB_31_23_port, Z => 
                           n72);
   U73 : XOR2_X1 port map( A => CARRYB_31_24_port, B => SUMB_31_25_port, Z => 
                           n73);
   U74 : XOR2_X1 port map( A => CARRYB_31_26_port, B => SUMB_31_27_port, Z => 
                           n74);
   U75 : XOR2_X1 port map( A => CARRYB_31_28_port, B => SUMB_31_29_port, Z => 
                           n75);
   U76 : XOR2_X1 port map( A => CARRYB_31_1_port, B => SUMB_31_2_port, Z => n76
                           );
   U77 : XOR2_X1 port map( A => CARRYB_31_3_port, B => SUMB_31_4_port, Z => n77
                           );
   U78 : XOR2_X1 port map( A => CARRYB_31_7_port, B => SUMB_31_8_port, Z => n78
                           );
   U79 : XOR2_X1 port map( A => CARRYB_31_9_port, B => SUMB_31_10_port, Z => 
                           n79);
   U80 : XOR2_X1 port map( A => CARRYB_31_15_port, B => SUMB_31_16_port, Z => 
                           n80);
   U81 : XOR2_X1 port map( A => CARRYB_31_17_port, B => SUMB_31_18_port, Z => 
                           n81);
   U82 : AND2_X1 port map( A1 => CARRYB_31_4_port, A2 => SUMB_31_5_port, ZN => 
                           n82);
   U83 : AND2_X1 port map( A1 => CARRYB_31_1_port, A2 => SUMB_31_2_port, ZN => 
                           n83);
   U84 : AND2_X1 port map( A1 => CARRYB_31_5_port, A2 => SUMB_31_6_port, ZN => 
                           n84);
   U85 : AND2_X1 port map( A1 => CARRYB_31_10_port, A2 => SUMB_31_11_port, ZN 
                           => n85);
   U86 : AND2_X1 port map( A1 => CARRYB_31_9_port, A2 => SUMB_31_10_port, ZN =>
                           n86);
   U87 : AND2_X1 port map( A1 => CARRYB_31_12_port, A2 => SUMB_31_13_port, ZN 
                           => n87);
   U88 : AND2_X1 port map( A1 => CARRYB_31_17_port, A2 => SUMB_31_18_port, ZN 
                           => n88);
   U89 : AND2_X1 port map( A1 => CARRYB_31_19_port, A2 => SUMB_31_20_port, ZN 
                           => n89);
   U90 : AND2_X1 port map( A1 => CARRYB_31_21_port, A2 => SUMB_31_22_port, ZN 
                           => n90);
   U91 : AND2_X1 port map( A1 => CARRYB_31_23_port, A2 => SUMB_31_24_port, ZN 
                           => n91);
   U92 : AND2_X1 port map( A1 => CARRYB_31_25_port, A2 => SUMB_31_26_port, ZN 
                           => n92);
   U93 : AND2_X1 port map( A1 => CARRYB_31_27_port, A2 => SUMB_31_28_port, ZN 
                           => n93);
   U94 : AND2_X1 port map( A1 => CARRYB_31_0_port, A2 => SUMB_31_1_port, ZN => 
                           n94);
   U95 : AND2_X1 port map( A1 => CARRYB_31_2_port, A2 => SUMB_31_3_port, ZN => 
                           n95);
   U96 : AND2_X1 port map( A1 => CARRYB_31_6_port, A2 => SUMB_31_7_port, ZN => 
                           n96);
   U97 : AND2_X1 port map( A1 => CARRYB_31_8_port, A2 => SUMB_31_9_port, ZN => 
                           n97);
   U98 : AND2_X1 port map( A1 => CARRYB_31_14_port, A2 => SUMB_31_15_port, ZN 
                           => n98);
   U99 : AND2_X1 port map( A1 => CARRYB_31_16_port, A2 => SUMB_31_17_port, ZN 
                           => n99);
   U100 : AND2_X1 port map( A1 => CARRYB_31_29_port, A2 => SUMB_31_30_port, ZN 
                           => n100);
   U101 : XOR2_X1 port map( A => CARRYB_31_4_port, B => SUMB_31_5_port, Z => 
                           n101);
   U102 : XOR2_X1 port map( A => CARRYB_31_12_port, B => SUMB_31_13_port, Z => 
                           n102);
   U103 : XOR2_X1 port map( A => CARRYB_31_14_port, B => SUMB_31_15_port, Z => 
                           n103);
   U104 : XOR2_X1 port map( A => CARRYB_31_19_port, B => SUMB_31_20_port, Z => 
                           n104);
   U105 : XOR2_X1 port map( A => CARRYB_31_21_port, B => SUMB_31_22_port, Z => 
                           n105);
   U106 : XOR2_X1 port map( A => CARRYB_31_23_port, B => SUMB_31_24_port, Z => 
                           n106);
   U107 : XOR2_X1 port map( A => CARRYB_31_25_port, B => SUMB_31_26_port, Z => 
                           n107);
   U108 : XOR2_X1 port map( A => CARRYB_31_27_port, B => SUMB_31_28_port, Z => 
                           n108);
   U109 : XOR2_X1 port map( A => CARRYB_31_29_port, B => SUMB_31_30_port, Z => 
                           n109);
   U110 : XOR2_X1 port map( A => CARRYB_31_8_port, B => SUMB_31_9_port, Z => 
                           n110);
   U111 : XOR2_X1 port map( A => CARRYB_31_16_port, B => SUMB_31_17_port, Z => 
                           n111);
   U112 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1)
                           );
   U113 : AND2_X1 port map( A1 => CARRYB_31_3_port, A2 => SUMB_31_4_port, ZN =>
                           n113);
   U114 : AND2_X1 port map( A1 => CARRYB_31_11_port, A2 => SUMB_31_12_port, ZN 
                           => n114);
   U115 : AND2_X1 port map( A1 => CARRYB_31_13_port, A2 => SUMB_31_14_port, ZN 
                           => n115);
   U116 : AND2_X1 port map( A1 => CARRYB_31_18_port, A2 => SUMB_31_19_port, ZN 
                           => n116);
   U117 : AND2_X1 port map( A1 => CARRYB_31_20_port, A2 => SUMB_31_21_port, ZN 
                           => n117);
   U118 : AND2_X1 port map( A1 => CARRYB_31_22_port, A2 => SUMB_31_23_port, ZN 
                           => n118);
   U119 : AND2_X1 port map( A1 => CARRYB_31_24_port, A2 => SUMB_31_25_port, ZN 
                           => n119);
   U120 : AND2_X1 port map( A1 => CARRYB_31_26_port, A2 => SUMB_31_27_port, ZN 
                           => n120);
   U121 : AND2_X1 port map( A1 => CARRYB_31_28_port, A2 => SUMB_31_29_port, ZN 
                           => n121);
   U122 : AND2_X1 port map( A1 => CARRYB_31_7_port, A2 => SUMB_31_8_port, ZN =>
                           n122);
   U123 : AND2_X1 port map( A1 => CARRYB_31_15_port, A2 => SUMB_31_16_port, ZN 
                           => n123);
   U124 : AND2_X1 port map( A1 => CARRYB_31_30_port, A2 => ab_31_31_port, ZN =>
                           n124);
   U125 : XOR2_X1 port map( A => CARRYB_31_0_port, B => SUMB_31_1_port, Z => 
                           n125);
   U126 : INV_X2 port map( A => A(31), ZN => n126);
   U127 : INV_X2 port map( A => A(30), ZN => n127);
   U128 : INV_X2 port map( A => A(29), ZN => n128);
   U129 : INV_X2 port map( A => A(28), ZN => n129);
   U130 : INV_X2 port map( A => A(27), ZN => n130);
   U131 : INV_X2 port map( A => A(26), ZN => n131);
   U132 : INV_X2 port map( A => A(25), ZN => n132);
   U133 : INV_X2 port map( A => A(24), ZN => n133);
   U134 : INV_X2 port map( A => A(23), ZN => n134);
   U135 : INV_X2 port map( A => A(22), ZN => n135);
   U136 : INV_X2 port map( A => A(21), ZN => n136);
   U137 : INV_X2 port map( A => A(20), ZN => n137);
   U138 : INV_X2 port map( A => A(19), ZN => n138);
   U139 : INV_X2 port map( A => A(18), ZN => n139);
   U140 : INV_X2 port map( A => A(17), ZN => n140);
   U141 : INV_X2 port map( A => A(16), ZN => n141);
   U142 : INV_X2 port map( A => A(15), ZN => n142);
   U143 : INV_X2 port map( A => A(14), ZN => n143);
   U144 : INV_X2 port map( A => A(13), ZN => n144);
   U145 : INV_X2 port map( A => A(12), ZN => n145);
   U146 : INV_X2 port map( A => A(11), ZN => n146);
   U147 : INV_X2 port map( A => A(10), ZN => n147);
   U148 : INV_X2 port map( A => A(9), ZN => n148);
   U149 : INV_X2 port map( A => A(8), ZN => n149);
   U150 : INV_X2 port map( A => A(7), ZN => n150);
   U151 : INV_X2 port map( A => A(6), ZN => n151);
   U152 : INV_X2 port map( A => A(5), ZN => n152);
   U153 : INV_X2 port map( A => A(4), ZN => n153);
   U154 : INV_X2 port map( A => A(3), ZN => n154);
   U155 : INV_X2 port map( A => A(2), ZN => n155);
   U156 : INV_X2 port map( A => A(1), ZN => n156);
   U157 : INV_X2 port map( A => A(0), ZN => n157);
   U158 : INV_X2 port map( A => B(31), ZN => n158);
   U159 : INV_X2 port map( A => B(30), ZN => n159);
   U160 : INV_X2 port map( A => B(29), ZN => n160);
   U161 : INV_X2 port map( A => B(28), ZN => n161);
   U162 : INV_X2 port map( A => B(27), ZN => n162);
   U163 : INV_X2 port map( A => B(26), ZN => n163);
   U164 : INV_X2 port map( A => B(25), ZN => n164);
   U165 : INV_X2 port map( A => B(24), ZN => n165);
   U166 : INV_X2 port map( A => B(23), ZN => n166);
   U167 : INV_X2 port map( A => B(22), ZN => n167);
   U168 : INV_X2 port map( A => B(21), ZN => n168);
   U169 : INV_X2 port map( A => B(20), ZN => n169);
   U170 : INV_X2 port map( A => B(19), ZN => n170);
   U171 : INV_X2 port map( A => B(18), ZN => n171);
   U172 : INV_X2 port map( A => B(17), ZN => n172);
   U173 : INV_X2 port map( A => B(16), ZN => n173);
   U174 : INV_X2 port map( A => B(15), ZN => n174);
   U175 : INV_X2 port map( A => B(14), ZN => n175);
   U176 : INV_X2 port map( A => B(13), ZN => n176);
   U177 : INV_X2 port map( A => B(12), ZN => n177);
   U178 : INV_X2 port map( A => B(11), ZN => n178);
   U179 : INV_X2 port map( A => B(10), ZN => n179);
   U180 : INV_X2 port map( A => B(9), ZN => n180);
   U181 : INV_X2 port map( A => B(8), ZN => n181);
   U182 : INV_X2 port map( A => B(7), ZN => n182);
   U183 : INV_X2 port map( A => B(6), ZN => n183);
   U184 : INV_X2 port map( A => B(5), ZN => n184);
   U185 : INV_X2 port map( A => B(4), ZN => n185);
   U186 : INV_X2 port map( A => B(3), ZN => n186);
   U187 : INV_X2 port map( A => B(2), ZN => n187);
   U188 : INV_X2 port map( A => B(1), ZN => n188);
   U189 : INV_X2 port map( A => B(0), ZN => n189);
   n190 <= '0';
   U191 : NOR2_X1 port map( A1 => n148, A2 => n180, ZN => ab_9_9_port);
   U192 : NOR2_X1 port map( A1 => n148, A2 => n181, ZN => ab_9_8_port);
   U193 : NOR2_X1 port map( A1 => n148, A2 => n182, ZN => ab_9_7_port);
   U194 : NOR2_X1 port map( A1 => n148, A2 => n183, ZN => ab_9_6_port);
   U195 : NOR2_X1 port map( A1 => n148, A2 => n184, ZN => ab_9_5_port);
   U196 : NOR2_X1 port map( A1 => n148, A2 => n185, ZN => ab_9_4_port);
   U197 : NOR2_X1 port map( A1 => n148, A2 => n186, ZN => ab_9_3_port);
   U198 : NOR2_X1 port map( A1 => n148, A2 => n158, ZN => ab_9_31_port);
   U199 : NOR2_X1 port map( A1 => n148, A2 => n159, ZN => ab_9_30_port);
   U200 : NOR2_X1 port map( A1 => n148, A2 => n187, ZN => ab_9_2_port);
   U201 : NOR2_X1 port map( A1 => n148, A2 => n160, ZN => ab_9_29_port);
   U202 : NOR2_X1 port map( A1 => n148, A2 => n161, ZN => ab_9_28_port);
   U203 : NOR2_X1 port map( A1 => n148, A2 => n162, ZN => ab_9_27_port);
   U204 : NOR2_X1 port map( A1 => n148, A2 => n163, ZN => ab_9_26_port);
   U205 : NOR2_X1 port map( A1 => n148, A2 => n164, ZN => ab_9_25_port);
   U206 : NOR2_X1 port map( A1 => n148, A2 => n165, ZN => ab_9_24_port);
   U207 : NOR2_X1 port map( A1 => n148, A2 => n166, ZN => ab_9_23_port);
   U208 : NOR2_X1 port map( A1 => n148, A2 => n167, ZN => ab_9_22_port);
   U209 : NOR2_X1 port map( A1 => n148, A2 => n168, ZN => ab_9_21_port);
   U210 : NOR2_X1 port map( A1 => n148, A2 => n169, ZN => ab_9_20_port);
   U211 : NOR2_X1 port map( A1 => n148, A2 => n188, ZN => ab_9_1_port);
   U212 : NOR2_X1 port map( A1 => n148, A2 => n170, ZN => ab_9_19_port);
   U213 : NOR2_X1 port map( A1 => n148, A2 => n171, ZN => ab_9_18_port);
   U214 : NOR2_X1 port map( A1 => n148, A2 => n172, ZN => ab_9_17_port);
   U215 : NOR2_X1 port map( A1 => n148, A2 => n173, ZN => ab_9_16_port);
   U216 : NOR2_X1 port map( A1 => n148, A2 => n174, ZN => ab_9_15_port);
   U217 : NOR2_X1 port map( A1 => n148, A2 => n175, ZN => ab_9_14_port);
   U218 : NOR2_X1 port map( A1 => n148, A2 => n176, ZN => ab_9_13_port);
   U219 : NOR2_X1 port map( A1 => n148, A2 => n177, ZN => ab_9_12_port);
   U220 : NOR2_X1 port map( A1 => n148, A2 => n178, ZN => ab_9_11_port);
   U221 : NOR2_X1 port map( A1 => n148, A2 => n179, ZN => ab_9_10_port);
   U222 : NOR2_X1 port map( A1 => n148, A2 => n189, ZN => ab_9_0_port);
   U223 : NOR2_X1 port map( A1 => n180, A2 => n149, ZN => ab_8_9_port);
   U224 : NOR2_X1 port map( A1 => n181, A2 => n149, ZN => ab_8_8_port);
   U225 : NOR2_X1 port map( A1 => n182, A2 => n149, ZN => ab_8_7_port);
   U226 : NOR2_X1 port map( A1 => n183, A2 => n149, ZN => ab_8_6_port);
   U227 : NOR2_X1 port map( A1 => n184, A2 => n149, ZN => ab_8_5_port);
   U228 : NOR2_X1 port map( A1 => n185, A2 => n149, ZN => ab_8_4_port);
   U229 : NOR2_X1 port map( A1 => n186, A2 => n149, ZN => ab_8_3_port);
   U230 : NOR2_X1 port map( A1 => n158, A2 => n149, ZN => ab_8_31_port);
   U231 : NOR2_X1 port map( A1 => n159, A2 => n149, ZN => ab_8_30_port);
   U232 : NOR2_X1 port map( A1 => n187, A2 => n149, ZN => ab_8_2_port);
   U233 : NOR2_X1 port map( A1 => n160, A2 => n149, ZN => ab_8_29_port);
   U234 : NOR2_X1 port map( A1 => n161, A2 => n149, ZN => ab_8_28_port);
   U235 : NOR2_X1 port map( A1 => n162, A2 => n149, ZN => ab_8_27_port);
   U236 : NOR2_X1 port map( A1 => n163, A2 => n149, ZN => ab_8_26_port);
   U237 : NOR2_X1 port map( A1 => n164, A2 => n149, ZN => ab_8_25_port);
   U238 : NOR2_X1 port map( A1 => n165, A2 => n149, ZN => ab_8_24_port);
   U239 : NOR2_X1 port map( A1 => n166, A2 => n149, ZN => ab_8_23_port);
   U240 : NOR2_X1 port map( A1 => n167, A2 => n149, ZN => ab_8_22_port);
   U241 : NOR2_X1 port map( A1 => n168, A2 => n149, ZN => ab_8_21_port);
   U242 : NOR2_X1 port map( A1 => n169, A2 => n149, ZN => ab_8_20_port);
   U243 : NOR2_X1 port map( A1 => n188, A2 => n149, ZN => ab_8_1_port);
   U244 : NOR2_X1 port map( A1 => n170, A2 => n149, ZN => ab_8_19_port);
   U245 : NOR2_X1 port map( A1 => n171, A2 => n149, ZN => ab_8_18_port);
   U246 : NOR2_X1 port map( A1 => n172, A2 => n149, ZN => ab_8_17_port);
   U247 : NOR2_X1 port map( A1 => n173, A2 => n149, ZN => ab_8_16_port);
   U248 : NOR2_X1 port map( A1 => n174, A2 => n149, ZN => ab_8_15_port);
   U249 : NOR2_X1 port map( A1 => n175, A2 => n149, ZN => ab_8_14_port);
   U250 : NOR2_X1 port map( A1 => n176, A2 => n149, ZN => ab_8_13_port);
   U251 : NOR2_X1 port map( A1 => n177, A2 => n149, ZN => ab_8_12_port);
   U252 : NOR2_X1 port map( A1 => n178, A2 => n149, ZN => ab_8_11_port);
   U253 : NOR2_X1 port map( A1 => n179, A2 => n149, ZN => ab_8_10_port);
   U254 : NOR2_X1 port map( A1 => n189, A2 => n149, ZN => ab_8_0_port);
   U255 : NOR2_X1 port map( A1 => n180, A2 => n150, ZN => ab_7_9_port);
   U256 : NOR2_X1 port map( A1 => n181, A2 => n150, ZN => ab_7_8_port);
   U257 : NOR2_X1 port map( A1 => n182, A2 => n150, ZN => ab_7_7_port);
   U258 : NOR2_X1 port map( A1 => n183, A2 => n150, ZN => ab_7_6_port);
   U259 : NOR2_X1 port map( A1 => n184, A2 => n150, ZN => ab_7_5_port);
   U260 : NOR2_X1 port map( A1 => n185, A2 => n150, ZN => ab_7_4_port);
   U261 : NOR2_X1 port map( A1 => n186, A2 => n150, ZN => ab_7_3_port);
   U262 : NOR2_X1 port map( A1 => n158, A2 => n150, ZN => ab_7_31_port);
   U263 : NOR2_X1 port map( A1 => n159, A2 => n150, ZN => ab_7_30_port);
   U264 : NOR2_X1 port map( A1 => n187, A2 => n150, ZN => ab_7_2_port);
   U265 : NOR2_X1 port map( A1 => n160, A2 => n150, ZN => ab_7_29_port);
   U266 : NOR2_X1 port map( A1 => n161, A2 => n150, ZN => ab_7_28_port);
   U267 : NOR2_X1 port map( A1 => n162, A2 => n150, ZN => ab_7_27_port);
   U268 : NOR2_X1 port map( A1 => n163, A2 => n150, ZN => ab_7_26_port);
   U269 : NOR2_X1 port map( A1 => n164, A2 => n150, ZN => ab_7_25_port);
   U270 : NOR2_X1 port map( A1 => n165, A2 => n150, ZN => ab_7_24_port);
   U271 : NOR2_X1 port map( A1 => n166, A2 => n150, ZN => ab_7_23_port);
   U272 : NOR2_X1 port map( A1 => n167, A2 => n150, ZN => ab_7_22_port);
   U273 : NOR2_X1 port map( A1 => n168, A2 => n150, ZN => ab_7_21_port);
   U274 : NOR2_X1 port map( A1 => n169, A2 => n150, ZN => ab_7_20_port);
   U275 : NOR2_X1 port map( A1 => n188, A2 => n150, ZN => ab_7_1_port);
   U276 : NOR2_X1 port map( A1 => n170, A2 => n150, ZN => ab_7_19_port);
   U277 : NOR2_X1 port map( A1 => n171, A2 => n150, ZN => ab_7_18_port);
   U278 : NOR2_X1 port map( A1 => n172, A2 => n150, ZN => ab_7_17_port);
   U279 : NOR2_X1 port map( A1 => n173, A2 => n150, ZN => ab_7_16_port);
   U280 : NOR2_X1 port map( A1 => n174, A2 => n150, ZN => ab_7_15_port);
   U281 : NOR2_X1 port map( A1 => n175, A2 => n150, ZN => ab_7_14_port);
   U282 : NOR2_X1 port map( A1 => n176, A2 => n150, ZN => ab_7_13_port);
   U283 : NOR2_X1 port map( A1 => n177, A2 => n150, ZN => ab_7_12_port);
   U284 : NOR2_X1 port map( A1 => n178, A2 => n150, ZN => ab_7_11_port);
   U285 : NOR2_X1 port map( A1 => n179, A2 => n150, ZN => ab_7_10_port);
   U286 : NOR2_X1 port map( A1 => n189, A2 => n150, ZN => ab_7_0_port);
   U287 : NOR2_X1 port map( A1 => n180, A2 => n151, ZN => ab_6_9_port);
   U288 : NOR2_X1 port map( A1 => n181, A2 => n151, ZN => ab_6_8_port);
   U289 : NOR2_X1 port map( A1 => n182, A2 => n151, ZN => ab_6_7_port);
   U290 : NOR2_X1 port map( A1 => n183, A2 => n151, ZN => ab_6_6_port);
   U291 : NOR2_X1 port map( A1 => n184, A2 => n151, ZN => ab_6_5_port);
   U292 : NOR2_X1 port map( A1 => n185, A2 => n151, ZN => ab_6_4_port);
   U293 : NOR2_X1 port map( A1 => n186, A2 => n151, ZN => ab_6_3_port);
   U294 : NOR2_X1 port map( A1 => n158, A2 => n151, ZN => ab_6_31_port);
   U295 : NOR2_X1 port map( A1 => n159, A2 => n151, ZN => ab_6_30_port);
   U296 : NOR2_X1 port map( A1 => n187, A2 => n151, ZN => ab_6_2_port);
   U297 : NOR2_X1 port map( A1 => n160, A2 => n151, ZN => ab_6_29_port);
   U298 : NOR2_X1 port map( A1 => n161, A2 => n151, ZN => ab_6_28_port);
   U299 : NOR2_X1 port map( A1 => n162, A2 => n151, ZN => ab_6_27_port);
   U300 : NOR2_X1 port map( A1 => n163, A2 => n151, ZN => ab_6_26_port);
   U301 : NOR2_X1 port map( A1 => n164, A2 => n151, ZN => ab_6_25_port);
   U302 : NOR2_X1 port map( A1 => n165, A2 => n151, ZN => ab_6_24_port);
   U303 : NOR2_X1 port map( A1 => n166, A2 => n151, ZN => ab_6_23_port);
   U304 : NOR2_X1 port map( A1 => n167, A2 => n151, ZN => ab_6_22_port);
   U305 : NOR2_X1 port map( A1 => n168, A2 => n151, ZN => ab_6_21_port);
   U306 : NOR2_X1 port map( A1 => n169, A2 => n151, ZN => ab_6_20_port);
   U307 : NOR2_X1 port map( A1 => n188, A2 => n151, ZN => ab_6_1_port);
   U308 : NOR2_X1 port map( A1 => n170, A2 => n151, ZN => ab_6_19_port);
   U309 : NOR2_X1 port map( A1 => n171, A2 => n151, ZN => ab_6_18_port);
   U310 : NOR2_X1 port map( A1 => n172, A2 => n151, ZN => ab_6_17_port);
   U311 : NOR2_X1 port map( A1 => n173, A2 => n151, ZN => ab_6_16_port);
   U312 : NOR2_X1 port map( A1 => n174, A2 => n151, ZN => ab_6_15_port);
   U313 : NOR2_X1 port map( A1 => n175, A2 => n151, ZN => ab_6_14_port);
   U314 : NOR2_X1 port map( A1 => n176, A2 => n151, ZN => ab_6_13_port);
   U315 : NOR2_X1 port map( A1 => n177, A2 => n151, ZN => ab_6_12_port);
   U316 : NOR2_X1 port map( A1 => n178, A2 => n151, ZN => ab_6_11_port);
   U317 : NOR2_X1 port map( A1 => n179, A2 => n151, ZN => ab_6_10_port);
   U318 : NOR2_X1 port map( A1 => n189, A2 => n151, ZN => ab_6_0_port);
   U319 : NOR2_X1 port map( A1 => n180, A2 => n152, ZN => ab_5_9_port);
   U320 : NOR2_X1 port map( A1 => n181, A2 => n152, ZN => ab_5_8_port);
   U321 : NOR2_X1 port map( A1 => n182, A2 => n152, ZN => ab_5_7_port);
   U322 : NOR2_X1 port map( A1 => n183, A2 => n152, ZN => ab_5_6_port);
   U323 : NOR2_X1 port map( A1 => n184, A2 => n152, ZN => ab_5_5_port);
   U324 : NOR2_X1 port map( A1 => n185, A2 => n152, ZN => ab_5_4_port);
   U325 : NOR2_X1 port map( A1 => n186, A2 => n152, ZN => ab_5_3_port);
   U326 : NOR2_X1 port map( A1 => n158, A2 => n152, ZN => ab_5_31_port);
   U327 : NOR2_X1 port map( A1 => n159, A2 => n152, ZN => ab_5_30_port);
   U328 : NOR2_X1 port map( A1 => n187, A2 => n152, ZN => ab_5_2_port);
   U329 : NOR2_X1 port map( A1 => n160, A2 => n152, ZN => ab_5_29_port);
   U330 : NOR2_X1 port map( A1 => n161, A2 => n152, ZN => ab_5_28_port);
   U331 : NOR2_X1 port map( A1 => n162, A2 => n152, ZN => ab_5_27_port);
   U332 : NOR2_X1 port map( A1 => n163, A2 => n152, ZN => ab_5_26_port);
   U333 : NOR2_X1 port map( A1 => n164, A2 => n152, ZN => ab_5_25_port);
   U334 : NOR2_X1 port map( A1 => n165, A2 => n152, ZN => ab_5_24_port);
   U335 : NOR2_X1 port map( A1 => n166, A2 => n152, ZN => ab_5_23_port);
   U336 : NOR2_X1 port map( A1 => n167, A2 => n152, ZN => ab_5_22_port);
   U337 : NOR2_X1 port map( A1 => n168, A2 => n152, ZN => ab_5_21_port);
   U338 : NOR2_X1 port map( A1 => n169, A2 => n152, ZN => ab_5_20_port);
   U339 : NOR2_X1 port map( A1 => n188, A2 => n152, ZN => ab_5_1_port);
   U340 : NOR2_X1 port map( A1 => n170, A2 => n152, ZN => ab_5_19_port);
   U341 : NOR2_X1 port map( A1 => n171, A2 => n152, ZN => ab_5_18_port);
   U342 : NOR2_X1 port map( A1 => n172, A2 => n152, ZN => ab_5_17_port);
   U343 : NOR2_X1 port map( A1 => n173, A2 => n152, ZN => ab_5_16_port);
   U344 : NOR2_X1 port map( A1 => n174, A2 => n152, ZN => ab_5_15_port);
   U345 : NOR2_X1 port map( A1 => n175, A2 => n152, ZN => ab_5_14_port);
   U346 : NOR2_X1 port map( A1 => n176, A2 => n152, ZN => ab_5_13_port);
   U347 : NOR2_X1 port map( A1 => n177, A2 => n152, ZN => ab_5_12_port);
   U348 : NOR2_X1 port map( A1 => n178, A2 => n152, ZN => ab_5_11_port);
   U349 : NOR2_X1 port map( A1 => n179, A2 => n152, ZN => ab_5_10_port);
   U350 : NOR2_X1 port map( A1 => n189, A2 => n152, ZN => ab_5_0_port);
   U351 : NOR2_X1 port map( A1 => n180, A2 => n153, ZN => ab_4_9_port);
   U352 : NOR2_X1 port map( A1 => n181, A2 => n153, ZN => ab_4_8_port);
   U353 : NOR2_X1 port map( A1 => n182, A2 => n153, ZN => ab_4_7_port);
   U354 : NOR2_X1 port map( A1 => n183, A2 => n153, ZN => ab_4_6_port);
   U355 : NOR2_X1 port map( A1 => n184, A2 => n153, ZN => ab_4_5_port);
   U356 : NOR2_X1 port map( A1 => n185, A2 => n153, ZN => ab_4_4_port);
   U357 : NOR2_X1 port map( A1 => n186, A2 => n153, ZN => ab_4_3_port);
   U358 : NOR2_X1 port map( A1 => n158, A2 => n153, ZN => ab_4_31_port);
   U359 : NOR2_X1 port map( A1 => n159, A2 => n153, ZN => ab_4_30_port);
   U360 : NOR2_X1 port map( A1 => n187, A2 => n153, ZN => ab_4_2_port);
   U361 : NOR2_X1 port map( A1 => n160, A2 => n153, ZN => ab_4_29_port);
   U362 : NOR2_X1 port map( A1 => n161, A2 => n153, ZN => ab_4_28_port);
   U363 : NOR2_X1 port map( A1 => n162, A2 => n153, ZN => ab_4_27_port);
   U364 : NOR2_X1 port map( A1 => n163, A2 => n153, ZN => ab_4_26_port);
   U365 : NOR2_X1 port map( A1 => n164, A2 => n153, ZN => ab_4_25_port);
   U366 : NOR2_X1 port map( A1 => n165, A2 => n153, ZN => ab_4_24_port);
   U367 : NOR2_X1 port map( A1 => n166, A2 => n153, ZN => ab_4_23_port);
   U368 : NOR2_X1 port map( A1 => n167, A2 => n153, ZN => ab_4_22_port);
   U369 : NOR2_X1 port map( A1 => n168, A2 => n153, ZN => ab_4_21_port);
   U370 : NOR2_X1 port map( A1 => n169, A2 => n153, ZN => ab_4_20_port);
   U371 : NOR2_X1 port map( A1 => n188, A2 => n153, ZN => ab_4_1_port);
   U372 : NOR2_X1 port map( A1 => n170, A2 => n153, ZN => ab_4_19_port);
   U373 : NOR2_X1 port map( A1 => n171, A2 => n153, ZN => ab_4_18_port);
   U374 : NOR2_X1 port map( A1 => n172, A2 => n153, ZN => ab_4_17_port);
   U375 : NOR2_X1 port map( A1 => n173, A2 => n153, ZN => ab_4_16_port);
   U376 : NOR2_X1 port map( A1 => n174, A2 => n153, ZN => ab_4_15_port);
   U377 : NOR2_X1 port map( A1 => n175, A2 => n153, ZN => ab_4_14_port);
   U378 : NOR2_X1 port map( A1 => n176, A2 => n153, ZN => ab_4_13_port);
   U379 : NOR2_X1 port map( A1 => n177, A2 => n153, ZN => ab_4_12_port);
   U380 : NOR2_X1 port map( A1 => n178, A2 => n153, ZN => ab_4_11_port);
   U381 : NOR2_X1 port map( A1 => n179, A2 => n153, ZN => ab_4_10_port);
   U382 : NOR2_X1 port map( A1 => n189, A2 => n153, ZN => ab_4_0_port);
   U383 : NOR2_X1 port map( A1 => n180, A2 => n154, ZN => ab_3_9_port);
   U384 : NOR2_X1 port map( A1 => n181, A2 => n154, ZN => ab_3_8_port);
   U385 : NOR2_X1 port map( A1 => n182, A2 => n154, ZN => ab_3_7_port);
   U386 : NOR2_X1 port map( A1 => n183, A2 => n154, ZN => ab_3_6_port);
   U387 : NOR2_X1 port map( A1 => n184, A2 => n154, ZN => ab_3_5_port);
   U388 : NOR2_X1 port map( A1 => n185, A2 => n154, ZN => ab_3_4_port);
   U389 : NOR2_X1 port map( A1 => n186, A2 => n154, ZN => ab_3_3_port);
   U390 : NOR2_X1 port map( A1 => n158, A2 => n154, ZN => ab_3_31_port);
   U391 : NOR2_X1 port map( A1 => n159, A2 => n154, ZN => ab_3_30_port);
   U392 : NOR2_X1 port map( A1 => n187, A2 => n154, ZN => ab_3_2_port);
   U393 : NOR2_X1 port map( A1 => n160, A2 => n154, ZN => ab_3_29_port);
   U394 : NOR2_X1 port map( A1 => n161, A2 => n154, ZN => ab_3_28_port);
   U395 : NOR2_X1 port map( A1 => n162, A2 => n154, ZN => ab_3_27_port);
   U396 : NOR2_X1 port map( A1 => n163, A2 => n154, ZN => ab_3_26_port);
   U397 : NOR2_X1 port map( A1 => n164, A2 => n154, ZN => ab_3_25_port);
   U398 : NOR2_X1 port map( A1 => n165, A2 => n154, ZN => ab_3_24_port);
   U399 : NOR2_X1 port map( A1 => n166, A2 => n154, ZN => ab_3_23_port);
   U400 : NOR2_X1 port map( A1 => n167, A2 => n154, ZN => ab_3_22_port);
   U401 : NOR2_X1 port map( A1 => n168, A2 => n154, ZN => ab_3_21_port);
   U402 : NOR2_X1 port map( A1 => n169, A2 => n154, ZN => ab_3_20_port);
   U403 : NOR2_X1 port map( A1 => n188, A2 => n154, ZN => ab_3_1_port);
   U404 : NOR2_X1 port map( A1 => n170, A2 => n154, ZN => ab_3_19_port);
   U405 : NOR2_X1 port map( A1 => n171, A2 => n154, ZN => ab_3_18_port);
   U406 : NOR2_X1 port map( A1 => n172, A2 => n154, ZN => ab_3_17_port);
   U407 : NOR2_X1 port map( A1 => n173, A2 => n154, ZN => ab_3_16_port);
   U408 : NOR2_X1 port map( A1 => n174, A2 => n154, ZN => ab_3_15_port);
   U409 : NOR2_X1 port map( A1 => n175, A2 => n154, ZN => ab_3_14_port);
   U410 : NOR2_X1 port map( A1 => n176, A2 => n154, ZN => ab_3_13_port);
   U411 : NOR2_X1 port map( A1 => n177, A2 => n154, ZN => ab_3_12_port);
   U412 : NOR2_X1 port map( A1 => n178, A2 => n154, ZN => ab_3_11_port);
   U413 : NOR2_X1 port map( A1 => n179, A2 => n154, ZN => ab_3_10_port);
   U414 : NOR2_X1 port map( A1 => n189, A2 => n154, ZN => ab_3_0_port);
   U415 : NOR2_X1 port map( A1 => n180, A2 => n126, ZN => ab_31_9_port);
   U416 : NOR2_X1 port map( A1 => n181, A2 => n126, ZN => ab_31_8_port);
   U417 : NOR2_X1 port map( A1 => n182, A2 => n126, ZN => ab_31_7_port);
   U418 : NOR2_X1 port map( A1 => n183, A2 => n126, ZN => ab_31_6_port);
   U419 : NOR2_X1 port map( A1 => n184, A2 => n126, ZN => ab_31_5_port);
   U420 : NOR2_X1 port map( A1 => n185, A2 => n126, ZN => ab_31_4_port);
   U421 : NOR2_X1 port map( A1 => n186, A2 => n126, ZN => ab_31_3_port);
   U422 : NOR2_X1 port map( A1 => n158, A2 => n126, ZN => ab_31_31_port);
   U423 : NOR2_X1 port map( A1 => n159, A2 => n126, ZN => ab_31_30_port);
   U424 : NOR2_X1 port map( A1 => n187, A2 => n126, ZN => ab_31_2_port);
   U425 : NOR2_X1 port map( A1 => n160, A2 => n126, ZN => ab_31_29_port);
   U426 : NOR2_X1 port map( A1 => n161, A2 => n126, ZN => ab_31_28_port);
   U427 : NOR2_X1 port map( A1 => n162, A2 => n126, ZN => ab_31_27_port);
   U428 : NOR2_X1 port map( A1 => n163, A2 => n126, ZN => ab_31_26_port);
   U429 : NOR2_X1 port map( A1 => n164, A2 => n126, ZN => ab_31_25_port);
   U430 : NOR2_X1 port map( A1 => n165, A2 => n126, ZN => ab_31_24_port);
   U431 : NOR2_X1 port map( A1 => n166, A2 => n126, ZN => ab_31_23_port);
   U432 : NOR2_X1 port map( A1 => n167, A2 => n126, ZN => ab_31_22_port);
   U433 : NOR2_X1 port map( A1 => n168, A2 => n126, ZN => ab_31_21_port);
   U434 : NOR2_X1 port map( A1 => n169, A2 => n126, ZN => ab_31_20_port);
   U435 : NOR2_X1 port map( A1 => n188, A2 => n126, ZN => ab_31_1_port);
   U436 : NOR2_X1 port map( A1 => n170, A2 => n126, ZN => ab_31_19_port);
   U437 : NOR2_X1 port map( A1 => n171, A2 => n126, ZN => ab_31_18_port);
   U438 : NOR2_X1 port map( A1 => n172, A2 => n126, ZN => ab_31_17_port);
   U439 : NOR2_X1 port map( A1 => n173, A2 => n126, ZN => ab_31_16_port);
   U440 : NOR2_X1 port map( A1 => n174, A2 => n126, ZN => ab_31_15_port);
   U441 : NOR2_X1 port map( A1 => n175, A2 => n126, ZN => ab_31_14_port);
   U442 : NOR2_X1 port map( A1 => n176, A2 => n126, ZN => ab_31_13_port);
   U443 : NOR2_X1 port map( A1 => n177, A2 => n126, ZN => ab_31_12_port);
   U444 : NOR2_X1 port map( A1 => n178, A2 => n126, ZN => ab_31_11_port);
   U445 : NOR2_X1 port map( A1 => n179, A2 => n126, ZN => ab_31_10_port);
   U446 : NOR2_X1 port map( A1 => n189, A2 => n126, ZN => ab_31_0_port);
   U447 : NOR2_X1 port map( A1 => n180, A2 => n127, ZN => ab_30_9_port);
   U448 : NOR2_X1 port map( A1 => n181, A2 => n127, ZN => ab_30_8_port);
   U449 : NOR2_X1 port map( A1 => n182, A2 => n127, ZN => ab_30_7_port);
   U450 : NOR2_X1 port map( A1 => n183, A2 => n127, ZN => ab_30_6_port);
   U451 : NOR2_X1 port map( A1 => n184, A2 => n127, ZN => ab_30_5_port);
   U452 : NOR2_X1 port map( A1 => n185, A2 => n127, ZN => ab_30_4_port);
   U453 : NOR2_X1 port map( A1 => n186, A2 => n127, ZN => ab_30_3_port);
   U454 : NOR2_X1 port map( A1 => n158, A2 => n127, ZN => ab_30_31_port);
   U455 : NOR2_X1 port map( A1 => n159, A2 => n127, ZN => ab_30_30_port);
   U456 : NOR2_X1 port map( A1 => n187, A2 => n127, ZN => ab_30_2_port);
   U457 : NOR2_X1 port map( A1 => n160, A2 => n127, ZN => ab_30_29_port);
   U458 : NOR2_X1 port map( A1 => n161, A2 => n127, ZN => ab_30_28_port);
   U459 : NOR2_X1 port map( A1 => n162, A2 => n127, ZN => ab_30_27_port);
   U460 : NOR2_X1 port map( A1 => n163, A2 => n127, ZN => ab_30_26_port);
   U461 : NOR2_X1 port map( A1 => n164, A2 => n127, ZN => ab_30_25_port);
   U462 : NOR2_X1 port map( A1 => n165, A2 => n127, ZN => ab_30_24_port);
   U463 : NOR2_X1 port map( A1 => n166, A2 => n127, ZN => ab_30_23_port);
   U464 : NOR2_X1 port map( A1 => n167, A2 => n127, ZN => ab_30_22_port);
   U465 : NOR2_X1 port map( A1 => n168, A2 => n127, ZN => ab_30_21_port);
   U466 : NOR2_X1 port map( A1 => n169, A2 => n127, ZN => ab_30_20_port);
   U467 : NOR2_X1 port map( A1 => n188, A2 => n127, ZN => ab_30_1_port);
   U468 : NOR2_X1 port map( A1 => n170, A2 => n127, ZN => ab_30_19_port);
   U469 : NOR2_X1 port map( A1 => n171, A2 => n127, ZN => ab_30_18_port);
   U470 : NOR2_X1 port map( A1 => n172, A2 => n127, ZN => ab_30_17_port);
   U471 : NOR2_X1 port map( A1 => n173, A2 => n127, ZN => ab_30_16_port);
   U472 : NOR2_X1 port map( A1 => n174, A2 => n127, ZN => ab_30_15_port);
   U473 : NOR2_X1 port map( A1 => n175, A2 => n127, ZN => ab_30_14_port);
   U474 : NOR2_X1 port map( A1 => n176, A2 => n127, ZN => ab_30_13_port);
   U475 : NOR2_X1 port map( A1 => n177, A2 => n127, ZN => ab_30_12_port);
   U476 : NOR2_X1 port map( A1 => n178, A2 => n127, ZN => ab_30_11_port);
   U477 : NOR2_X1 port map( A1 => n179, A2 => n127, ZN => ab_30_10_port);
   U478 : NOR2_X1 port map( A1 => n189, A2 => n127, ZN => ab_30_0_port);
   U479 : NOR2_X1 port map( A1 => n180, A2 => n155, ZN => ab_2_9_port);
   U480 : NOR2_X1 port map( A1 => n181, A2 => n155, ZN => ab_2_8_port);
   U481 : NOR2_X1 port map( A1 => n182, A2 => n155, ZN => ab_2_7_port);
   U482 : NOR2_X1 port map( A1 => n183, A2 => n155, ZN => ab_2_6_port);
   U483 : NOR2_X1 port map( A1 => n184, A2 => n155, ZN => ab_2_5_port);
   U484 : NOR2_X1 port map( A1 => n185, A2 => n155, ZN => ab_2_4_port);
   U485 : NOR2_X1 port map( A1 => n186, A2 => n155, ZN => ab_2_3_port);
   U486 : NOR2_X1 port map( A1 => n158, A2 => n155, ZN => ab_2_31_port);
   U487 : NOR2_X1 port map( A1 => n159, A2 => n155, ZN => ab_2_30_port);
   U488 : NOR2_X1 port map( A1 => n187, A2 => n155, ZN => ab_2_2_port);
   U489 : NOR2_X1 port map( A1 => n160, A2 => n155, ZN => ab_2_29_port);
   U490 : NOR2_X1 port map( A1 => n161, A2 => n155, ZN => ab_2_28_port);
   U491 : NOR2_X1 port map( A1 => n162, A2 => n155, ZN => ab_2_27_port);
   U492 : NOR2_X1 port map( A1 => n163, A2 => n155, ZN => ab_2_26_port);
   U493 : NOR2_X1 port map( A1 => n164, A2 => n155, ZN => ab_2_25_port);
   U494 : NOR2_X1 port map( A1 => n165, A2 => n155, ZN => ab_2_24_port);
   U495 : NOR2_X1 port map( A1 => n166, A2 => n155, ZN => ab_2_23_port);
   U496 : NOR2_X1 port map( A1 => n167, A2 => n155, ZN => ab_2_22_port);
   U497 : NOR2_X1 port map( A1 => n168, A2 => n155, ZN => ab_2_21_port);
   U498 : NOR2_X1 port map( A1 => n169, A2 => n155, ZN => ab_2_20_port);
   U499 : NOR2_X1 port map( A1 => n188, A2 => n155, ZN => ab_2_1_port);
   U500 : NOR2_X1 port map( A1 => n170, A2 => n155, ZN => ab_2_19_port);
   U501 : NOR2_X1 port map( A1 => n171, A2 => n155, ZN => ab_2_18_port);
   U502 : NOR2_X1 port map( A1 => n172, A2 => n155, ZN => ab_2_17_port);
   U503 : NOR2_X1 port map( A1 => n173, A2 => n155, ZN => ab_2_16_port);
   U504 : NOR2_X1 port map( A1 => n174, A2 => n155, ZN => ab_2_15_port);
   U505 : NOR2_X1 port map( A1 => n175, A2 => n155, ZN => ab_2_14_port);
   U506 : NOR2_X1 port map( A1 => n176, A2 => n155, ZN => ab_2_13_port);
   U507 : NOR2_X1 port map( A1 => n177, A2 => n155, ZN => ab_2_12_port);
   U508 : NOR2_X1 port map( A1 => n178, A2 => n155, ZN => ab_2_11_port);
   U509 : NOR2_X1 port map( A1 => n179, A2 => n155, ZN => ab_2_10_port);
   U510 : NOR2_X1 port map( A1 => n189, A2 => n155, ZN => ab_2_0_port);
   U511 : NOR2_X1 port map( A1 => n180, A2 => n128, ZN => ab_29_9_port);
   U512 : NOR2_X1 port map( A1 => n181, A2 => n128, ZN => ab_29_8_port);
   U513 : NOR2_X1 port map( A1 => n182, A2 => n128, ZN => ab_29_7_port);
   U514 : NOR2_X1 port map( A1 => n183, A2 => n128, ZN => ab_29_6_port);
   U515 : NOR2_X1 port map( A1 => n184, A2 => n128, ZN => ab_29_5_port);
   U516 : NOR2_X1 port map( A1 => n185, A2 => n128, ZN => ab_29_4_port);
   U517 : NOR2_X1 port map( A1 => n186, A2 => n128, ZN => ab_29_3_port);
   U518 : NOR2_X1 port map( A1 => n158, A2 => n128, ZN => ab_29_31_port);
   U519 : NOR2_X1 port map( A1 => n159, A2 => n128, ZN => ab_29_30_port);
   U520 : NOR2_X1 port map( A1 => n187, A2 => n128, ZN => ab_29_2_port);
   U521 : NOR2_X1 port map( A1 => n160, A2 => n128, ZN => ab_29_29_port);
   U522 : NOR2_X1 port map( A1 => n161, A2 => n128, ZN => ab_29_28_port);
   U523 : NOR2_X1 port map( A1 => n162, A2 => n128, ZN => ab_29_27_port);
   U524 : NOR2_X1 port map( A1 => n163, A2 => n128, ZN => ab_29_26_port);
   U525 : NOR2_X1 port map( A1 => n164, A2 => n128, ZN => ab_29_25_port);
   U526 : NOR2_X1 port map( A1 => n165, A2 => n128, ZN => ab_29_24_port);
   U527 : NOR2_X1 port map( A1 => n166, A2 => n128, ZN => ab_29_23_port);
   U528 : NOR2_X1 port map( A1 => n167, A2 => n128, ZN => ab_29_22_port);
   U529 : NOR2_X1 port map( A1 => n168, A2 => n128, ZN => ab_29_21_port);
   U530 : NOR2_X1 port map( A1 => n169, A2 => n128, ZN => ab_29_20_port);
   U531 : NOR2_X1 port map( A1 => n188, A2 => n128, ZN => ab_29_1_port);
   U532 : NOR2_X1 port map( A1 => n170, A2 => n128, ZN => ab_29_19_port);
   U533 : NOR2_X1 port map( A1 => n171, A2 => n128, ZN => ab_29_18_port);
   U534 : NOR2_X1 port map( A1 => n172, A2 => n128, ZN => ab_29_17_port);
   U535 : NOR2_X1 port map( A1 => n173, A2 => n128, ZN => ab_29_16_port);
   U536 : NOR2_X1 port map( A1 => n174, A2 => n128, ZN => ab_29_15_port);
   U537 : NOR2_X1 port map( A1 => n175, A2 => n128, ZN => ab_29_14_port);
   U538 : NOR2_X1 port map( A1 => n176, A2 => n128, ZN => ab_29_13_port);
   U539 : NOR2_X1 port map( A1 => n177, A2 => n128, ZN => ab_29_12_port);
   U540 : NOR2_X1 port map( A1 => n178, A2 => n128, ZN => ab_29_11_port);
   U541 : NOR2_X1 port map( A1 => n179, A2 => n128, ZN => ab_29_10_port);
   U542 : NOR2_X1 port map( A1 => n189, A2 => n128, ZN => ab_29_0_port);
   U543 : NOR2_X1 port map( A1 => n180, A2 => n129, ZN => ab_28_9_port);
   U544 : NOR2_X1 port map( A1 => n181, A2 => n129, ZN => ab_28_8_port);
   U545 : NOR2_X1 port map( A1 => n182, A2 => n129, ZN => ab_28_7_port);
   U546 : NOR2_X1 port map( A1 => n183, A2 => n129, ZN => ab_28_6_port);
   U547 : NOR2_X1 port map( A1 => n184, A2 => n129, ZN => ab_28_5_port);
   U548 : NOR2_X1 port map( A1 => n185, A2 => n129, ZN => ab_28_4_port);
   U549 : NOR2_X1 port map( A1 => n186, A2 => n129, ZN => ab_28_3_port);
   U550 : NOR2_X1 port map( A1 => n158, A2 => n129, ZN => ab_28_31_port);
   U551 : NOR2_X1 port map( A1 => n159, A2 => n129, ZN => ab_28_30_port);
   U552 : NOR2_X1 port map( A1 => n187, A2 => n129, ZN => ab_28_2_port);
   U553 : NOR2_X1 port map( A1 => n160, A2 => n129, ZN => ab_28_29_port);
   U554 : NOR2_X1 port map( A1 => n161, A2 => n129, ZN => ab_28_28_port);
   U555 : NOR2_X1 port map( A1 => n162, A2 => n129, ZN => ab_28_27_port);
   U556 : NOR2_X1 port map( A1 => n163, A2 => n129, ZN => ab_28_26_port);
   U557 : NOR2_X1 port map( A1 => n164, A2 => n129, ZN => ab_28_25_port);
   U558 : NOR2_X1 port map( A1 => n165, A2 => n129, ZN => ab_28_24_port);
   U559 : NOR2_X1 port map( A1 => n166, A2 => n129, ZN => ab_28_23_port);
   U560 : NOR2_X1 port map( A1 => n167, A2 => n129, ZN => ab_28_22_port);
   U561 : NOR2_X1 port map( A1 => n168, A2 => n129, ZN => ab_28_21_port);
   U562 : NOR2_X1 port map( A1 => n169, A2 => n129, ZN => ab_28_20_port);
   U563 : NOR2_X1 port map( A1 => n188, A2 => n129, ZN => ab_28_1_port);
   U564 : NOR2_X1 port map( A1 => n170, A2 => n129, ZN => ab_28_19_port);
   U565 : NOR2_X1 port map( A1 => n171, A2 => n129, ZN => ab_28_18_port);
   U566 : NOR2_X1 port map( A1 => n172, A2 => n129, ZN => ab_28_17_port);
   U567 : NOR2_X1 port map( A1 => n173, A2 => n129, ZN => ab_28_16_port);
   U568 : NOR2_X1 port map( A1 => n174, A2 => n129, ZN => ab_28_15_port);
   U569 : NOR2_X1 port map( A1 => n175, A2 => n129, ZN => ab_28_14_port);
   U570 : NOR2_X1 port map( A1 => n176, A2 => n129, ZN => ab_28_13_port);
   U571 : NOR2_X1 port map( A1 => n177, A2 => n129, ZN => ab_28_12_port);
   U572 : NOR2_X1 port map( A1 => n178, A2 => n129, ZN => ab_28_11_port);
   U573 : NOR2_X1 port map( A1 => n179, A2 => n129, ZN => ab_28_10_port);
   U574 : NOR2_X1 port map( A1 => n189, A2 => n129, ZN => ab_28_0_port);
   U575 : NOR2_X1 port map( A1 => n180, A2 => n130, ZN => ab_27_9_port);
   U576 : NOR2_X1 port map( A1 => n181, A2 => n130, ZN => ab_27_8_port);
   U577 : NOR2_X1 port map( A1 => n182, A2 => n130, ZN => ab_27_7_port);
   U578 : NOR2_X1 port map( A1 => n183, A2 => n130, ZN => ab_27_6_port);
   U579 : NOR2_X1 port map( A1 => n184, A2 => n130, ZN => ab_27_5_port);
   U580 : NOR2_X1 port map( A1 => n185, A2 => n130, ZN => ab_27_4_port);
   U581 : NOR2_X1 port map( A1 => n186, A2 => n130, ZN => ab_27_3_port);
   U582 : NOR2_X1 port map( A1 => n158, A2 => n130, ZN => ab_27_31_port);
   U583 : NOR2_X1 port map( A1 => n159, A2 => n130, ZN => ab_27_30_port);
   U584 : NOR2_X1 port map( A1 => n187, A2 => n130, ZN => ab_27_2_port);
   U585 : NOR2_X1 port map( A1 => n160, A2 => n130, ZN => ab_27_29_port);
   U586 : NOR2_X1 port map( A1 => n161, A2 => n130, ZN => ab_27_28_port);
   U587 : NOR2_X1 port map( A1 => n162, A2 => n130, ZN => ab_27_27_port);
   U588 : NOR2_X1 port map( A1 => n163, A2 => n130, ZN => ab_27_26_port);
   U589 : NOR2_X1 port map( A1 => n164, A2 => n130, ZN => ab_27_25_port);
   U590 : NOR2_X1 port map( A1 => n165, A2 => n130, ZN => ab_27_24_port);
   U591 : NOR2_X1 port map( A1 => n166, A2 => n130, ZN => ab_27_23_port);
   U592 : NOR2_X1 port map( A1 => n167, A2 => n130, ZN => ab_27_22_port);
   U593 : NOR2_X1 port map( A1 => n168, A2 => n130, ZN => ab_27_21_port);
   U594 : NOR2_X1 port map( A1 => n169, A2 => n130, ZN => ab_27_20_port);
   U595 : NOR2_X1 port map( A1 => n188, A2 => n130, ZN => ab_27_1_port);
   U596 : NOR2_X1 port map( A1 => n170, A2 => n130, ZN => ab_27_19_port);
   U597 : NOR2_X1 port map( A1 => n171, A2 => n130, ZN => ab_27_18_port);
   U598 : NOR2_X1 port map( A1 => n172, A2 => n130, ZN => ab_27_17_port);
   U599 : NOR2_X1 port map( A1 => n173, A2 => n130, ZN => ab_27_16_port);
   U600 : NOR2_X1 port map( A1 => n174, A2 => n130, ZN => ab_27_15_port);
   U601 : NOR2_X1 port map( A1 => n175, A2 => n130, ZN => ab_27_14_port);
   U602 : NOR2_X1 port map( A1 => n176, A2 => n130, ZN => ab_27_13_port);
   U603 : NOR2_X1 port map( A1 => n177, A2 => n130, ZN => ab_27_12_port);
   U604 : NOR2_X1 port map( A1 => n178, A2 => n130, ZN => ab_27_11_port);
   U605 : NOR2_X1 port map( A1 => n179, A2 => n130, ZN => ab_27_10_port);
   U606 : NOR2_X1 port map( A1 => n189, A2 => n130, ZN => ab_27_0_port);
   U607 : NOR2_X1 port map( A1 => n180, A2 => n131, ZN => ab_26_9_port);
   U608 : NOR2_X1 port map( A1 => n181, A2 => n131, ZN => ab_26_8_port);
   U609 : NOR2_X1 port map( A1 => n182, A2 => n131, ZN => ab_26_7_port);
   U610 : NOR2_X1 port map( A1 => n183, A2 => n131, ZN => ab_26_6_port);
   U611 : NOR2_X1 port map( A1 => n184, A2 => n131, ZN => ab_26_5_port);
   U612 : NOR2_X1 port map( A1 => n185, A2 => n131, ZN => ab_26_4_port);
   U613 : NOR2_X1 port map( A1 => n186, A2 => n131, ZN => ab_26_3_port);
   U614 : NOR2_X1 port map( A1 => n158, A2 => n131, ZN => ab_26_31_port);
   U615 : NOR2_X1 port map( A1 => n159, A2 => n131, ZN => ab_26_30_port);
   U616 : NOR2_X1 port map( A1 => n187, A2 => n131, ZN => ab_26_2_port);
   U617 : NOR2_X1 port map( A1 => n160, A2 => n131, ZN => ab_26_29_port);
   U618 : NOR2_X1 port map( A1 => n161, A2 => n131, ZN => ab_26_28_port);
   U619 : NOR2_X1 port map( A1 => n162, A2 => n131, ZN => ab_26_27_port);
   U620 : NOR2_X1 port map( A1 => n163, A2 => n131, ZN => ab_26_26_port);
   U621 : NOR2_X1 port map( A1 => n164, A2 => n131, ZN => ab_26_25_port);
   U622 : NOR2_X1 port map( A1 => n165, A2 => n131, ZN => ab_26_24_port);
   U623 : NOR2_X1 port map( A1 => n166, A2 => n131, ZN => ab_26_23_port);
   U624 : NOR2_X1 port map( A1 => n167, A2 => n131, ZN => ab_26_22_port);
   U625 : NOR2_X1 port map( A1 => n168, A2 => n131, ZN => ab_26_21_port);
   U626 : NOR2_X1 port map( A1 => n169, A2 => n131, ZN => ab_26_20_port);
   U627 : NOR2_X1 port map( A1 => n188, A2 => n131, ZN => ab_26_1_port);
   U628 : NOR2_X1 port map( A1 => n170, A2 => n131, ZN => ab_26_19_port);
   U629 : NOR2_X1 port map( A1 => n171, A2 => n131, ZN => ab_26_18_port);
   U630 : NOR2_X1 port map( A1 => n172, A2 => n131, ZN => ab_26_17_port);
   U631 : NOR2_X1 port map( A1 => n173, A2 => n131, ZN => ab_26_16_port);
   U632 : NOR2_X1 port map( A1 => n174, A2 => n131, ZN => ab_26_15_port);
   U633 : NOR2_X1 port map( A1 => n175, A2 => n131, ZN => ab_26_14_port);
   U634 : NOR2_X1 port map( A1 => n176, A2 => n131, ZN => ab_26_13_port);
   U635 : NOR2_X1 port map( A1 => n177, A2 => n131, ZN => ab_26_12_port);
   U636 : NOR2_X1 port map( A1 => n178, A2 => n131, ZN => ab_26_11_port);
   U637 : NOR2_X1 port map( A1 => n179, A2 => n131, ZN => ab_26_10_port);
   U638 : NOR2_X1 port map( A1 => n189, A2 => n131, ZN => ab_26_0_port);
   U639 : NOR2_X1 port map( A1 => n180, A2 => n132, ZN => ab_25_9_port);
   U640 : NOR2_X1 port map( A1 => n181, A2 => n132, ZN => ab_25_8_port);
   U641 : NOR2_X1 port map( A1 => n182, A2 => n132, ZN => ab_25_7_port);
   U642 : NOR2_X1 port map( A1 => n183, A2 => n132, ZN => ab_25_6_port);
   U643 : NOR2_X1 port map( A1 => n184, A2 => n132, ZN => ab_25_5_port);
   U644 : NOR2_X1 port map( A1 => n185, A2 => n132, ZN => ab_25_4_port);
   U645 : NOR2_X1 port map( A1 => n186, A2 => n132, ZN => ab_25_3_port);
   U646 : NOR2_X1 port map( A1 => n158, A2 => n132, ZN => ab_25_31_port);
   U647 : NOR2_X1 port map( A1 => n159, A2 => n132, ZN => ab_25_30_port);
   U648 : NOR2_X1 port map( A1 => n187, A2 => n132, ZN => ab_25_2_port);
   U649 : NOR2_X1 port map( A1 => n160, A2 => n132, ZN => ab_25_29_port);
   U650 : NOR2_X1 port map( A1 => n161, A2 => n132, ZN => ab_25_28_port);
   U651 : NOR2_X1 port map( A1 => n162, A2 => n132, ZN => ab_25_27_port);
   U652 : NOR2_X1 port map( A1 => n163, A2 => n132, ZN => ab_25_26_port);
   U653 : NOR2_X1 port map( A1 => n164, A2 => n132, ZN => ab_25_25_port);
   U654 : NOR2_X1 port map( A1 => n165, A2 => n132, ZN => ab_25_24_port);
   U655 : NOR2_X1 port map( A1 => n166, A2 => n132, ZN => ab_25_23_port);
   U656 : NOR2_X1 port map( A1 => n167, A2 => n132, ZN => ab_25_22_port);
   U657 : NOR2_X1 port map( A1 => n168, A2 => n132, ZN => ab_25_21_port);
   U658 : NOR2_X1 port map( A1 => n169, A2 => n132, ZN => ab_25_20_port);
   U659 : NOR2_X1 port map( A1 => n188, A2 => n132, ZN => ab_25_1_port);
   U660 : NOR2_X1 port map( A1 => n170, A2 => n132, ZN => ab_25_19_port);
   U661 : NOR2_X1 port map( A1 => n171, A2 => n132, ZN => ab_25_18_port);
   U662 : NOR2_X1 port map( A1 => n172, A2 => n132, ZN => ab_25_17_port);
   U663 : NOR2_X1 port map( A1 => n173, A2 => n132, ZN => ab_25_16_port);
   U664 : NOR2_X1 port map( A1 => n174, A2 => n132, ZN => ab_25_15_port);
   U665 : NOR2_X1 port map( A1 => n175, A2 => n132, ZN => ab_25_14_port);
   U666 : NOR2_X1 port map( A1 => n176, A2 => n132, ZN => ab_25_13_port);
   U667 : NOR2_X1 port map( A1 => n177, A2 => n132, ZN => ab_25_12_port);
   U668 : NOR2_X1 port map( A1 => n178, A2 => n132, ZN => ab_25_11_port);
   U669 : NOR2_X1 port map( A1 => n179, A2 => n132, ZN => ab_25_10_port);
   U670 : NOR2_X1 port map( A1 => n189, A2 => n132, ZN => ab_25_0_port);
   U671 : NOR2_X1 port map( A1 => n180, A2 => n133, ZN => ab_24_9_port);
   U672 : NOR2_X1 port map( A1 => n181, A2 => n133, ZN => ab_24_8_port);
   U673 : NOR2_X1 port map( A1 => n182, A2 => n133, ZN => ab_24_7_port);
   U674 : NOR2_X1 port map( A1 => n183, A2 => n133, ZN => ab_24_6_port);
   U675 : NOR2_X1 port map( A1 => n184, A2 => n133, ZN => ab_24_5_port);
   U676 : NOR2_X1 port map( A1 => n185, A2 => n133, ZN => ab_24_4_port);
   U677 : NOR2_X1 port map( A1 => n186, A2 => n133, ZN => ab_24_3_port);
   U678 : NOR2_X1 port map( A1 => n158, A2 => n133, ZN => ab_24_31_port);
   U679 : NOR2_X1 port map( A1 => n159, A2 => n133, ZN => ab_24_30_port);
   U680 : NOR2_X1 port map( A1 => n187, A2 => n133, ZN => ab_24_2_port);
   U681 : NOR2_X1 port map( A1 => n160, A2 => n133, ZN => ab_24_29_port);
   U682 : NOR2_X1 port map( A1 => n161, A2 => n133, ZN => ab_24_28_port);
   U683 : NOR2_X1 port map( A1 => n162, A2 => n133, ZN => ab_24_27_port);
   U684 : NOR2_X1 port map( A1 => n163, A2 => n133, ZN => ab_24_26_port);
   U685 : NOR2_X1 port map( A1 => n164, A2 => n133, ZN => ab_24_25_port);
   U686 : NOR2_X1 port map( A1 => n165, A2 => n133, ZN => ab_24_24_port);
   U687 : NOR2_X1 port map( A1 => n166, A2 => n133, ZN => ab_24_23_port);
   U688 : NOR2_X1 port map( A1 => n167, A2 => n133, ZN => ab_24_22_port);
   U689 : NOR2_X1 port map( A1 => n168, A2 => n133, ZN => ab_24_21_port);
   U690 : NOR2_X1 port map( A1 => n169, A2 => n133, ZN => ab_24_20_port);
   U691 : NOR2_X1 port map( A1 => n188, A2 => n133, ZN => ab_24_1_port);
   U692 : NOR2_X1 port map( A1 => n170, A2 => n133, ZN => ab_24_19_port);
   U693 : NOR2_X1 port map( A1 => n171, A2 => n133, ZN => ab_24_18_port);
   U694 : NOR2_X1 port map( A1 => n172, A2 => n133, ZN => ab_24_17_port);
   U695 : NOR2_X1 port map( A1 => n173, A2 => n133, ZN => ab_24_16_port);
   U696 : NOR2_X1 port map( A1 => n174, A2 => n133, ZN => ab_24_15_port);
   U697 : NOR2_X1 port map( A1 => n175, A2 => n133, ZN => ab_24_14_port);
   U698 : NOR2_X1 port map( A1 => n176, A2 => n133, ZN => ab_24_13_port);
   U699 : NOR2_X1 port map( A1 => n177, A2 => n133, ZN => ab_24_12_port);
   U700 : NOR2_X1 port map( A1 => n178, A2 => n133, ZN => ab_24_11_port);
   U701 : NOR2_X1 port map( A1 => n179, A2 => n133, ZN => ab_24_10_port);
   U702 : NOR2_X1 port map( A1 => n189, A2 => n133, ZN => ab_24_0_port);
   U703 : NOR2_X1 port map( A1 => n180, A2 => n134, ZN => ab_23_9_port);
   U704 : NOR2_X1 port map( A1 => n181, A2 => n134, ZN => ab_23_8_port);
   U705 : NOR2_X1 port map( A1 => n182, A2 => n134, ZN => ab_23_7_port);
   U706 : NOR2_X1 port map( A1 => n183, A2 => n134, ZN => ab_23_6_port);
   U707 : NOR2_X1 port map( A1 => n184, A2 => n134, ZN => ab_23_5_port);
   U708 : NOR2_X1 port map( A1 => n185, A2 => n134, ZN => ab_23_4_port);
   U709 : NOR2_X1 port map( A1 => n186, A2 => n134, ZN => ab_23_3_port);
   U710 : NOR2_X1 port map( A1 => n158, A2 => n134, ZN => ab_23_31_port);
   U711 : NOR2_X1 port map( A1 => n159, A2 => n134, ZN => ab_23_30_port);
   U712 : NOR2_X1 port map( A1 => n187, A2 => n134, ZN => ab_23_2_port);
   U713 : NOR2_X1 port map( A1 => n160, A2 => n134, ZN => ab_23_29_port);
   U714 : NOR2_X1 port map( A1 => n161, A2 => n134, ZN => ab_23_28_port);
   U715 : NOR2_X1 port map( A1 => n162, A2 => n134, ZN => ab_23_27_port);
   U716 : NOR2_X1 port map( A1 => n163, A2 => n134, ZN => ab_23_26_port);
   U717 : NOR2_X1 port map( A1 => n164, A2 => n134, ZN => ab_23_25_port);
   U718 : NOR2_X1 port map( A1 => n165, A2 => n134, ZN => ab_23_24_port);
   U719 : NOR2_X1 port map( A1 => n166, A2 => n134, ZN => ab_23_23_port);
   U720 : NOR2_X1 port map( A1 => n167, A2 => n134, ZN => ab_23_22_port);
   U721 : NOR2_X1 port map( A1 => n168, A2 => n134, ZN => ab_23_21_port);
   U722 : NOR2_X1 port map( A1 => n169, A2 => n134, ZN => ab_23_20_port);
   U723 : NOR2_X1 port map( A1 => n188, A2 => n134, ZN => ab_23_1_port);
   U724 : NOR2_X1 port map( A1 => n170, A2 => n134, ZN => ab_23_19_port);
   U725 : NOR2_X1 port map( A1 => n171, A2 => n134, ZN => ab_23_18_port);
   U726 : NOR2_X1 port map( A1 => n172, A2 => n134, ZN => ab_23_17_port);
   U727 : NOR2_X1 port map( A1 => n173, A2 => n134, ZN => ab_23_16_port);
   U728 : NOR2_X1 port map( A1 => n174, A2 => n134, ZN => ab_23_15_port);
   U729 : NOR2_X1 port map( A1 => n175, A2 => n134, ZN => ab_23_14_port);
   U730 : NOR2_X1 port map( A1 => n176, A2 => n134, ZN => ab_23_13_port);
   U731 : NOR2_X1 port map( A1 => n177, A2 => n134, ZN => ab_23_12_port);
   U732 : NOR2_X1 port map( A1 => n178, A2 => n134, ZN => ab_23_11_port);
   U733 : NOR2_X1 port map( A1 => n179, A2 => n134, ZN => ab_23_10_port);
   U734 : NOR2_X1 port map( A1 => n189, A2 => n134, ZN => ab_23_0_port);
   U735 : NOR2_X1 port map( A1 => n180, A2 => n135, ZN => ab_22_9_port);
   U736 : NOR2_X1 port map( A1 => n181, A2 => n135, ZN => ab_22_8_port);
   U737 : NOR2_X1 port map( A1 => n182, A2 => n135, ZN => ab_22_7_port);
   U738 : NOR2_X1 port map( A1 => n183, A2 => n135, ZN => ab_22_6_port);
   U739 : NOR2_X1 port map( A1 => n184, A2 => n135, ZN => ab_22_5_port);
   U740 : NOR2_X1 port map( A1 => n185, A2 => n135, ZN => ab_22_4_port);
   U741 : NOR2_X1 port map( A1 => n186, A2 => n135, ZN => ab_22_3_port);
   U742 : NOR2_X1 port map( A1 => n158, A2 => n135, ZN => ab_22_31_port);
   U743 : NOR2_X1 port map( A1 => n159, A2 => n135, ZN => ab_22_30_port);
   U744 : NOR2_X1 port map( A1 => n187, A2 => n135, ZN => ab_22_2_port);
   U745 : NOR2_X1 port map( A1 => n160, A2 => n135, ZN => ab_22_29_port);
   U746 : NOR2_X1 port map( A1 => n161, A2 => n135, ZN => ab_22_28_port);
   U747 : NOR2_X1 port map( A1 => n162, A2 => n135, ZN => ab_22_27_port);
   U748 : NOR2_X1 port map( A1 => n163, A2 => n135, ZN => ab_22_26_port);
   U749 : NOR2_X1 port map( A1 => n164, A2 => n135, ZN => ab_22_25_port);
   U750 : NOR2_X1 port map( A1 => n165, A2 => n135, ZN => ab_22_24_port);
   U751 : NOR2_X1 port map( A1 => n166, A2 => n135, ZN => ab_22_23_port);
   U752 : NOR2_X1 port map( A1 => n167, A2 => n135, ZN => ab_22_22_port);
   U753 : NOR2_X1 port map( A1 => n168, A2 => n135, ZN => ab_22_21_port);
   U754 : NOR2_X1 port map( A1 => n169, A2 => n135, ZN => ab_22_20_port);
   U755 : NOR2_X1 port map( A1 => n188, A2 => n135, ZN => ab_22_1_port);
   U756 : NOR2_X1 port map( A1 => n170, A2 => n135, ZN => ab_22_19_port);
   U757 : NOR2_X1 port map( A1 => n171, A2 => n135, ZN => ab_22_18_port);
   U758 : NOR2_X1 port map( A1 => n172, A2 => n135, ZN => ab_22_17_port);
   U759 : NOR2_X1 port map( A1 => n173, A2 => n135, ZN => ab_22_16_port);
   U760 : NOR2_X1 port map( A1 => n174, A2 => n135, ZN => ab_22_15_port);
   U761 : NOR2_X1 port map( A1 => n175, A2 => n135, ZN => ab_22_14_port);
   U762 : NOR2_X1 port map( A1 => n176, A2 => n135, ZN => ab_22_13_port);
   U763 : NOR2_X1 port map( A1 => n177, A2 => n135, ZN => ab_22_12_port);
   U764 : NOR2_X1 port map( A1 => n178, A2 => n135, ZN => ab_22_11_port);
   U765 : NOR2_X1 port map( A1 => n179, A2 => n135, ZN => ab_22_10_port);
   U766 : NOR2_X1 port map( A1 => n189, A2 => n135, ZN => ab_22_0_port);
   U767 : NOR2_X1 port map( A1 => n180, A2 => n136, ZN => ab_21_9_port);
   U768 : NOR2_X1 port map( A1 => n181, A2 => n136, ZN => ab_21_8_port);
   U769 : NOR2_X1 port map( A1 => n182, A2 => n136, ZN => ab_21_7_port);
   U770 : NOR2_X1 port map( A1 => n183, A2 => n136, ZN => ab_21_6_port);
   U771 : NOR2_X1 port map( A1 => n184, A2 => n136, ZN => ab_21_5_port);
   U772 : NOR2_X1 port map( A1 => n185, A2 => n136, ZN => ab_21_4_port);
   U773 : NOR2_X1 port map( A1 => n186, A2 => n136, ZN => ab_21_3_port);
   U774 : NOR2_X1 port map( A1 => n158, A2 => n136, ZN => ab_21_31_port);
   U775 : NOR2_X1 port map( A1 => n159, A2 => n136, ZN => ab_21_30_port);
   U776 : NOR2_X1 port map( A1 => n187, A2 => n136, ZN => ab_21_2_port);
   U777 : NOR2_X1 port map( A1 => n160, A2 => n136, ZN => ab_21_29_port);
   U778 : NOR2_X1 port map( A1 => n161, A2 => n136, ZN => ab_21_28_port);
   U779 : NOR2_X1 port map( A1 => n162, A2 => n136, ZN => ab_21_27_port);
   U780 : NOR2_X1 port map( A1 => n163, A2 => n136, ZN => ab_21_26_port);
   U781 : NOR2_X1 port map( A1 => n164, A2 => n136, ZN => ab_21_25_port);
   U782 : NOR2_X1 port map( A1 => n165, A2 => n136, ZN => ab_21_24_port);
   U783 : NOR2_X1 port map( A1 => n166, A2 => n136, ZN => ab_21_23_port);
   U784 : NOR2_X1 port map( A1 => n167, A2 => n136, ZN => ab_21_22_port);
   U785 : NOR2_X1 port map( A1 => n168, A2 => n136, ZN => ab_21_21_port);
   U786 : NOR2_X1 port map( A1 => n169, A2 => n136, ZN => ab_21_20_port);
   U787 : NOR2_X1 port map( A1 => n188, A2 => n136, ZN => ab_21_1_port);
   U788 : NOR2_X1 port map( A1 => n170, A2 => n136, ZN => ab_21_19_port);
   U789 : NOR2_X1 port map( A1 => n171, A2 => n136, ZN => ab_21_18_port);
   U790 : NOR2_X1 port map( A1 => n172, A2 => n136, ZN => ab_21_17_port);
   U791 : NOR2_X1 port map( A1 => n173, A2 => n136, ZN => ab_21_16_port);
   U792 : NOR2_X1 port map( A1 => n174, A2 => n136, ZN => ab_21_15_port);
   U793 : NOR2_X1 port map( A1 => n175, A2 => n136, ZN => ab_21_14_port);
   U794 : NOR2_X1 port map( A1 => n176, A2 => n136, ZN => ab_21_13_port);
   U795 : NOR2_X1 port map( A1 => n177, A2 => n136, ZN => ab_21_12_port);
   U796 : NOR2_X1 port map( A1 => n178, A2 => n136, ZN => ab_21_11_port);
   U797 : NOR2_X1 port map( A1 => n179, A2 => n136, ZN => ab_21_10_port);
   U798 : NOR2_X1 port map( A1 => n189, A2 => n136, ZN => ab_21_0_port);
   U799 : NOR2_X1 port map( A1 => n180, A2 => n137, ZN => ab_20_9_port);
   U800 : NOR2_X1 port map( A1 => n181, A2 => n137, ZN => ab_20_8_port);
   U801 : NOR2_X1 port map( A1 => n182, A2 => n137, ZN => ab_20_7_port);
   U802 : NOR2_X1 port map( A1 => n183, A2 => n137, ZN => ab_20_6_port);
   U803 : NOR2_X1 port map( A1 => n184, A2 => n137, ZN => ab_20_5_port);
   U804 : NOR2_X1 port map( A1 => n185, A2 => n137, ZN => ab_20_4_port);
   U805 : NOR2_X1 port map( A1 => n186, A2 => n137, ZN => ab_20_3_port);
   U806 : NOR2_X1 port map( A1 => n158, A2 => n137, ZN => ab_20_31_port);
   U807 : NOR2_X1 port map( A1 => n159, A2 => n137, ZN => ab_20_30_port);
   U808 : NOR2_X1 port map( A1 => n187, A2 => n137, ZN => ab_20_2_port);
   U809 : NOR2_X1 port map( A1 => n160, A2 => n137, ZN => ab_20_29_port);
   U810 : NOR2_X1 port map( A1 => n161, A2 => n137, ZN => ab_20_28_port);
   U811 : NOR2_X1 port map( A1 => n162, A2 => n137, ZN => ab_20_27_port);
   U812 : NOR2_X1 port map( A1 => n163, A2 => n137, ZN => ab_20_26_port);
   U813 : NOR2_X1 port map( A1 => n164, A2 => n137, ZN => ab_20_25_port);
   U814 : NOR2_X1 port map( A1 => n165, A2 => n137, ZN => ab_20_24_port);
   U815 : NOR2_X1 port map( A1 => n166, A2 => n137, ZN => ab_20_23_port);
   U816 : NOR2_X1 port map( A1 => n167, A2 => n137, ZN => ab_20_22_port);
   U817 : NOR2_X1 port map( A1 => n168, A2 => n137, ZN => ab_20_21_port);
   U818 : NOR2_X1 port map( A1 => n169, A2 => n137, ZN => ab_20_20_port);
   U819 : NOR2_X1 port map( A1 => n188, A2 => n137, ZN => ab_20_1_port);
   U820 : NOR2_X1 port map( A1 => n170, A2 => n137, ZN => ab_20_19_port);
   U821 : NOR2_X1 port map( A1 => n171, A2 => n137, ZN => ab_20_18_port);
   U822 : NOR2_X1 port map( A1 => n172, A2 => n137, ZN => ab_20_17_port);
   U823 : NOR2_X1 port map( A1 => n173, A2 => n137, ZN => ab_20_16_port);
   U824 : NOR2_X1 port map( A1 => n174, A2 => n137, ZN => ab_20_15_port);
   U825 : NOR2_X1 port map( A1 => n175, A2 => n137, ZN => ab_20_14_port);
   U826 : NOR2_X1 port map( A1 => n176, A2 => n137, ZN => ab_20_13_port);
   U827 : NOR2_X1 port map( A1 => n177, A2 => n137, ZN => ab_20_12_port);
   U828 : NOR2_X1 port map( A1 => n178, A2 => n137, ZN => ab_20_11_port);
   U829 : NOR2_X1 port map( A1 => n179, A2 => n137, ZN => ab_20_10_port);
   U830 : NOR2_X1 port map( A1 => n189, A2 => n137, ZN => ab_20_0_port);
   U831 : NOR2_X1 port map( A1 => n180, A2 => n156, ZN => ab_1_9_port);
   U832 : NOR2_X1 port map( A1 => n181, A2 => n156, ZN => ab_1_8_port);
   U833 : NOR2_X1 port map( A1 => n182, A2 => n156, ZN => ab_1_7_port);
   U834 : NOR2_X1 port map( A1 => n183, A2 => n156, ZN => ab_1_6_port);
   U835 : NOR2_X1 port map( A1 => n184, A2 => n156, ZN => ab_1_5_port);
   U836 : NOR2_X1 port map( A1 => n185, A2 => n156, ZN => ab_1_4_port);
   U837 : NOR2_X1 port map( A1 => n186, A2 => n156, ZN => ab_1_3_port);
   U838 : NOR2_X1 port map( A1 => n158, A2 => n156, ZN => ab_1_31_port);
   U839 : NOR2_X1 port map( A1 => n159, A2 => n156, ZN => ab_1_30_port);
   U840 : NOR2_X1 port map( A1 => n187, A2 => n156, ZN => ab_1_2_port);
   U841 : NOR2_X1 port map( A1 => n160, A2 => n156, ZN => ab_1_29_port);
   U842 : NOR2_X1 port map( A1 => n161, A2 => n156, ZN => ab_1_28_port);
   U843 : NOR2_X1 port map( A1 => n162, A2 => n156, ZN => ab_1_27_port);
   U844 : NOR2_X1 port map( A1 => n163, A2 => n156, ZN => ab_1_26_port);
   U845 : NOR2_X1 port map( A1 => n164, A2 => n156, ZN => ab_1_25_port);
   U846 : NOR2_X1 port map( A1 => n165, A2 => n156, ZN => ab_1_24_port);
   U847 : NOR2_X1 port map( A1 => n166, A2 => n156, ZN => ab_1_23_port);
   U848 : NOR2_X1 port map( A1 => n167, A2 => n156, ZN => ab_1_22_port);
   U849 : NOR2_X1 port map( A1 => n168, A2 => n156, ZN => ab_1_21_port);
   U850 : NOR2_X1 port map( A1 => n169, A2 => n156, ZN => ab_1_20_port);
   U851 : NOR2_X1 port map( A1 => n188, A2 => n156, ZN => ab_1_1_port);
   U852 : NOR2_X1 port map( A1 => n170, A2 => n156, ZN => ab_1_19_port);
   U853 : NOR2_X1 port map( A1 => n171, A2 => n156, ZN => ab_1_18_port);
   U854 : NOR2_X1 port map( A1 => n172, A2 => n156, ZN => ab_1_17_port);
   U855 : NOR2_X1 port map( A1 => n173, A2 => n156, ZN => ab_1_16_port);
   U856 : NOR2_X1 port map( A1 => n174, A2 => n156, ZN => ab_1_15_port);
   U857 : NOR2_X1 port map( A1 => n175, A2 => n156, ZN => ab_1_14_port);
   U858 : NOR2_X1 port map( A1 => n176, A2 => n156, ZN => ab_1_13_port);
   U859 : NOR2_X1 port map( A1 => n177, A2 => n156, ZN => ab_1_12_port);
   U860 : NOR2_X1 port map( A1 => n178, A2 => n156, ZN => ab_1_11_port);
   U861 : NOR2_X1 port map( A1 => n179, A2 => n156, ZN => ab_1_10_port);
   U862 : NOR2_X1 port map( A1 => n189, A2 => n156, ZN => ab_1_0_port);
   U863 : NOR2_X1 port map( A1 => n180, A2 => n138, ZN => ab_19_9_port);
   U864 : NOR2_X1 port map( A1 => n181, A2 => n138, ZN => ab_19_8_port);
   U865 : NOR2_X1 port map( A1 => n182, A2 => n138, ZN => ab_19_7_port);
   U866 : NOR2_X1 port map( A1 => n183, A2 => n138, ZN => ab_19_6_port);
   U867 : NOR2_X1 port map( A1 => n184, A2 => n138, ZN => ab_19_5_port);
   U868 : NOR2_X1 port map( A1 => n185, A2 => n138, ZN => ab_19_4_port);
   U869 : NOR2_X1 port map( A1 => n186, A2 => n138, ZN => ab_19_3_port);
   U870 : NOR2_X1 port map( A1 => n158, A2 => n138, ZN => ab_19_31_port);
   U871 : NOR2_X1 port map( A1 => n159, A2 => n138, ZN => ab_19_30_port);
   U872 : NOR2_X1 port map( A1 => n187, A2 => n138, ZN => ab_19_2_port);
   U873 : NOR2_X1 port map( A1 => n160, A2 => n138, ZN => ab_19_29_port);
   U874 : NOR2_X1 port map( A1 => n161, A2 => n138, ZN => ab_19_28_port);
   U875 : NOR2_X1 port map( A1 => n162, A2 => n138, ZN => ab_19_27_port);
   U876 : NOR2_X1 port map( A1 => n163, A2 => n138, ZN => ab_19_26_port);
   U877 : NOR2_X1 port map( A1 => n164, A2 => n138, ZN => ab_19_25_port);
   U878 : NOR2_X1 port map( A1 => n165, A2 => n138, ZN => ab_19_24_port);
   U879 : NOR2_X1 port map( A1 => n166, A2 => n138, ZN => ab_19_23_port);
   U880 : NOR2_X1 port map( A1 => n167, A2 => n138, ZN => ab_19_22_port);
   U881 : NOR2_X1 port map( A1 => n168, A2 => n138, ZN => ab_19_21_port);
   U882 : NOR2_X1 port map( A1 => n169, A2 => n138, ZN => ab_19_20_port);
   U883 : NOR2_X1 port map( A1 => n188, A2 => n138, ZN => ab_19_1_port);
   U884 : NOR2_X1 port map( A1 => n170, A2 => n138, ZN => ab_19_19_port);
   U885 : NOR2_X1 port map( A1 => n171, A2 => n138, ZN => ab_19_18_port);
   U886 : NOR2_X1 port map( A1 => n172, A2 => n138, ZN => ab_19_17_port);
   U887 : NOR2_X1 port map( A1 => n173, A2 => n138, ZN => ab_19_16_port);
   U888 : NOR2_X1 port map( A1 => n174, A2 => n138, ZN => ab_19_15_port);
   U889 : NOR2_X1 port map( A1 => n175, A2 => n138, ZN => ab_19_14_port);
   U890 : NOR2_X1 port map( A1 => n176, A2 => n138, ZN => ab_19_13_port);
   U891 : NOR2_X1 port map( A1 => n177, A2 => n138, ZN => ab_19_12_port);
   U892 : NOR2_X1 port map( A1 => n178, A2 => n138, ZN => ab_19_11_port);
   U893 : NOR2_X1 port map( A1 => n179, A2 => n138, ZN => ab_19_10_port);
   U894 : NOR2_X1 port map( A1 => n189, A2 => n138, ZN => ab_19_0_port);
   U895 : NOR2_X1 port map( A1 => n180, A2 => n139, ZN => ab_18_9_port);
   U896 : NOR2_X1 port map( A1 => n181, A2 => n139, ZN => ab_18_8_port);
   U897 : NOR2_X1 port map( A1 => n182, A2 => n139, ZN => ab_18_7_port);
   U898 : NOR2_X1 port map( A1 => n183, A2 => n139, ZN => ab_18_6_port);
   U899 : NOR2_X1 port map( A1 => n184, A2 => n139, ZN => ab_18_5_port);
   U900 : NOR2_X1 port map( A1 => n185, A2 => n139, ZN => ab_18_4_port);
   U901 : NOR2_X1 port map( A1 => n186, A2 => n139, ZN => ab_18_3_port);
   U902 : NOR2_X1 port map( A1 => n158, A2 => n139, ZN => ab_18_31_port);
   U903 : NOR2_X1 port map( A1 => n159, A2 => n139, ZN => ab_18_30_port);
   U904 : NOR2_X1 port map( A1 => n187, A2 => n139, ZN => ab_18_2_port);
   U905 : NOR2_X1 port map( A1 => n160, A2 => n139, ZN => ab_18_29_port);
   U906 : NOR2_X1 port map( A1 => n161, A2 => n139, ZN => ab_18_28_port);
   U907 : NOR2_X1 port map( A1 => n162, A2 => n139, ZN => ab_18_27_port);
   U908 : NOR2_X1 port map( A1 => n163, A2 => n139, ZN => ab_18_26_port);
   U909 : NOR2_X1 port map( A1 => n164, A2 => n139, ZN => ab_18_25_port);
   U910 : NOR2_X1 port map( A1 => n165, A2 => n139, ZN => ab_18_24_port);
   U911 : NOR2_X1 port map( A1 => n166, A2 => n139, ZN => ab_18_23_port);
   U912 : NOR2_X1 port map( A1 => n167, A2 => n139, ZN => ab_18_22_port);
   U913 : NOR2_X1 port map( A1 => n168, A2 => n139, ZN => ab_18_21_port);
   U914 : NOR2_X1 port map( A1 => n169, A2 => n139, ZN => ab_18_20_port);
   U915 : NOR2_X1 port map( A1 => n188, A2 => n139, ZN => ab_18_1_port);
   U916 : NOR2_X1 port map( A1 => n170, A2 => n139, ZN => ab_18_19_port);
   U917 : NOR2_X1 port map( A1 => n171, A2 => n139, ZN => ab_18_18_port);
   U918 : NOR2_X1 port map( A1 => n172, A2 => n139, ZN => ab_18_17_port);
   U919 : NOR2_X1 port map( A1 => n173, A2 => n139, ZN => ab_18_16_port);
   U920 : NOR2_X1 port map( A1 => n174, A2 => n139, ZN => ab_18_15_port);
   U921 : NOR2_X1 port map( A1 => n175, A2 => n139, ZN => ab_18_14_port);
   U922 : NOR2_X1 port map( A1 => n176, A2 => n139, ZN => ab_18_13_port);
   U923 : NOR2_X1 port map( A1 => n177, A2 => n139, ZN => ab_18_12_port);
   U924 : NOR2_X1 port map( A1 => n178, A2 => n139, ZN => ab_18_11_port);
   U925 : NOR2_X1 port map( A1 => n179, A2 => n139, ZN => ab_18_10_port);
   U926 : NOR2_X1 port map( A1 => n189, A2 => n139, ZN => ab_18_0_port);
   U927 : NOR2_X1 port map( A1 => n180, A2 => n140, ZN => ab_17_9_port);
   U928 : NOR2_X1 port map( A1 => n181, A2 => n140, ZN => ab_17_8_port);
   U929 : NOR2_X1 port map( A1 => n182, A2 => n140, ZN => ab_17_7_port);
   U930 : NOR2_X1 port map( A1 => n183, A2 => n140, ZN => ab_17_6_port);
   U931 : NOR2_X1 port map( A1 => n184, A2 => n140, ZN => ab_17_5_port);
   U932 : NOR2_X1 port map( A1 => n185, A2 => n140, ZN => ab_17_4_port);
   U933 : NOR2_X1 port map( A1 => n186, A2 => n140, ZN => ab_17_3_port);
   U934 : NOR2_X1 port map( A1 => n158, A2 => n140, ZN => ab_17_31_port);
   U935 : NOR2_X1 port map( A1 => n159, A2 => n140, ZN => ab_17_30_port);
   U936 : NOR2_X1 port map( A1 => n187, A2 => n140, ZN => ab_17_2_port);
   U937 : NOR2_X1 port map( A1 => n160, A2 => n140, ZN => ab_17_29_port);
   U938 : NOR2_X1 port map( A1 => n161, A2 => n140, ZN => ab_17_28_port);
   U939 : NOR2_X1 port map( A1 => n162, A2 => n140, ZN => ab_17_27_port);
   U940 : NOR2_X1 port map( A1 => n163, A2 => n140, ZN => ab_17_26_port);
   U941 : NOR2_X1 port map( A1 => n164, A2 => n140, ZN => ab_17_25_port);
   U942 : NOR2_X1 port map( A1 => n165, A2 => n140, ZN => ab_17_24_port);
   U943 : NOR2_X1 port map( A1 => n166, A2 => n140, ZN => ab_17_23_port);
   U944 : NOR2_X1 port map( A1 => n167, A2 => n140, ZN => ab_17_22_port);
   U945 : NOR2_X1 port map( A1 => n168, A2 => n140, ZN => ab_17_21_port);
   U946 : NOR2_X1 port map( A1 => n169, A2 => n140, ZN => ab_17_20_port);
   U947 : NOR2_X1 port map( A1 => n188, A2 => n140, ZN => ab_17_1_port);
   U948 : NOR2_X1 port map( A1 => n170, A2 => n140, ZN => ab_17_19_port);
   U949 : NOR2_X1 port map( A1 => n171, A2 => n140, ZN => ab_17_18_port);
   U950 : NOR2_X1 port map( A1 => n172, A2 => n140, ZN => ab_17_17_port);
   U951 : NOR2_X1 port map( A1 => n173, A2 => n140, ZN => ab_17_16_port);
   U952 : NOR2_X1 port map( A1 => n174, A2 => n140, ZN => ab_17_15_port);
   U953 : NOR2_X1 port map( A1 => n175, A2 => n140, ZN => ab_17_14_port);
   U954 : NOR2_X1 port map( A1 => n176, A2 => n140, ZN => ab_17_13_port);
   U955 : NOR2_X1 port map( A1 => n177, A2 => n140, ZN => ab_17_12_port);
   U956 : NOR2_X1 port map( A1 => n178, A2 => n140, ZN => ab_17_11_port);
   U957 : NOR2_X1 port map( A1 => n179, A2 => n140, ZN => ab_17_10_port);
   U958 : NOR2_X1 port map( A1 => n189, A2 => n140, ZN => ab_17_0_port);
   U959 : NOR2_X1 port map( A1 => n180, A2 => n141, ZN => ab_16_9_port);
   U960 : NOR2_X1 port map( A1 => n181, A2 => n141, ZN => ab_16_8_port);
   U961 : NOR2_X1 port map( A1 => n182, A2 => n141, ZN => ab_16_7_port);
   U962 : NOR2_X1 port map( A1 => n183, A2 => n141, ZN => ab_16_6_port);
   U963 : NOR2_X1 port map( A1 => n184, A2 => n141, ZN => ab_16_5_port);
   U964 : NOR2_X1 port map( A1 => n185, A2 => n141, ZN => ab_16_4_port);
   U965 : NOR2_X1 port map( A1 => n186, A2 => n141, ZN => ab_16_3_port);
   U966 : NOR2_X1 port map( A1 => n158, A2 => n141, ZN => ab_16_31_port);
   U967 : NOR2_X1 port map( A1 => n159, A2 => n141, ZN => ab_16_30_port);
   U968 : NOR2_X1 port map( A1 => n187, A2 => n141, ZN => ab_16_2_port);
   U969 : NOR2_X1 port map( A1 => n160, A2 => n141, ZN => ab_16_29_port);
   U970 : NOR2_X1 port map( A1 => n161, A2 => n141, ZN => ab_16_28_port);
   U971 : NOR2_X1 port map( A1 => n162, A2 => n141, ZN => ab_16_27_port);
   U972 : NOR2_X1 port map( A1 => n163, A2 => n141, ZN => ab_16_26_port);
   U973 : NOR2_X1 port map( A1 => n164, A2 => n141, ZN => ab_16_25_port);
   U974 : NOR2_X1 port map( A1 => n165, A2 => n141, ZN => ab_16_24_port);
   U975 : NOR2_X1 port map( A1 => n166, A2 => n141, ZN => ab_16_23_port);
   U976 : NOR2_X1 port map( A1 => n167, A2 => n141, ZN => ab_16_22_port);
   U977 : NOR2_X1 port map( A1 => n168, A2 => n141, ZN => ab_16_21_port);
   U978 : NOR2_X1 port map( A1 => n169, A2 => n141, ZN => ab_16_20_port);
   U979 : NOR2_X1 port map( A1 => n188, A2 => n141, ZN => ab_16_1_port);
   U980 : NOR2_X1 port map( A1 => n170, A2 => n141, ZN => ab_16_19_port);
   U981 : NOR2_X1 port map( A1 => n171, A2 => n141, ZN => ab_16_18_port);
   U982 : NOR2_X1 port map( A1 => n172, A2 => n141, ZN => ab_16_17_port);
   U983 : NOR2_X1 port map( A1 => n173, A2 => n141, ZN => ab_16_16_port);
   U984 : NOR2_X1 port map( A1 => n174, A2 => n141, ZN => ab_16_15_port);
   U985 : NOR2_X1 port map( A1 => n175, A2 => n141, ZN => ab_16_14_port);
   U986 : NOR2_X1 port map( A1 => n176, A2 => n141, ZN => ab_16_13_port);
   U987 : NOR2_X1 port map( A1 => n177, A2 => n141, ZN => ab_16_12_port);
   U988 : NOR2_X1 port map( A1 => n178, A2 => n141, ZN => ab_16_11_port);
   U989 : NOR2_X1 port map( A1 => n179, A2 => n141, ZN => ab_16_10_port);
   U990 : NOR2_X1 port map( A1 => n189, A2 => n141, ZN => ab_16_0_port);
   U991 : NOR2_X1 port map( A1 => n180, A2 => n142, ZN => ab_15_9_port);
   U992 : NOR2_X1 port map( A1 => n181, A2 => n142, ZN => ab_15_8_port);
   U993 : NOR2_X1 port map( A1 => n182, A2 => n142, ZN => ab_15_7_port);
   U994 : NOR2_X1 port map( A1 => n183, A2 => n142, ZN => ab_15_6_port);
   U995 : NOR2_X1 port map( A1 => n184, A2 => n142, ZN => ab_15_5_port);
   U996 : NOR2_X1 port map( A1 => n185, A2 => n142, ZN => ab_15_4_port);
   U997 : NOR2_X1 port map( A1 => n186, A2 => n142, ZN => ab_15_3_port);
   U998 : NOR2_X1 port map( A1 => n158, A2 => n142, ZN => ab_15_31_port);
   U999 : NOR2_X1 port map( A1 => n159, A2 => n142, ZN => ab_15_30_port);
   U1000 : NOR2_X1 port map( A1 => n187, A2 => n142, ZN => ab_15_2_port);
   U1001 : NOR2_X1 port map( A1 => n160, A2 => n142, ZN => ab_15_29_port);
   U1002 : NOR2_X1 port map( A1 => n161, A2 => n142, ZN => ab_15_28_port);
   U1003 : NOR2_X1 port map( A1 => n162, A2 => n142, ZN => ab_15_27_port);
   U1004 : NOR2_X1 port map( A1 => n163, A2 => n142, ZN => ab_15_26_port);
   U1005 : NOR2_X1 port map( A1 => n164, A2 => n142, ZN => ab_15_25_port);
   U1006 : NOR2_X1 port map( A1 => n165, A2 => n142, ZN => ab_15_24_port);
   U1007 : NOR2_X1 port map( A1 => n166, A2 => n142, ZN => ab_15_23_port);
   U1008 : NOR2_X1 port map( A1 => n167, A2 => n142, ZN => ab_15_22_port);
   U1009 : NOR2_X1 port map( A1 => n168, A2 => n142, ZN => ab_15_21_port);
   U1010 : NOR2_X1 port map( A1 => n169, A2 => n142, ZN => ab_15_20_port);
   U1011 : NOR2_X1 port map( A1 => n188, A2 => n142, ZN => ab_15_1_port);
   U1012 : NOR2_X1 port map( A1 => n170, A2 => n142, ZN => ab_15_19_port);
   U1013 : NOR2_X1 port map( A1 => n171, A2 => n142, ZN => ab_15_18_port);
   U1014 : NOR2_X1 port map( A1 => n172, A2 => n142, ZN => ab_15_17_port);
   U1015 : NOR2_X1 port map( A1 => n173, A2 => n142, ZN => ab_15_16_port);
   U1016 : NOR2_X1 port map( A1 => n174, A2 => n142, ZN => ab_15_15_port);
   U1017 : NOR2_X1 port map( A1 => n175, A2 => n142, ZN => ab_15_14_port);
   U1018 : NOR2_X1 port map( A1 => n176, A2 => n142, ZN => ab_15_13_port);
   U1019 : NOR2_X1 port map( A1 => n177, A2 => n142, ZN => ab_15_12_port);
   U1020 : NOR2_X1 port map( A1 => n178, A2 => n142, ZN => ab_15_11_port);
   U1021 : NOR2_X1 port map( A1 => n179, A2 => n142, ZN => ab_15_10_port);
   U1022 : NOR2_X1 port map( A1 => n189, A2 => n142, ZN => ab_15_0_port);
   U1023 : NOR2_X1 port map( A1 => n180, A2 => n143, ZN => ab_14_9_port);
   U1024 : NOR2_X1 port map( A1 => n181, A2 => n143, ZN => ab_14_8_port);
   U1025 : NOR2_X1 port map( A1 => n182, A2 => n143, ZN => ab_14_7_port);
   U1026 : NOR2_X1 port map( A1 => n183, A2 => n143, ZN => ab_14_6_port);
   U1027 : NOR2_X1 port map( A1 => n184, A2 => n143, ZN => ab_14_5_port);
   U1028 : NOR2_X1 port map( A1 => n185, A2 => n143, ZN => ab_14_4_port);
   U1029 : NOR2_X1 port map( A1 => n186, A2 => n143, ZN => ab_14_3_port);
   U1030 : NOR2_X1 port map( A1 => n158, A2 => n143, ZN => ab_14_31_port);
   U1031 : NOR2_X1 port map( A1 => n159, A2 => n143, ZN => ab_14_30_port);
   U1032 : NOR2_X1 port map( A1 => n187, A2 => n143, ZN => ab_14_2_port);
   U1033 : NOR2_X1 port map( A1 => n160, A2 => n143, ZN => ab_14_29_port);
   U1034 : NOR2_X1 port map( A1 => n161, A2 => n143, ZN => ab_14_28_port);
   U1035 : NOR2_X1 port map( A1 => n162, A2 => n143, ZN => ab_14_27_port);
   U1036 : NOR2_X1 port map( A1 => n163, A2 => n143, ZN => ab_14_26_port);
   U1037 : NOR2_X1 port map( A1 => n164, A2 => n143, ZN => ab_14_25_port);
   U1038 : NOR2_X1 port map( A1 => n165, A2 => n143, ZN => ab_14_24_port);
   U1039 : NOR2_X1 port map( A1 => n166, A2 => n143, ZN => ab_14_23_port);
   U1040 : NOR2_X1 port map( A1 => n167, A2 => n143, ZN => ab_14_22_port);
   U1041 : NOR2_X1 port map( A1 => n168, A2 => n143, ZN => ab_14_21_port);
   U1042 : NOR2_X1 port map( A1 => n169, A2 => n143, ZN => ab_14_20_port);
   U1043 : NOR2_X1 port map( A1 => n188, A2 => n143, ZN => ab_14_1_port);
   U1044 : NOR2_X1 port map( A1 => n170, A2 => n143, ZN => ab_14_19_port);
   U1045 : NOR2_X1 port map( A1 => n171, A2 => n143, ZN => ab_14_18_port);
   U1046 : NOR2_X1 port map( A1 => n172, A2 => n143, ZN => ab_14_17_port);
   U1047 : NOR2_X1 port map( A1 => n173, A2 => n143, ZN => ab_14_16_port);
   U1048 : NOR2_X1 port map( A1 => n174, A2 => n143, ZN => ab_14_15_port);
   U1049 : NOR2_X1 port map( A1 => n175, A2 => n143, ZN => ab_14_14_port);
   U1050 : NOR2_X1 port map( A1 => n176, A2 => n143, ZN => ab_14_13_port);
   U1051 : NOR2_X1 port map( A1 => n177, A2 => n143, ZN => ab_14_12_port);
   U1052 : NOR2_X1 port map( A1 => n178, A2 => n143, ZN => ab_14_11_port);
   U1053 : NOR2_X1 port map( A1 => n179, A2 => n143, ZN => ab_14_10_port);
   U1054 : NOR2_X1 port map( A1 => n189, A2 => n143, ZN => ab_14_0_port);
   U1055 : NOR2_X1 port map( A1 => n180, A2 => n144, ZN => ab_13_9_port);
   U1056 : NOR2_X1 port map( A1 => n181, A2 => n144, ZN => ab_13_8_port);
   U1057 : NOR2_X1 port map( A1 => n182, A2 => n144, ZN => ab_13_7_port);
   U1058 : NOR2_X1 port map( A1 => n183, A2 => n144, ZN => ab_13_6_port);
   U1059 : NOR2_X1 port map( A1 => n184, A2 => n144, ZN => ab_13_5_port);
   U1060 : NOR2_X1 port map( A1 => n185, A2 => n144, ZN => ab_13_4_port);
   U1061 : NOR2_X1 port map( A1 => n186, A2 => n144, ZN => ab_13_3_port);
   U1062 : NOR2_X1 port map( A1 => n158, A2 => n144, ZN => ab_13_31_port);
   U1063 : NOR2_X1 port map( A1 => n159, A2 => n144, ZN => ab_13_30_port);
   U1064 : NOR2_X1 port map( A1 => n187, A2 => n144, ZN => ab_13_2_port);
   U1065 : NOR2_X1 port map( A1 => n160, A2 => n144, ZN => ab_13_29_port);
   U1066 : NOR2_X1 port map( A1 => n161, A2 => n144, ZN => ab_13_28_port);
   U1067 : NOR2_X1 port map( A1 => n162, A2 => n144, ZN => ab_13_27_port);
   U1068 : NOR2_X1 port map( A1 => n163, A2 => n144, ZN => ab_13_26_port);
   U1069 : NOR2_X1 port map( A1 => n164, A2 => n144, ZN => ab_13_25_port);
   U1070 : NOR2_X1 port map( A1 => n165, A2 => n144, ZN => ab_13_24_port);
   U1071 : NOR2_X1 port map( A1 => n166, A2 => n144, ZN => ab_13_23_port);
   U1072 : NOR2_X1 port map( A1 => n167, A2 => n144, ZN => ab_13_22_port);
   U1073 : NOR2_X1 port map( A1 => n168, A2 => n144, ZN => ab_13_21_port);
   U1074 : NOR2_X1 port map( A1 => n169, A2 => n144, ZN => ab_13_20_port);
   U1075 : NOR2_X1 port map( A1 => n188, A2 => n144, ZN => ab_13_1_port);
   U1076 : NOR2_X1 port map( A1 => n170, A2 => n144, ZN => ab_13_19_port);
   U1077 : NOR2_X1 port map( A1 => n171, A2 => n144, ZN => ab_13_18_port);
   U1078 : NOR2_X1 port map( A1 => n172, A2 => n144, ZN => ab_13_17_port);
   U1079 : NOR2_X1 port map( A1 => n173, A2 => n144, ZN => ab_13_16_port);
   U1080 : NOR2_X1 port map( A1 => n174, A2 => n144, ZN => ab_13_15_port);
   U1081 : NOR2_X1 port map( A1 => n175, A2 => n144, ZN => ab_13_14_port);
   U1082 : NOR2_X1 port map( A1 => n176, A2 => n144, ZN => ab_13_13_port);
   U1083 : NOR2_X1 port map( A1 => n177, A2 => n144, ZN => ab_13_12_port);
   U1084 : NOR2_X1 port map( A1 => n178, A2 => n144, ZN => ab_13_11_port);
   U1085 : NOR2_X1 port map( A1 => n179, A2 => n144, ZN => ab_13_10_port);
   U1086 : NOR2_X1 port map( A1 => n189, A2 => n144, ZN => ab_13_0_port);
   U1087 : NOR2_X1 port map( A1 => n180, A2 => n145, ZN => ab_12_9_port);
   U1088 : NOR2_X1 port map( A1 => n181, A2 => n145, ZN => ab_12_8_port);
   U1089 : NOR2_X1 port map( A1 => n182, A2 => n145, ZN => ab_12_7_port);
   U1090 : NOR2_X1 port map( A1 => n183, A2 => n145, ZN => ab_12_6_port);
   U1091 : NOR2_X1 port map( A1 => n184, A2 => n145, ZN => ab_12_5_port);
   U1092 : NOR2_X1 port map( A1 => n185, A2 => n145, ZN => ab_12_4_port);
   U1093 : NOR2_X1 port map( A1 => n186, A2 => n145, ZN => ab_12_3_port);
   U1094 : NOR2_X1 port map( A1 => n158, A2 => n145, ZN => ab_12_31_port);
   U1095 : NOR2_X1 port map( A1 => n159, A2 => n145, ZN => ab_12_30_port);
   U1096 : NOR2_X1 port map( A1 => n187, A2 => n145, ZN => ab_12_2_port);
   U1097 : NOR2_X1 port map( A1 => n160, A2 => n145, ZN => ab_12_29_port);
   U1098 : NOR2_X1 port map( A1 => n161, A2 => n145, ZN => ab_12_28_port);
   U1099 : NOR2_X1 port map( A1 => n162, A2 => n145, ZN => ab_12_27_port);
   U1100 : NOR2_X1 port map( A1 => n163, A2 => n145, ZN => ab_12_26_port);
   U1101 : NOR2_X1 port map( A1 => n164, A2 => n145, ZN => ab_12_25_port);
   U1102 : NOR2_X1 port map( A1 => n165, A2 => n145, ZN => ab_12_24_port);
   U1103 : NOR2_X1 port map( A1 => n166, A2 => n145, ZN => ab_12_23_port);
   U1104 : NOR2_X1 port map( A1 => n167, A2 => n145, ZN => ab_12_22_port);
   U1105 : NOR2_X1 port map( A1 => n168, A2 => n145, ZN => ab_12_21_port);
   U1106 : NOR2_X1 port map( A1 => n169, A2 => n145, ZN => ab_12_20_port);
   U1107 : NOR2_X1 port map( A1 => n188, A2 => n145, ZN => ab_12_1_port);
   U1108 : NOR2_X1 port map( A1 => n170, A2 => n145, ZN => ab_12_19_port);
   U1109 : NOR2_X1 port map( A1 => n171, A2 => n145, ZN => ab_12_18_port);
   U1110 : NOR2_X1 port map( A1 => n172, A2 => n145, ZN => ab_12_17_port);
   U1111 : NOR2_X1 port map( A1 => n173, A2 => n145, ZN => ab_12_16_port);
   U1112 : NOR2_X1 port map( A1 => n174, A2 => n145, ZN => ab_12_15_port);
   U1113 : NOR2_X1 port map( A1 => n175, A2 => n145, ZN => ab_12_14_port);
   U1114 : NOR2_X1 port map( A1 => n176, A2 => n145, ZN => ab_12_13_port);
   U1115 : NOR2_X1 port map( A1 => n177, A2 => n145, ZN => ab_12_12_port);
   U1116 : NOR2_X1 port map( A1 => n178, A2 => n145, ZN => ab_12_11_port);
   U1117 : NOR2_X1 port map( A1 => n179, A2 => n145, ZN => ab_12_10_port);
   U1118 : NOR2_X1 port map( A1 => n189, A2 => n145, ZN => ab_12_0_port);
   U1119 : NOR2_X1 port map( A1 => n180, A2 => n146, ZN => ab_11_9_port);
   U1120 : NOR2_X1 port map( A1 => n181, A2 => n146, ZN => ab_11_8_port);
   U1121 : NOR2_X1 port map( A1 => n182, A2 => n146, ZN => ab_11_7_port);
   U1122 : NOR2_X1 port map( A1 => n183, A2 => n146, ZN => ab_11_6_port);
   U1123 : NOR2_X1 port map( A1 => n184, A2 => n146, ZN => ab_11_5_port);
   U1124 : NOR2_X1 port map( A1 => n185, A2 => n146, ZN => ab_11_4_port);
   U1125 : NOR2_X1 port map( A1 => n186, A2 => n146, ZN => ab_11_3_port);
   U1126 : NOR2_X1 port map( A1 => n158, A2 => n146, ZN => ab_11_31_port);
   U1127 : NOR2_X1 port map( A1 => n159, A2 => n146, ZN => ab_11_30_port);
   U1128 : NOR2_X1 port map( A1 => n187, A2 => n146, ZN => ab_11_2_port);
   U1129 : NOR2_X1 port map( A1 => n160, A2 => n146, ZN => ab_11_29_port);
   U1130 : NOR2_X1 port map( A1 => n161, A2 => n146, ZN => ab_11_28_port);
   U1131 : NOR2_X1 port map( A1 => n162, A2 => n146, ZN => ab_11_27_port);
   U1132 : NOR2_X1 port map( A1 => n163, A2 => n146, ZN => ab_11_26_port);
   U1133 : NOR2_X1 port map( A1 => n164, A2 => n146, ZN => ab_11_25_port);
   U1134 : NOR2_X1 port map( A1 => n165, A2 => n146, ZN => ab_11_24_port);
   U1135 : NOR2_X1 port map( A1 => n166, A2 => n146, ZN => ab_11_23_port);
   U1136 : NOR2_X1 port map( A1 => n167, A2 => n146, ZN => ab_11_22_port);
   U1137 : NOR2_X1 port map( A1 => n168, A2 => n146, ZN => ab_11_21_port);
   U1138 : NOR2_X1 port map( A1 => n169, A2 => n146, ZN => ab_11_20_port);
   U1139 : NOR2_X1 port map( A1 => n188, A2 => n146, ZN => ab_11_1_port);
   U1140 : NOR2_X1 port map( A1 => n170, A2 => n146, ZN => ab_11_19_port);
   U1141 : NOR2_X1 port map( A1 => n171, A2 => n146, ZN => ab_11_18_port);
   U1142 : NOR2_X1 port map( A1 => n172, A2 => n146, ZN => ab_11_17_port);
   U1143 : NOR2_X1 port map( A1 => n173, A2 => n146, ZN => ab_11_16_port);
   U1144 : NOR2_X1 port map( A1 => n174, A2 => n146, ZN => ab_11_15_port);
   U1145 : NOR2_X1 port map( A1 => n175, A2 => n146, ZN => ab_11_14_port);
   U1146 : NOR2_X1 port map( A1 => n176, A2 => n146, ZN => ab_11_13_port);
   U1147 : NOR2_X1 port map( A1 => n177, A2 => n146, ZN => ab_11_12_port);
   U1148 : NOR2_X1 port map( A1 => n178, A2 => n146, ZN => ab_11_11_port);
   U1149 : NOR2_X1 port map( A1 => n179, A2 => n146, ZN => ab_11_10_port);
   U1150 : NOR2_X1 port map( A1 => n189, A2 => n146, ZN => ab_11_0_port);
   U1151 : NOR2_X1 port map( A1 => n180, A2 => n147, ZN => ab_10_9_port);
   U1152 : NOR2_X1 port map( A1 => n181, A2 => n147, ZN => ab_10_8_port);
   U1153 : NOR2_X1 port map( A1 => n182, A2 => n147, ZN => ab_10_7_port);
   U1154 : NOR2_X1 port map( A1 => n183, A2 => n147, ZN => ab_10_6_port);
   U1155 : NOR2_X1 port map( A1 => n184, A2 => n147, ZN => ab_10_5_port);
   U1156 : NOR2_X1 port map( A1 => n185, A2 => n147, ZN => ab_10_4_port);
   U1157 : NOR2_X1 port map( A1 => n186, A2 => n147, ZN => ab_10_3_port);
   U1158 : NOR2_X1 port map( A1 => n158, A2 => n147, ZN => ab_10_31_port);
   U1159 : NOR2_X1 port map( A1 => n159, A2 => n147, ZN => ab_10_30_port);
   U1160 : NOR2_X1 port map( A1 => n187, A2 => n147, ZN => ab_10_2_port);
   U1161 : NOR2_X1 port map( A1 => n160, A2 => n147, ZN => ab_10_29_port);
   U1162 : NOR2_X1 port map( A1 => n161, A2 => n147, ZN => ab_10_28_port);
   U1163 : NOR2_X1 port map( A1 => n162, A2 => n147, ZN => ab_10_27_port);
   U1164 : NOR2_X1 port map( A1 => n163, A2 => n147, ZN => ab_10_26_port);
   U1165 : NOR2_X1 port map( A1 => n164, A2 => n147, ZN => ab_10_25_port);
   U1166 : NOR2_X1 port map( A1 => n165, A2 => n147, ZN => ab_10_24_port);
   U1167 : NOR2_X1 port map( A1 => n166, A2 => n147, ZN => ab_10_23_port);
   U1168 : NOR2_X1 port map( A1 => n167, A2 => n147, ZN => ab_10_22_port);
   U1169 : NOR2_X1 port map( A1 => n168, A2 => n147, ZN => ab_10_21_port);
   U1170 : NOR2_X1 port map( A1 => n169, A2 => n147, ZN => ab_10_20_port);
   U1171 : NOR2_X1 port map( A1 => n188, A2 => n147, ZN => ab_10_1_port);
   U1172 : NOR2_X1 port map( A1 => n170, A2 => n147, ZN => ab_10_19_port);
   U1173 : NOR2_X1 port map( A1 => n171, A2 => n147, ZN => ab_10_18_port);
   U1174 : NOR2_X1 port map( A1 => n172, A2 => n147, ZN => ab_10_17_port);
   U1175 : NOR2_X1 port map( A1 => n173, A2 => n147, ZN => ab_10_16_port);
   U1176 : NOR2_X1 port map( A1 => n174, A2 => n147, ZN => ab_10_15_port);
   U1177 : NOR2_X1 port map( A1 => n175, A2 => n147, ZN => ab_10_14_port);
   U1178 : NOR2_X1 port map( A1 => n176, A2 => n147, ZN => ab_10_13_port);
   U1179 : NOR2_X1 port map( A1 => n177, A2 => n147, ZN => ab_10_12_port);
   U1180 : NOR2_X1 port map( A1 => n178, A2 => n147, ZN => ab_10_11_port);
   U1181 : NOR2_X1 port map( A1 => n179, A2 => n147, ZN => ab_10_10_port);
   U1182 : NOR2_X1 port map( A1 => n189, A2 => n147, ZN => ab_10_0_port);
   U1183 : NOR2_X1 port map( A1 => n180, A2 => n157, ZN => ab_0_9_port);
   U1184 : NOR2_X1 port map( A1 => n181, A2 => n157, ZN => ab_0_8_port);
   U1185 : NOR2_X1 port map( A1 => n182, A2 => n157, ZN => ab_0_7_port);
   U1186 : NOR2_X1 port map( A1 => n183, A2 => n157, ZN => ab_0_6_port);
   U1187 : NOR2_X1 port map( A1 => n184, A2 => n157, ZN => ab_0_5_port);
   U1188 : NOR2_X1 port map( A1 => n185, A2 => n157, ZN => ab_0_4_port);
   U1189 : NOR2_X1 port map( A1 => n186, A2 => n157, ZN => ab_0_3_port);
   U1190 : NOR2_X1 port map( A1 => n158, A2 => n157, ZN => ab_0_31_port);
   U1191 : NOR2_X1 port map( A1 => n159, A2 => n157, ZN => ab_0_30_port);
   U1192 : NOR2_X1 port map( A1 => n187, A2 => n157, ZN => ab_0_2_port);
   U1193 : NOR2_X1 port map( A1 => n160, A2 => n157, ZN => ab_0_29_port);
   U1194 : NOR2_X1 port map( A1 => n161, A2 => n157, ZN => ab_0_28_port);
   U1195 : NOR2_X1 port map( A1 => n162, A2 => n157, ZN => ab_0_27_port);
   U1196 : NOR2_X1 port map( A1 => n163, A2 => n157, ZN => ab_0_26_port);
   U1197 : NOR2_X1 port map( A1 => n164, A2 => n157, ZN => ab_0_25_port);
   U1198 : NOR2_X1 port map( A1 => n165, A2 => n157, ZN => ab_0_24_port);
   U1199 : NOR2_X1 port map( A1 => n166, A2 => n157, ZN => ab_0_23_port);
   U1200 : NOR2_X1 port map( A1 => n167, A2 => n157, ZN => ab_0_22_port);
   U1201 : NOR2_X1 port map( A1 => n168, A2 => n157, ZN => ab_0_21_port);
   U1202 : NOR2_X1 port map( A1 => n169, A2 => n157, ZN => ab_0_20_port);
   U1203 : NOR2_X1 port map( A1 => n188, A2 => n157, ZN => ab_0_1_port);
   U1204 : NOR2_X1 port map( A1 => n170, A2 => n157, ZN => ab_0_19_port);
   U1205 : NOR2_X1 port map( A1 => n171, A2 => n157, ZN => ab_0_18_port);
   U1206 : NOR2_X1 port map( A1 => n172, A2 => n157, ZN => ab_0_17_port);
   U1207 : NOR2_X1 port map( A1 => n173, A2 => n157, ZN => ab_0_16_port);
   U1208 : NOR2_X1 port map( A1 => n174, A2 => n157, ZN => ab_0_15_port);
   U1209 : NOR2_X1 port map( A1 => n175, A2 => n157, ZN => ab_0_14_port);
   U1210 : NOR2_X1 port map( A1 => n176, A2 => n157, ZN => ab_0_13_port);
   U1211 : NOR2_X1 port map( A1 => n177, A2 => n157, ZN => ab_0_12_port);
   U1212 : NOR2_X1 port map( A1 => n178, A2 => n157, ZN => ab_0_11_port);
   U1213 : NOR2_X1 port map( A1 => n179, A2 => n157, ZN => ab_0_10_port);
   U1214 : NOR2_X1 port map( A1 => n189, A2 => n157, ZN => PRODUCT(0));
   n191 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_N64.all;

entity ALU_N64_DW01_addsub_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (64 downto 0);  CO : out std_logic);

end ALU_N64_DW01_addsub_0;

architecture SYN_rpl of ALU_N64_DW01_addsub_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_64_port, carry_63_port, carry_62_port, carry_61_port, 
      carry_60_port, carry_59_port, carry_58_port, carry_57_port, carry_56_port
      , carry_55_port, carry_54_port, carry_53_port, carry_52_port, 
      carry_51_port, carry_50_port, carry_49_port, carry_48_port, carry_47_port
      , carry_46_port, carry_45_port, carry_44_port, carry_43_port, 
      carry_42_port, carry_41_port, carry_40_port, carry_39_port, carry_38_port
      , carry_37_port, carry_36_port, carry_35_port, carry_34_port, 
      carry_33_port, carry_32_port, carry_31_port, carry_30_port, carry_29_port
      , carry_28_port, carry_27_port, carry_26_port, carry_25_port, 
      carry_24_port, carry_23_port, carry_22_port, carry_21_port, carry_20_port
      , carry_19_port, carry_18_port, carry_17_port, carry_16_port, 
      carry_15_port, carry_14_port, carry_13_port, carry_12_port, carry_11_port
      , carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      B_AS_63_port, B_AS_62_port, B_AS_61_port, B_AS_60_port, B_AS_59_port, 
      B_AS_58_port, B_AS_57_port, B_AS_56_port, B_AS_55_port, B_AS_54_port, 
      B_AS_53_port, B_AS_52_port, B_AS_51_port, B_AS_50_port, B_AS_49_port, 
      B_AS_48_port, B_AS_47_port, B_AS_46_port, B_AS_45_port, B_AS_44_port, 
      B_AS_43_port, B_AS_42_port, B_AS_41_port, B_AS_40_port, B_AS_39_port, 
      B_AS_38_port, B_AS_37_port, B_AS_36_port, B_AS_35_port, B_AS_34_port, 
      B_AS_33_port, B_AS_32_port, B_AS_31_port, B_AS_30_port, B_AS_29_port, 
      B_AS_28_port, B_AS_27_port, B_AS_26_port, B_AS_25_port, B_AS_24_port, 
      B_AS_23_port, B_AS_22_port, B_AS_21_port, B_AS_20_port, B_AS_19_port, 
      B_AS_18_port, B_AS_17_port, B_AS_16_port, B_AS_15_port, B_AS_14_port, 
      B_AS_13_port, B_AS_12_port, B_AS_11_port, B_AS_10_port, B_AS_9_port, 
      B_AS_8_port, B_AS_7_port, B_AS_6_port, B_AS_5_port, B_AS_4_port, 
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B_AS_63_port, CI => carry_63_port, 
                           CO => carry_64_port, S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B_AS_62_port, CI => carry_62_port, 
                           CO => carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B_AS_61_port, CI => carry_61_port, 
                           CO => carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B_AS_60_port, CI => carry_60_port, 
                           CO => carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B_AS_59_port, CI => carry_59_port, 
                           CO => carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B_AS_58_port, CI => carry_58_port, 
                           CO => carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B_AS_57_port, CI => carry_57_port, 
                           CO => carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B_AS_56_port, CI => carry_56_port, 
                           CO => carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B_AS_55_port, CI => carry_55_port, 
                           CO => carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B_AS_54_port, CI => carry_54_port, 
                           CO => carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B_AS_53_port, CI => carry_53_port, 
                           CO => carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B_AS_52_port, CI => carry_52_port, 
                           CO => carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B_AS_51_port, CI => carry_51_port, 
                           CO => carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B_AS_50_port, CI => carry_50_port, 
                           CO => carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B_AS_49_port, CI => carry_49_port, 
                           CO => carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B_AS_48_port, CI => carry_48_port, 
                           CO => carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B_AS_47_port, CI => carry_47_port, 
                           CO => carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B_AS_46_port, CI => carry_46_port, 
                           CO => carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B_AS_45_port, CI => carry_45_port, 
                           CO => carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B_AS_44_port, CI => carry_44_port, 
                           CO => carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B_AS_43_port, CI => carry_43_port, 
                           CO => carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B_AS_42_port, CI => carry_42_port, 
                           CO => carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B_AS_41_port, CI => carry_41_port, 
                           CO => carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B_AS_40_port, CI => carry_40_port, 
                           CO => carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B_AS_39_port, CI => carry_39_port, 
                           CO => carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B_AS_38_port, CI => carry_38_port, 
                           CO => carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B_AS_37_port, CI => carry_37_port, 
                           CO => carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B_AS_36_port, CI => carry_36_port, 
                           CO => carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B_AS_35_port, CI => carry_35_port, 
                           CO => carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B_AS_34_port, CI => carry_34_port, 
                           CO => carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B_AS_33_port, CI => carry_33_port, 
                           CO => carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B_AS_32_port, CI => carry_32_port, 
                           CO => carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B_AS_31_port, CI => carry_31_port, 
                           CO => carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B_AS_30_port, CI => carry_30_port, 
                           CO => carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B_AS_29_port, CI => carry_29_port, 
                           CO => carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B_AS_28_port, CI => carry_28_port, 
                           CO => carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B_AS_27_port, CI => carry_27_port, 
                           CO => carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B_AS_26_port, CI => carry_26_port, 
                           CO => carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B_AS_25_port, CI => carry_25_port, 
                           CO => carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B_AS_24_port, CI => carry_24_port, 
                           CO => carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B_AS_23_port, CI => carry_23_port, 
                           CO => carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B_AS_22_port, CI => carry_22_port, 
                           CO => carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B_AS_21_port, CI => carry_21_port, 
                           CO => carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B_AS_20_port, CI => carry_20_port, 
                           CO => carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B_AS_19_port, CI => carry_19_port, 
                           CO => carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B_AS_18_port, CI => carry_18_port, 
                           CO => carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B_AS_17_port, CI => carry_17_port, 
                           CO => carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B_AS_16_port, CI => carry_16_port, 
                           CO => carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B_AS_15_port, CI => carry_15_port, 
                           CO => carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B_AS_14_port, CI => carry_14_port, 
                           CO => carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B_AS_13_port, CI => carry_13_port, 
                           CO => carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B_AS_12_port, CI => carry_12_port, 
                           CO => carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B_AS_11_port, CI => carry_11_port, 
                           CO => carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B_AS_10_port, CI => carry_10_port, 
                           CO => carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B_AS_9_port, CI => carry_9_port, CO 
                           => carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B_AS_8_port, CI => carry_8_port, CO 
                           => carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B_AS_7_port, CI => carry_7_port, CO 
                           => carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B_AS_6_port, CI => carry_6_port, CO 
                           => carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B_AS_5_port, CI => carry_5_port, CO 
                           => carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B_AS_4_port, CI => carry_4_port, CO 
                           => carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => ADD_SUB, B => carry_64_port, Z => SUM(64));
   U2 : XOR2_X1 port map( A => B(9), B => ADD_SUB, Z => B_AS_9_port);
   U3 : XOR2_X1 port map( A => B(8), B => ADD_SUB, Z => B_AS_8_port);
   U4 : XOR2_X1 port map( A => B(7), B => ADD_SUB, Z => B_AS_7_port);
   U5 : XOR2_X1 port map( A => B(6), B => ADD_SUB, Z => B_AS_6_port);
   U6 : XOR2_X1 port map( A => B(63), B => ADD_SUB, Z => B_AS_63_port);
   U7 : XOR2_X1 port map( A => B(62), B => ADD_SUB, Z => B_AS_62_port);
   U8 : XOR2_X1 port map( A => B(61), B => ADD_SUB, Z => B_AS_61_port);
   U9 : XOR2_X1 port map( A => B(60), B => ADD_SUB, Z => B_AS_60_port);
   U10 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_AS_5_port);
   U11 : XOR2_X1 port map( A => B(59), B => ADD_SUB, Z => B_AS_59_port);
   U12 : XOR2_X1 port map( A => B(58), B => ADD_SUB, Z => B_AS_58_port);
   U13 : XOR2_X1 port map( A => B(57), B => ADD_SUB, Z => B_AS_57_port);
   U14 : XOR2_X1 port map( A => B(56), B => ADD_SUB, Z => B_AS_56_port);
   U15 : XOR2_X1 port map( A => B(55), B => ADD_SUB, Z => B_AS_55_port);
   U16 : XOR2_X1 port map( A => B(54), B => ADD_SUB, Z => B_AS_54_port);
   U17 : XOR2_X1 port map( A => B(53), B => ADD_SUB, Z => B_AS_53_port);
   U18 : XOR2_X1 port map( A => B(52), B => ADD_SUB, Z => B_AS_52_port);
   U19 : XOR2_X1 port map( A => B(51), B => ADD_SUB, Z => B_AS_51_port);
   U20 : XOR2_X1 port map( A => B(50), B => ADD_SUB, Z => B_AS_50_port);
   U21 : XOR2_X1 port map( A => B(4), B => ADD_SUB, Z => B_AS_4_port);
   U22 : XOR2_X1 port map( A => B(49), B => ADD_SUB, Z => B_AS_49_port);
   U23 : XOR2_X1 port map( A => B(48), B => ADD_SUB, Z => B_AS_48_port);
   U24 : XOR2_X1 port map( A => B(47), B => ADD_SUB, Z => B_AS_47_port);
   U25 : XOR2_X1 port map( A => B(46), B => ADD_SUB, Z => B_AS_46_port);
   U26 : XOR2_X1 port map( A => B(45), B => ADD_SUB, Z => B_AS_45_port);
   U27 : XOR2_X1 port map( A => B(44), B => ADD_SUB, Z => B_AS_44_port);
   U28 : XOR2_X1 port map( A => B(43), B => ADD_SUB, Z => B_AS_43_port);
   U29 : XOR2_X1 port map( A => B(42), B => ADD_SUB, Z => B_AS_42_port);
   U30 : XOR2_X1 port map( A => B(41), B => ADD_SUB, Z => B_AS_41_port);
   U31 : XOR2_X1 port map( A => B(40), B => ADD_SUB, Z => B_AS_40_port);
   U32 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U33 : XOR2_X1 port map( A => B(39), B => ADD_SUB, Z => B_AS_39_port);
   U34 : XOR2_X1 port map( A => B(38), B => ADD_SUB, Z => B_AS_38_port);
   U35 : XOR2_X1 port map( A => B(37), B => ADD_SUB, Z => B_AS_37_port);
   U36 : XOR2_X1 port map( A => B(36), B => ADD_SUB, Z => B_AS_36_port);
   U37 : XOR2_X1 port map( A => B(35), B => ADD_SUB, Z => B_AS_35_port);
   U38 : XOR2_X1 port map( A => B(34), B => ADD_SUB, Z => B_AS_34_port);
   U39 : XOR2_X1 port map( A => B(33), B => ADD_SUB, Z => B_AS_33_port);
   U40 : XOR2_X1 port map( A => B(32), B => ADD_SUB, Z => B_AS_32_port);
   U41 : XOR2_X1 port map( A => B(31), B => ADD_SUB, Z => B_AS_31_port);
   U42 : XOR2_X1 port map( A => B(30), B => ADD_SUB, Z => B_AS_30_port);
   U43 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U44 : XOR2_X1 port map( A => B(29), B => ADD_SUB, Z => B_AS_29_port);
   U45 : XOR2_X1 port map( A => B(28), B => ADD_SUB, Z => B_AS_28_port);
   U46 : XOR2_X1 port map( A => B(27), B => ADD_SUB, Z => B_AS_27_port);
   U47 : XOR2_X1 port map( A => B(26), B => ADD_SUB, Z => B_AS_26_port);
   U48 : XOR2_X1 port map( A => B(25), B => ADD_SUB, Z => B_AS_25_port);
   U49 : XOR2_X1 port map( A => B(24), B => ADD_SUB, Z => B_AS_24_port);
   U50 : XOR2_X1 port map( A => B(23), B => ADD_SUB, Z => B_AS_23_port);
   U51 : XOR2_X1 port map( A => B(22), B => ADD_SUB, Z => B_AS_22_port);
   U52 : XOR2_X1 port map( A => B(21), B => ADD_SUB, Z => B_AS_21_port);
   U53 : XOR2_X1 port map( A => B(20), B => ADD_SUB, Z => B_AS_20_port);
   U54 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U55 : XOR2_X1 port map( A => B(19), B => ADD_SUB, Z => B_AS_19_port);
   U56 : XOR2_X1 port map( A => B(18), B => ADD_SUB, Z => B_AS_18_port);
   U57 : XOR2_X1 port map( A => B(17), B => ADD_SUB, Z => B_AS_17_port);
   U58 : XOR2_X1 port map( A => B(16), B => ADD_SUB, Z => B_AS_16_port);
   U59 : XOR2_X1 port map( A => B(15), B => ADD_SUB, Z => B_AS_15_port);
   U60 : XOR2_X1 port map( A => B(14), B => ADD_SUB, Z => B_AS_14_port);
   U61 : XOR2_X1 port map( A => B(13), B => ADD_SUB, Z => B_AS_13_port);
   U62 : XOR2_X1 port map( A => B(12), B => ADD_SUB, Z => B_AS_12_port);
   U63 : XOR2_X1 port map( A => B(11), B => ADD_SUB, Z => B_AS_11_port);
   U64 : XOR2_X1 port map( A => B(10), B => ADD_SUB, Z => B_AS_10_port);
   U65 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_N64.all;

entity ALU_N64 is

   port( FUNC : in TYPE_OP;  DATA1, DATA2 : in std_logic_vector (63 downto 0); 
         OUTALU : out std_logic_vector (63 downto 0));

end ALU_N64;

architecture SYN_BEHAVIOR_1 of ALU_N64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N64_DW01_cmp2_0
      port( A, B : in std_logic_vector (63 downto 0);  LEQ, TC : in std_logic; 
            LT_LE, GE_GT : out std_logic);
   end component;
   
   component ALU_N64_DW02_mult_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (63 downto 0));
   end component;
   
   component ALU_N64_DW01_addsub_0
      port( A, B : in std_logic_vector (64 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (64 downto 0);  CO : out 
            std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal FUNC_3_port, FUNC_2_port, FUNC_1_port, FUNC_0_port, N46, N47, N48, 
      N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63
      , N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, 
      N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92
      , N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N177, N307, N308, N309, N310, N311, N312, 
      N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, 
      N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, 
      N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, 
      N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, 
      N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N564, N565, 
      N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, 
      N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, 
      N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, 
      N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, 
      N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, 
      N626, N627, n13, n16, n17, n447, n448, n449, n450, n451, n452, n453, n454
      , n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564_port, n565_port, n566_port, n567_port, n568_port, n569_port, 
      n570_port, n571_port, n572_port, n573_port, n574_port, n575_port, 
      n576_port, n577_port, n578_port, n579_port, n580_port, n581_port, 
      n582_port, n583_port, n584_port, n585_port, n586_port, n587_port, 
      n588_port, n589_port, n590_port, n591_port, n592_port, n593_port, 
      n594_port, n595_port, n596_port, n597_port, n598_port, n599_port, 
      n600_port, n601_port, n602_port, n603_port, n604_port, n605_port, 
      n606_port, n607_port, n608_port, n609_port, n610_port, n611_port, 
      n612_port, n613_port, n614_port, n615_port, n616_port, n617_port, 
      n618_port, n619_port, n620_port, n621_port, n622_port, n623_port, 
      n624_port, n625_port, n626_port, n627_port, n628, n629, n630, n631, n632,
      n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n_1043, n_1044 : 
      std_logic;

begin
   (FUNC_3_port, FUNC_2_port, FUNC_1_port, FUNC_0_port) <= 
      TYPE_OP_to_std_logic_vector(FUNC);
   
   n13 <= '0';
   n16 <= '0';
   n17 <= '0';
   OUTALU_reg_63_inst : DLH_X1 port map( G => n452, D => N627, Q => OUTALU(63))
                           ;
   OUTALU_reg_62_inst : DLH_X1 port map( G => n452, D => N626, Q => OUTALU(62))
                           ;
   OUTALU_reg_61_inst : DLH_X1 port map( G => n452, D => N625, Q => OUTALU(61))
                           ;
   OUTALU_reg_60_inst : DLH_X1 port map( G => n452, D => N624, Q => OUTALU(60))
                           ;
   OUTALU_reg_59_inst : DLH_X1 port map( G => n452, D => N623, Q => OUTALU(59))
                           ;
   OUTALU_reg_58_inst : DLH_X1 port map( G => n452, D => N622, Q => OUTALU(58))
                           ;
   OUTALU_reg_57_inst : DLH_X1 port map( G => n452, D => N621, Q => OUTALU(57))
                           ;
   OUTALU_reg_56_inst : DLH_X1 port map( G => n452, D => N620, Q => OUTALU(56))
                           ;
   OUTALU_reg_55_inst : DLH_X1 port map( G => n452, D => N619, Q => OUTALU(55))
                           ;
   OUTALU_reg_54_inst : DLH_X1 port map( G => n452, D => N618, Q => OUTALU(54))
                           ;
   OUTALU_reg_53_inst : DLH_X1 port map( G => n452, D => N617, Q => OUTALU(53))
                           ;
   OUTALU_reg_52_inst : DLH_X1 port map( G => n452, D => N616, Q => OUTALU(52))
                           ;
   OUTALU_reg_51_inst : DLH_X1 port map( G => n452, D => N615, Q => OUTALU(51))
                           ;
   OUTALU_reg_50_inst : DLH_X1 port map( G => n452, D => N614, Q => OUTALU(50))
                           ;
   OUTALU_reg_49_inst : DLH_X1 port map( G => n452, D => N613, Q => OUTALU(49))
                           ;
   OUTALU_reg_48_inst : DLH_X1 port map( G => n452, D => N612, Q => OUTALU(48))
                           ;
   OUTALU_reg_47_inst : DLH_X1 port map( G => n452, D => N611, Q => OUTALU(47))
                           ;
   OUTALU_reg_46_inst : DLH_X1 port map( G => n452, D => N610, Q => OUTALU(46))
                           ;
   OUTALU_reg_45_inst : DLH_X1 port map( G => n452, D => N609, Q => OUTALU(45))
                           ;
   OUTALU_reg_44_inst : DLH_X1 port map( G => n452, D => N608, Q => OUTALU(44))
                           ;
   OUTALU_reg_43_inst : DLH_X1 port map( G => n452, D => N607, Q => OUTALU(43))
                           ;
   OUTALU_reg_42_inst : DLH_X1 port map( G => n452, D => N606, Q => OUTALU(42))
                           ;
   OUTALU_reg_41_inst : DLH_X1 port map( G => n452, D => N605, Q => OUTALU(41))
                           ;
   OUTALU_reg_40_inst : DLH_X1 port map( G => n452, D => N604, Q => OUTALU(40))
                           ;
   OUTALU_reg_39_inst : DLH_X1 port map( G => n452, D => N603, Q => OUTALU(39))
                           ;
   OUTALU_reg_38_inst : DLH_X1 port map( G => n452, D => N602, Q => OUTALU(38))
                           ;
   OUTALU_reg_37_inst : DLH_X1 port map( G => n452, D => N601, Q => OUTALU(37))
                           ;
   OUTALU_reg_36_inst : DLH_X1 port map( G => n452, D => N600, Q => OUTALU(36))
                           ;
   OUTALU_reg_35_inst : DLH_X1 port map( G => n452, D => N599, Q => OUTALU(35))
                           ;
   OUTALU_reg_34_inst : DLH_X1 port map( G => n452, D => N598, Q => OUTALU(34))
                           ;
   OUTALU_reg_33_inst : DLH_X1 port map( G => n452, D => N597, Q => OUTALU(33))
                           ;
   OUTALU_reg_32_inst : DLH_X1 port map( G => n452, D => N596, Q => OUTALU(32))
                           ;
   OUTALU_reg_31_inst : DLH_X1 port map( G => n452, D => N595, Q => OUTALU(31))
                           ;
   OUTALU_reg_30_inst : DLH_X1 port map( G => n452, D => N594, Q => OUTALU(30))
                           ;
   OUTALU_reg_29_inst : DLH_X1 port map( G => n452, D => N593, Q => OUTALU(29))
                           ;
   OUTALU_reg_28_inst : DLH_X1 port map( G => n452, D => N592, Q => OUTALU(28))
                           ;
   OUTALU_reg_27_inst : DLH_X1 port map( G => n452, D => N591, Q => OUTALU(27))
                           ;
   OUTALU_reg_26_inst : DLH_X1 port map( G => n452, D => N590, Q => OUTALU(26))
                           ;
   OUTALU_reg_25_inst : DLH_X1 port map( G => n452, D => N589, Q => OUTALU(25))
                           ;
   OUTALU_reg_24_inst : DLH_X1 port map( G => n452, D => N588, Q => OUTALU(24))
                           ;
   OUTALU_reg_23_inst : DLH_X1 port map( G => n452, D => N587, Q => OUTALU(23))
                           ;
   OUTALU_reg_22_inst : DLH_X1 port map( G => n452, D => N586, Q => OUTALU(22))
                           ;
   OUTALU_reg_21_inst : DLH_X1 port map( G => n452, D => N585, Q => OUTALU(21))
                           ;
   OUTALU_reg_20_inst : DLH_X1 port map( G => n452, D => N584, Q => OUTALU(20))
                           ;
   OUTALU_reg_19_inst : DLH_X1 port map( G => n452, D => N583, Q => OUTALU(19))
                           ;
   OUTALU_reg_18_inst : DLH_X1 port map( G => n452, D => N582, Q => OUTALU(18))
                           ;
   OUTALU_reg_17_inst : DLH_X1 port map( G => n452, D => N581, Q => OUTALU(17))
                           ;
   OUTALU_reg_16_inst : DLH_X1 port map( G => n452, D => N580, Q => OUTALU(16))
                           ;
   OUTALU_reg_15_inst : DLH_X1 port map( G => n452, D => N579, Q => OUTALU(15))
                           ;
   OUTALU_reg_14_inst : DLH_X1 port map( G => n452, D => N578, Q => OUTALU(14))
                           ;
   OUTALU_reg_13_inst : DLH_X1 port map( G => n452, D => N577, Q => OUTALU(13))
                           ;
   OUTALU_reg_12_inst : DLH_X1 port map( G => n452, D => N576, Q => OUTALU(12))
                           ;
   OUTALU_reg_11_inst : DLH_X1 port map( G => n452, D => N575, Q => OUTALU(11))
                           ;
   OUTALU_reg_10_inst : DLH_X1 port map( G => n452, D => N574, Q => OUTALU(10))
                           ;
   OUTALU_reg_9_inst : DLH_X1 port map( G => n452, D => N573, Q => OUTALU(9));
   OUTALU_reg_8_inst : DLH_X1 port map( G => n452, D => N572, Q => OUTALU(8));
   OUTALU_reg_7_inst : DLH_X1 port map( G => n452, D => N571, Q => OUTALU(7));
   OUTALU_reg_6_inst : DLH_X1 port map( G => n452, D => N570, Q => OUTALU(6));
   OUTALU_reg_5_inst : DLH_X1 port map( G => n452, D => N569, Q => OUTALU(5));
   OUTALU_reg_4_inst : DLH_X1 port map( G => n452, D => N568, Q => OUTALU(4));
   OUTALU_reg_3_inst : DLH_X1 port map( G => n452, D => N567, Q => OUTALU(3));
   OUTALU_reg_2_inst : DLH_X1 port map( G => n452, D => N566, Q => OUTALU(2));
   OUTALU_reg_1_inst : DLH_X1 port map( G => n452, D => N565, Q => OUTALU(1));
   OUTALU_reg_0_inst : DLH_X1 port map( G => n452, D => N564, Q => OUTALU(0));
   r74 : ALU_N64_DW01_addsub_0 port map( A(64) => n13, A(63) => DATA1(63), 
                           A(62) => DATA1(62), A(61) => DATA1(61), A(60) => 
                           DATA1(60), A(59) => DATA1(59), A(58) => DATA1(58), 
                           A(57) => DATA1(57), A(56) => DATA1(56), A(55) => 
                           DATA1(55), A(54) => DATA1(54), A(53) => DATA1(53), 
                           A(52) => DATA1(52), A(51) => DATA1(51), A(50) => 
                           DATA1(50), A(49) => DATA1(49), A(48) => DATA1(48), 
                           A(47) => DATA1(47), A(46) => DATA1(46), A(45) => 
                           DATA1(45), A(44) => DATA1(44), A(43) => DATA1(43), 
                           A(42) => DATA1(42), A(41) => DATA1(41), A(40) => 
                           DATA1(40), A(39) => DATA1(39), A(38) => DATA1(38), 
                           A(37) => DATA1(37), A(36) => DATA1(36), A(35) => 
                           DATA1(35), A(34) => DATA1(34), A(33) => DATA1(33), 
                           A(32) => DATA1(32), A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(64) => n13, 
                           B(63) => DATA2(63), B(62) => DATA2(62), B(61) => 
                           DATA2(61), B(60) => DATA2(60), B(59) => DATA2(59), 
                           B(58) => DATA2(58), B(57) => DATA2(57), B(56) => 
                           DATA2(56), B(55) => DATA2(55), B(54) => DATA2(54), 
                           B(53) => DATA2(53), B(52) => DATA2(52), B(51) => 
                           DATA2(51), B(50) => DATA2(50), B(49) => DATA2(49), 
                           B(48) => DATA2(48), B(47) => DATA2(47), B(46) => 
                           DATA2(46), B(45) => DATA2(45), B(44) => DATA2(44), 
                           B(43) => DATA2(43), B(42) => DATA2(42), B(41) => 
                           DATA2(41), B(40) => DATA2(40), B(39) => DATA2(39), 
                           B(38) => DATA2(38), B(37) => DATA2(37), B(36) => 
                           DATA2(36), B(35) => DATA2(35), B(34) => DATA2(34), 
                           B(33) => DATA2(33), B(32) => DATA2(32), B(31) => 
                           DATA2(31), B(30) => DATA2(30), B(29) => DATA2(29), 
                           B(28) => DATA2(28), B(27) => DATA2(27), B(26) => 
                           DATA2(26), B(25) => DATA2(25), B(24) => DATA2(24), 
                           B(23) => DATA2(23), B(22) => DATA2(22), B(21) => 
                           DATA2(21), B(20) => DATA2(20), B(19) => DATA2(19), 
                           B(18) => DATA2(18), B(17) => DATA2(17), B(16) => 
                           DATA2(16), B(15) => DATA2(15), B(14) => DATA2(14), 
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), CI => n13, ADD_SUB => n456, SUM(64) => 
                           N110, SUM(63) => N109, SUM(62) => N108, SUM(61) => 
                           N107, SUM(60) => N106, SUM(59) => N105, SUM(58) => 
                           N104, SUM(57) => N103, SUM(56) => N102, SUM(55) => 
                           N101, SUM(54) => N100, SUM(53) => N99, SUM(52) => 
                           N98, SUM(51) => N97, SUM(50) => N96, SUM(49) => N95,
                           SUM(48) => N94, SUM(47) => N93, SUM(46) => N92, 
                           SUM(45) => N91, SUM(44) => N90, SUM(43) => N89, 
                           SUM(42) => N88, SUM(41) => N87, SUM(40) => N86, 
                           SUM(39) => N85, SUM(38) => N84, SUM(37) => N83, 
                           SUM(36) => N82, SUM(35) => N81, SUM(34) => N80, 
                           SUM(33) => N79, SUM(32) => N78, SUM(31) => N77, 
                           SUM(30) => N76, SUM(29) => N75, SUM(28) => N74, 
                           SUM(27) => N73, SUM(26) => N72, SUM(25) => N71, 
                           SUM(24) => N70, SUM(23) => N69, SUM(22) => N68, 
                           SUM(21) => N67, SUM(20) => N66, SUM(19) => N65, 
                           SUM(18) => N64, SUM(17) => N63, SUM(16) => N62, 
                           SUM(15) => N61, SUM(14) => N60, SUM(13) => N59, 
                           SUM(12) => N58, SUM(11) => N57, SUM(10) => N56, 
                           SUM(9) => N55, SUM(8) => N54, SUM(7) => N53, SUM(6) 
                           => N52, SUM(5) => N51, SUM(4) => N50, SUM(3) => N49,
                           SUM(2) => N48, SUM(1) => N47, SUM(0) => N46, CO => 
                           n_1043);
   mult_42_S2 : ALU_N64_DW02_mult_0 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(31) => 
                           DATA2(31), B(30) => DATA2(30), B(29) => DATA2(29), 
                           B(28) => DATA2(28), B(27) => DATA2(27), B(26) => 
                           DATA2(26), B(25) => DATA2(25), B(24) => DATA2(24), 
                           B(23) => DATA2(23), B(22) => DATA2(22), B(21) => 
                           DATA2(21), B(20) => DATA2(20), B(19) => DATA2(19), 
                           B(18) => DATA2(18), B(17) => DATA2(17), B(16) => 
                           DATA2(16), B(15) => DATA2(15), B(14) => DATA2(14), 
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), TC => n16, PRODUCT(63) => N370, 
                           PRODUCT(62) => N369, PRODUCT(61) => N368, 
                           PRODUCT(60) => N367, PRODUCT(59) => N366, 
                           PRODUCT(58) => N365, PRODUCT(57) => N364, 
                           PRODUCT(56) => N363, PRODUCT(55) => N362, 
                           PRODUCT(54) => N361, PRODUCT(53) => N360, 
                           PRODUCT(52) => N359, PRODUCT(51) => N358, 
                           PRODUCT(50) => N357, PRODUCT(49) => N356, 
                           PRODUCT(48) => N355, PRODUCT(47) => N354, 
                           PRODUCT(46) => N353, PRODUCT(45) => N352, 
                           PRODUCT(44) => N351, PRODUCT(43) => N350, 
                           PRODUCT(42) => N349, PRODUCT(41) => N348, 
                           PRODUCT(40) => N347, PRODUCT(39) => N346, 
                           PRODUCT(38) => N345, PRODUCT(37) => N344, 
                           PRODUCT(36) => N343, PRODUCT(35) => N342, 
                           PRODUCT(34) => N341, PRODUCT(33) => N340, 
                           PRODUCT(32) => N339, PRODUCT(31) => N338, 
                           PRODUCT(30) => N337, PRODUCT(29) => N336, 
                           PRODUCT(28) => N335, PRODUCT(27) => N334, 
                           PRODUCT(26) => N333, PRODUCT(25) => N332, 
                           PRODUCT(24) => N331, PRODUCT(23) => N330, 
                           PRODUCT(22) => N329, PRODUCT(21) => N328, 
                           PRODUCT(20) => N327, PRODUCT(19) => N326, 
                           PRODUCT(18) => N325, PRODUCT(17) => N324, 
                           PRODUCT(16) => N323, PRODUCT(15) => N322, 
                           PRODUCT(14) => N321, PRODUCT(13) => N320, 
                           PRODUCT(12) => N319, PRODUCT(11) => N318, 
                           PRODUCT(10) => N317, PRODUCT(9) => N316, PRODUCT(8) 
                           => N315, PRODUCT(7) => N314, PRODUCT(6) => N313, 
                           PRODUCT(5) => N312, PRODUCT(4) => N311, PRODUCT(3) 
                           => N310, PRODUCT(2) => N309, PRODUCT(1) => N308, 
                           PRODUCT(0) => N307);
   lt_37 : ALU_N64_DW01_cmp2_0 port map( A(63) => DATA1(63), A(62) => DATA1(62)
                           , A(61) => DATA1(61), A(60) => DATA1(60), A(59) => 
                           DATA1(59), A(58) => DATA1(58), A(57) => DATA1(57), 
                           A(56) => DATA1(56), A(55) => DATA1(55), A(54) => 
                           DATA1(54), A(53) => DATA1(53), A(52) => DATA1(52), 
                           A(51) => DATA1(51), A(50) => DATA1(50), A(49) => 
                           DATA1(49), A(48) => DATA1(48), A(47) => DATA1(47), 
                           A(46) => DATA1(46), A(45) => DATA1(45), A(44) => 
                           DATA1(44), A(43) => DATA1(43), A(42) => DATA1(42), 
                           A(41) => DATA1(41), A(40) => DATA1(40), A(39) => 
                           DATA1(39), A(38) => DATA1(38), A(37) => DATA1(37), 
                           A(36) => DATA1(36), A(35) => DATA1(35), A(34) => 
                           DATA1(34), A(33) => DATA1(33), A(32) => DATA1(32), 
                           A(31) => DATA1(31), A(30) => DATA1(30), A(29) => 
                           DATA1(29), A(28) => DATA1(28), A(27) => DATA1(27), 
                           A(26) => DATA1(26), A(25) => DATA1(25), A(24) => 
                           DATA1(24), A(23) => DATA1(23), A(22) => DATA1(22), 
                           A(21) => DATA1(21), A(20) => DATA1(20), A(19) => 
                           DATA1(19), A(18) => DATA1(18), A(17) => DATA1(17), 
                           A(16) => DATA1(16), A(15) => DATA1(15), A(14) => 
                           DATA1(14), A(13) => DATA1(13), A(12) => DATA1(12), 
                           A(11) => DATA1(11), A(10) => DATA1(10), A(9) => 
                           DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7), A(6) 
                           => DATA1(6), A(5) => DATA1(5), A(4) => DATA1(4), 
                           A(3) => DATA1(3), A(2) => DATA1(2), A(1) => DATA1(1)
                           , A(0) => DATA1(0), B(63) => DATA2(63), B(62) => 
                           DATA2(62), B(61) => DATA2(61), B(60) => DATA2(60), 
                           B(59) => DATA2(59), B(58) => DATA2(58), B(57) => 
                           DATA2(57), B(56) => DATA2(56), B(55) => DATA2(55), 
                           B(54) => DATA2(54), B(53) => DATA2(53), B(52) => 
                           DATA2(52), B(51) => DATA2(51), B(50) => DATA2(50), 
                           B(49) => DATA2(49), B(48) => DATA2(48), B(47) => 
                           DATA2(47), B(46) => DATA2(46), B(45) => DATA2(45), 
                           B(44) => DATA2(44), B(43) => DATA2(43), B(42) => 
                           DATA2(42), B(41) => DATA2(41), B(40) => DATA2(40), 
                           B(39) => DATA2(39), B(38) => DATA2(38), B(37) => 
                           DATA2(37), B(36) => DATA2(36), B(35) => DATA2(35), 
                           B(34) => DATA2(34), B(33) => DATA2(33), B(32) => 
                           DATA2(32), B(31) => DATA2(31), B(30) => DATA2(30), 
                           B(29) => DATA2(29), B(28) => DATA2(28), B(27) => 
                           DATA2(27), B(26) => DATA2(26), B(25) => DATA2(25), 
                           B(24) => DATA2(24), B(23) => DATA2(23), B(22) => 
                           DATA2(22), B(21) => DATA2(21), B(20) => DATA2(20), 
                           B(19) => DATA2(19), B(18) => DATA2(18), B(17) => 
                           DATA2(17), B(16) => DATA2(16), B(15) => DATA2(15), 
                           B(14) => DATA2(14), B(13) => DATA2(13), B(12) => 
                           DATA2(12), B(11) => DATA2(11), B(10) => DATA2(10), 
                           B(9) => DATA2(9), B(8) => DATA2(8), B(7) => DATA2(7)
                           , B(6) => DATA2(6), B(5) => DATA2(5), B(4) => 
                           DATA2(4), B(3) => DATA2(3), B(2) => DATA2(2), B(1) 
                           => DATA2(1), B(0) => DATA2(0), LEQ => n17, TC => n17
                           , LT_LE => N177, GE_GT => n_1044);
   U507 : AND4_X1 port map( A1 => n847, A2 => n851, A3 => n867, A4 => n852, ZN 
                           => n447);
   U508 : OR4_X1 port map( A1 => N177, A2 => FUNC_3_port, A3 => n457, A4 => 
                           n458, ZN => n448);
   U509 : OR2_X1 port map( A1 => n852, A2 => FUNC_0_port, ZN => n449);
   U510 : OR2_X1 port map( A1 => n847, A2 => FUNC_0_port, ZN => n450);
   U511 : OR2_X1 port map( A1 => n458, A2 => n847, ZN => n451);
   U512 : INV_X2 port map( A => n447, ZN => n452);
   U513 : AND3_X4 port map( A1 => n858, A2 => n857, A3 => n471, ZN => n483);
   U514 : INV_X4 port map( A => n451, ZN => n453);
   U515 : INV_X4 port map( A => n450, ZN => n454);
   U516 : INV_X4 port map( A => n449, ZN => n455);
   U517 : AOI211_X4 port map( C1 => FUNC_0_port, C2 => N177, A => FUNC_3_port, 
                           B => n457, ZN => n464);
   U518 : INV_X4 port map( A => n448, ZN => n456);
   U519 : INV_X8 port map( A => n852, ZN => n481);
   U520 : INV_X2 port map( A => n851, ZN => n482);
   U521 : INV_X4 port map( A => n462, ZN => n477);
   U522 : NAND4_X1 port map( A1 => n459, A2 => n460, A3 => n461, A4 => n462, ZN
                           => N627);
   U523 : NAND3_X1 port map( A1 => n463, A2 => n458, A3 => DATA1(62), ZN => 
                           n461);
   U524 : NAND2_X1 port map( A1 => N109, A2 => n464, ZN => n460);
   U525 : MUX2_X1 port map( A => n465, B => n466, S => FUNC_2_port, Z => n459);
   U526 : NAND2_X1 port map( A1 => n467, A2 => n468, ZN => n466);
   U527 : MUX2_X1 port map( A => DATA1(63), B => n469, S => DATA2(63), Z => 
                           n467);
   U528 : NAND2_X1 port map( A1 => DATA1(63), A2 => FUNC_0_port, ZN => n469);
   U529 : AOI22_X1 port map( A1 => n470, A2 => FUNC_0_port, B1 => N370, B2 => 
                           n471, ZN => n465);
   U530 : MUX2_X1 port map( A => n472, B => n473, S => FUNC_1_port, Z => n470);
   U531 : AND2_X1 port map( A1 => DATA1(63), A2 => DATA2(63), ZN => n473);
   U532 : AND2_X1 port map( A1 => FUNC_3_port, A2 => DATA1(0), ZN => n472);
   U533 : NAND3_X1 port map( A1 => n474, A2 => n475, A3 => n476, ZN => N626);
   U534 : AOI221_X1 port map( B1 => n453, B2 => DATA1(63), C1 => DATA1(61), C2 
                           => n454, A => n477, ZN => n476);
   U535 : MUX2_X1 port map( A => n478, B => n479, S => DATA1(62), Z => n475);
   U536 : NOR2_X1 port map( A1 => n455, A2 => n480, ZN => n479);
   U537 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(62), Z => n480);
   U538 : NAND2_X1 port map( A1 => DATA2(62), A2 => n481, ZN => n478);
   U539 : AOI22_X1 port map( A1 => N108, A2 => n464, B1 => N369, B2 => n483, ZN
                           => n474);
   U540 : NAND3_X1 port map( A1 => n484, A2 => n485, A3 => n486, ZN => N625);
   U541 : AOI221_X1 port map( B1 => n453, B2 => DATA1(62), C1 => DATA1(60), C2 
                           => n454, A => n477, ZN => n486);
   U542 : MUX2_X1 port map( A => n487, B => n488, S => DATA1(61), Z => n485);
   U543 : NOR2_X1 port map( A1 => n455, A2 => n489, ZN => n488);
   U544 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(61), Z => n489);
   U545 : NAND2_X1 port map( A1 => DATA2(61), A2 => n481, ZN => n487);
   U546 : AOI22_X1 port map( A1 => N107, A2 => n464, B1 => N368, B2 => n483, ZN
                           => n484);
   U547 : NAND3_X1 port map( A1 => n490, A2 => n491, A3 => n492, ZN => N624);
   U548 : AOI221_X1 port map( B1 => n453, B2 => DATA1(61), C1 => DATA1(59), C2 
                           => n454, A => n477, ZN => n492);
   U549 : MUX2_X1 port map( A => n493, B => n494, S => DATA1(60), Z => n491);
   U550 : NOR2_X1 port map( A1 => n455, A2 => n495, ZN => n494);
   U551 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(60), Z => n495);
   U552 : NAND2_X1 port map( A1 => DATA2(60), A2 => n481, ZN => n493);
   U553 : AOI22_X1 port map( A1 => N106, A2 => n464, B1 => N367, B2 => n483, ZN
                           => n490);
   U554 : NAND3_X1 port map( A1 => n496, A2 => n497, A3 => n498, ZN => N623);
   U555 : AOI221_X1 port map( B1 => DATA1(60), B2 => n453, C1 => DATA1(58), C2 
                           => n454, A => n477, ZN => n498);
   U556 : MUX2_X1 port map( A => n499, B => n500, S => DATA1(59), Z => n497);
   U557 : NOR2_X1 port map( A1 => n455, A2 => n501, ZN => n500);
   U558 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(59), Z => n501);
   U559 : NAND2_X1 port map( A1 => DATA2(59), A2 => n481, ZN => n499);
   U560 : AOI22_X1 port map( A1 => N105, A2 => n464, B1 => N366, B2 => n483, ZN
                           => n496);
   U561 : NAND3_X1 port map( A1 => n502, A2 => n503, A3 => n504, ZN => N622);
   U562 : AOI221_X1 port map( B1 => DATA1(59), B2 => n453, C1 => DATA1(57), C2 
                           => n454, A => n477, ZN => n504);
   U563 : MUX2_X1 port map( A => n505, B => n506, S => DATA1(58), Z => n503);
   U564 : NOR2_X1 port map( A1 => n455, A2 => n507, ZN => n506);
   U565 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(58), Z => n507);
   U566 : NAND2_X1 port map( A1 => DATA2(58), A2 => n481, ZN => n505);
   U567 : AOI22_X1 port map( A1 => N104, A2 => n464, B1 => N365, B2 => n483, ZN
                           => n502);
   U568 : NAND3_X1 port map( A1 => n508, A2 => n509, A3 => n510, ZN => N621);
   U569 : AOI221_X1 port map( B1 => DATA1(58), B2 => n453, C1 => DATA1(56), C2 
                           => n454, A => n477, ZN => n510);
   U570 : MUX2_X1 port map( A => n511, B => n512, S => DATA1(57), Z => n509);
   U571 : NOR2_X1 port map( A1 => n455, A2 => n513, ZN => n512);
   U572 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(57), Z => n513);
   U573 : NAND2_X1 port map( A1 => DATA2(57), A2 => n481, ZN => n511);
   U574 : AOI22_X1 port map( A1 => N103, A2 => n464, B1 => N364, B2 => n483, ZN
                           => n508);
   U575 : NAND3_X1 port map( A1 => n514, A2 => n515, A3 => n516, ZN => N620);
   U576 : AOI221_X1 port map( B1 => DATA1(57), B2 => n453, C1 => DATA1(55), C2 
                           => n454, A => n477, ZN => n516);
   U577 : MUX2_X1 port map( A => n517, B => n518, S => DATA1(56), Z => n515);
   U578 : NOR2_X1 port map( A1 => n455, A2 => n519, ZN => n518);
   U579 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(56), Z => n519);
   U580 : NAND2_X1 port map( A1 => DATA2(56), A2 => n481, ZN => n517);
   U581 : AOI22_X1 port map( A1 => N102, A2 => n464, B1 => N363, B2 => n483, ZN
                           => n514);
   U582 : NAND3_X1 port map( A1 => n520, A2 => n521, A3 => n522, ZN => N619);
   U583 : AOI221_X1 port map( B1 => DATA1(56), B2 => n453, C1 => DATA1(54), C2 
                           => n454, A => n477, ZN => n522);
   U584 : MUX2_X1 port map( A => n523, B => n524, S => DATA1(55), Z => n521);
   U585 : NOR2_X1 port map( A1 => n455, A2 => n525, ZN => n524);
   U586 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(55), Z => n525);
   U587 : NAND2_X1 port map( A1 => DATA2(55), A2 => n481, ZN => n523);
   U588 : AOI22_X1 port map( A1 => N101, A2 => n464, B1 => N362, B2 => n483, ZN
                           => n520);
   U589 : NAND3_X1 port map( A1 => n526, A2 => n527, A3 => n528, ZN => N618);
   U590 : AOI221_X1 port map( B1 => DATA1(55), B2 => n453, C1 => DATA1(53), C2 
                           => n454, A => n477, ZN => n528);
   U591 : MUX2_X1 port map( A => n529, B => n530, S => DATA1(54), Z => n527);
   U592 : NOR2_X1 port map( A1 => n455, A2 => n531, ZN => n530);
   U593 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(54), Z => n531);
   U594 : NAND2_X1 port map( A1 => DATA2(54), A2 => n481, ZN => n529);
   U595 : AOI22_X1 port map( A1 => N100, A2 => n464, B1 => N361, B2 => n483, ZN
                           => n526);
   U596 : NAND3_X1 port map( A1 => n532, A2 => n533, A3 => n534, ZN => N617);
   U597 : AOI221_X1 port map( B1 => DATA1(54), B2 => n453, C1 => DATA1(52), C2 
                           => n454, A => n477, ZN => n534);
   U598 : MUX2_X1 port map( A => n535, B => n536, S => DATA1(53), Z => n533);
   U599 : NOR2_X1 port map( A1 => n455, A2 => n537, ZN => n536);
   U600 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(53), Z => n537);
   U601 : NAND2_X1 port map( A1 => DATA2(53), A2 => n481, ZN => n535);
   U602 : AOI22_X1 port map( A1 => N99, A2 => n464, B1 => N360, B2 => n483, ZN 
                           => n532);
   U603 : NAND3_X1 port map( A1 => n538, A2 => n539, A3 => n540, ZN => N616);
   U604 : AOI221_X1 port map( B1 => DATA1(53), B2 => n453, C1 => DATA1(51), C2 
                           => n454, A => n477, ZN => n540);
   U605 : MUX2_X1 port map( A => n541, B => n542, S => DATA1(52), Z => n539);
   U606 : NOR2_X1 port map( A1 => n455, A2 => n543, ZN => n542);
   U607 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(52), Z => n543);
   U608 : NAND2_X1 port map( A1 => DATA2(52), A2 => n481, ZN => n541);
   U609 : AOI22_X1 port map( A1 => N98, A2 => n464, B1 => N359, B2 => n483, ZN 
                           => n538);
   U610 : NAND3_X1 port map( A1 => n544, A2 => n545, A3 => n546, ZN => N615);
   U611 : AOI221_X1 port map( B1 => DATA1(52), B2 => n453, C1 => DATA1(50), C2 
                           => n454, A => n477, ZN => n546);
   U612 : MUX2_X1 port map( A => n547, B => n548, S => DATA1(51), Z => n545);
   U613 : NOR2_X1 port map( A1 => n455, A2 => n549, ZN => n548);
   U614 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(51), Z => n549);
   U615 : NAND2_X1 port map( A1 => DATA2(51), A2 => n481, ZN => n547);
   U616 : AOI22_X1 port map( A1 => N97, A2 => n464, B1 => N358, B2 => n483, ZN 
                           => n544);
   U617 : NAND3_X1 port map( A1 => n550, A2 => n551, A3 => n552, ZN => N614);
   U618 : AOI221_X1 port map( B1 => DATA1(51), B2 => n453, C1 => DATA1(49), C2 
                           => n454, A => n477, ZN => n552);
   U619 : MUX2_X1 port map( A => n553, B => n554, S => DATA1(50), Z => n551);
   U620 : NOR2_X1 port map( A1 => n455, A2 => n555, ZN => n554);
   U621 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(50), Z => n555);
   U622 : NAND2_X1 port map( A1 => DATA2(50), A2 => n481, ZN => n553);
   U623 : AOI22_X1 port map( A1 => N96, A2 => n464, B1 => N357, B2 => n483, ZN 
                           => n550);
   U624 : NAND3_X1 port map( A1 => n556, A2 => n557, A3 => n558, ZN => N613);
   U625 : AOI221_X1 port map( B1 => DATA1(50), B2 => n453, C1 => DATA1(48), C2 
                           => n454, A => n477, ZN => n558);
   U626 : MUX2_X1 port map( A => n559, B => n560, S => DATA1(49), Z => n557);
   U627 : NOR2_X1 port map( A1 => n455, A2 => n561, ZN => n560);
   U628 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(49), Z => n561);
   U629 : NAND2_X1 port map( A1 => DATA2(49), A2 => n481, ZN => n559);
   U630 : AOI22_X1 port map( A1 => N95, A2 => n464, B1 => N356, B2 => n483, ZN 
                           => n556);
   U631 : NAND3_X1 port map( A1 => n562, A2 => n563, A3 => n564_port, ZN => 
                           N612);
   U632 : AOI221_X1 port map( B1 => DATA1(49), B2 => n453, C1 => DATA1(47), C2 
                           => n454, A => n477, ZN => n564_port);
   U633 : MUX2_X1 port map( A => n565_port, B => n566_port, S => DATA1(48), Z 
                           => n563);
   U634 : NOR2_X1 port map( A1 => n455, A2 => n567_port, ZN => n566_port);
   U635 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(48), Z => 
                           n567_port);
   U636 : NAND2_X1 port map( A1 => DATA2(48), A2 => n481, ZN => n565_port);
   U637 : AOI22_X1 port map( A1 => N94, A2 => n464, B1 => N355, B2 => n483, ZN 
                           => n562);
   U638 : NAND3_X1 port map( A1 => n568_port, A2 => n569_port, A3 => n570_port,
                           ZN => N611);
   U639 : AOI221_X1 port map( B1 => DATA1(48), B2 => n453, C1 => DATA1(46), C2 
                           => n454, A => n477, ZN => n570_port);
   U640 : MUX2_X1 port map( A => n571_port, B => n572_port, S => DATA1(47), Z 
                           => n569_port);
   U641 : NOR2_X1 port map( A1 => n455, A2 => n573_port, ZN => n572_port);
   U642 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(47), Z => 
                           n573_port);
   U643 : NAND2_X1 port map( A1 => DATA2(47), A2 => n481, ZN => n571_port);
   U644 : AOI22_X1 port map( A1 => N93, A2 => n464, B1 => N354, B2 => n483, ZN 
                           => n568_port);
   U645 : NAND3_X1 port map( A1 => n574_port, A2 => n575_port, A3 => n576_port,
                           ZN => N610);
   U646 : AOI221_X1 port map( B1 => DATA1(47), B2 => n453, C1 => DATA1(45), C2 
                           => n454, A => n477, ZN => n576_port);
   U647 : MUX2_X1 port map( A => n577_port, B => n578_port, S => DATA1(46), Z 
                           => n575_port);
   U648 : NOR2_X1 port map( A1 => n455, A2 => n579_port, ZN => n578_port);
   U649 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(46), Z => 
                           n579_port);
   U650 : NAND2_X1 port map( A1 => DATA2(46), A2 => n481, ZN => n577_port);
   U651 : AOI22_X1 port map( A1 => N92, A2 => n464, B1 => N353, B2 => n483, ZN 
                           => n574_port);
   U652 : NAND3_X1 port map( A1 => n580_port, A2 => n581_port, A3 => n582_port,
                           ZN => N609);
   U653 : AOI221_X1 port map( B1 => DATA1(46), B2 => n453, C1 => DATA1(44), C2 
                           => n454, A => n477, ZN => n582_port);
   U654 : MUX2_X1 port map( A => n583_port, B => n584_port, S => DATA1(45), Z 
                           => n581_port);
   U655 : NOR2_X1 port map( A1 => n455, A2 => n585_port, ZN => n584_port);
   U656 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(45), Z => 
                           n585_port);
   U657 : NAND2_X1 port map( A1 => DATA2(45), A2 => n481, ZN => n583_port);
   U658 : AOI22_X1 port map( A1 => N91, A2 => n464, B1 => N352, B2 => n483, ZN 
                           => n580_port);
   U659 : NAND3_X1 port map( A1 => n586_port, A2 => n587_port, A3 => n588_port,
                           ZN => N608);
   U660 : AOI221_X1 port map( B1 => DATA1(45), B2 => n453, C1 => DATA1(43), C2 
                           => n454, A => n477, ZN => n588_port);
   U661 : MUX2_X1 port map( A => n589_port, B => n590_port, S => DATA1(44), Z 
                           => n587_port);
   U662 : NOR2_X1 port map( A1 => n455, A2 => n591_port, ZN => n590_port);
   U663 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(44), Z => 
                           n591_port);
   U664 : NAND2_X1 port map( A1 => DATA2(44), A2 => n481, ZN => n589_port);
   U665 : AOI22_X1 port map( A1 => N90, A2 => n464, B1 => N351, B2 => n483, ZN 
                           => n586_port);
   U666 : NAND3_X1 port map( A1 => n592_port, A2 => n593_port, A3 => n594_port,
                           ZN => N607);
   U667 : AOI221_X1 port map( B1 => DATA1(44), B2 => n453, C1 => DATA1(42), C2 
                           => n454, A => n477, ZN => n594_port);
   U668 : MUX2_X1 port map( A => n595_port, B => n596_port, S => DATA1(43), Z 
                           => n593_port);
   U669 : NOR2_X1 port map( A1 => n455, A2 => n597_port, ZN => n596_port);
   U670 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(43), Z => 
                           n597_port);
   U671 : NAND2_X1 port map( A1 => DATA2(43), A2 => n481, ZN => n595_port);
   U672 : AOI22_X1 port map( A1 => N89, A2 => n464, B1 => N350, B2 => n483, ZN 
                           => n592_port);
   U673 : NAND3_X1 port map( A1 => n598_port, A2 => n599_port, A3 => n600_port,
                           ZN => N606);
   U674 : AOI221_X1 port map( B1 => DATA1(43), B2 => n453, C1 => DATA1(41), C2 
                           => n454, A => n477, ZN => n600_port);
   U675 : MUX2_X1 port map( A => n601_port, B => n602_port, S => DATA1(42), Z 
                           => n599_port);
   U676 : NOR2_X1 port map( A1 => n455, A2 => n603_port, ZN => n602_port);
   U677 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(42), Z => 
                           n603_port);
   U678 : NAND2_X1 port map( A1 => DATA2(42), A2 => n481, ZN => n601_port);
   U679 : AOI22_X1 port map( A1 => N88, A2 => n464, B1 => N349, B2 => n483, ZN 
                           => n598_port);
   U680 : NAND3_X1 port map( A1 => n604_port, A2 => n605_port, A3 => n606_port,
                           ZN => N605);
   U681 : AOI221_X1 port map( B1 => DATA1(42), B2 => n453, C1 => DATA1(40), C2 
                           => n454, A => n477, ZN => n606_port);
   U682 : MUX2_X1 port map( A => n607_port, B => n608_port, S => DATA1(41), Z 
                           => n605_port);
   U683 : NOR2_X1 port map( A1 => n455, A2 => n609_port, ZN => n608_port);
   U684 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(41), Z => 
                           n609_port);
   U685 : NAND2_X1 port map( A1 => DATA2(41), A2 => n481, ZN => n607_port);
   U686 : AOI22_X1 port map( A1 => N87, A2 => n464, B1 => N348, B2 => n483, ZN 
                           => n604_port);
   U687 : NAND3_X1 port map( A1 => n610_port, A2 => n611_port, A3 => n612_port,
                           ZN => N604);
   U688 : AOI221_X1 port map( B1 => DATA1(41), B2 => n453, C1 => DATA1(39), C2 
                           => n454, A => n477, ZN => n612_port);
   U689 : MUX2_X1 port map( A => n613_port, B => n614_port, S => DATA1(40), Z 
                           => n611_port);
   U690 : NOR2_X1 port map( A1 => n455, A2 => n615_port, ZN => n614_port);
   U691 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(40), Z => 
                           n615_port);
   U692 : NAND2_X1 port map( A1 => DATA2(40), A2 => n481, ZN => n613_port);
   U693 : AOI22_X1 port map( A1 => N86, A2 => n464, B1 => N347, B2 => n483, ZN 
                           => n610_port);
   U694 : NAND3_X1 port map( A1 => n616_port, A2 => n617_port, A3 => n618_port,
                           ZN => N603);
   U695 : AOI221_X1 port map( B1 => DATA1(40), B2 => n453, C1 => DATA1(38), C2 
                           => n454, A => n477, ZN => n618_port);
   U696 : MUX2_X1 port map( A => n619_port, B => n620_port, S => DATA1(39), Z 
                           => n617_port);
   U697 : NOR2_X1 port map( A1 => n455, A2 => n621_port, ZN => n620_port);
   U698 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(39), Z => 
                           n621_port);
   U699 : NAND2_X1 port map( A1 => DATA2(39), A2 => n481, ZN => n619_port);
   U700 : AOI22_X1 port map( A1 => N85, A2 => n464, B1 => N346, B2 => n483, ZN 
                           => n616_port);
   U701 : NAND3_X1 port map( A1 => n622_port, A2 => n623_port, A3 => n624_port,
                           ZN => N602);
   U702 : AOI221_X1 port map( B1 => DATA1(39), B2 => n453, C1 => DATA1(37), C2 
                           => n454, A => n477, ZN => n624_port);
   U703 : MUX2_X1 port map( A => n625_port, B => n626_port, S => DATA1(38), Z 
                           => n623_port);
   U704 : NOR2_X1 port map( A1 => n455, A2 => n627_port, ZN => n626_port);
   U705 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(38), Z => 
                           n627_port);
   U706 : NAND2_X1 port map( A1 => DATA2(38), A2 => n481, ZN => n625_port);
   U707 : AOI22_X1 port map( A1 => N84, A2 => n464, B1 => N345, B2 => n483, ZN 
                           => n622_port);
   U708 : NAND3_X1 port map( A1 => n628, A2 => n629, A3 => n630, ZN => N601);
   U709 : AOI221_X1 port map( B1 => DATA1(38), B2 => n453, C1 => DATA1(36), C2 
                           => n454, A => n477, ZN => n630);
   U710 : MUX2_X1 port map( A => n631, B => n632, S => DATA1(37), Z => n629);
   U711 : NOR2_X1 port map( A1 => n455, A2 => n633, ZN => n632);
   U712 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(37), Z => n633);
   U713 : NAND2_X1 port map( A1 => DATA2(37), A2 => n481, ZN => n631);
   U714 : AOI22_X1 port map( A1 => N83, A2 => n464, B1 => N344, B2 => n483, ZN 
                           => n628);
   U715 : NAND3_X1 port map( A1 => n634, A2 => n635, A3 => n636, ZN => N600);
   U716 : AOI221_X1 port map( B1 => DATA1(37), B2 => n453, C1 => DATA1(35), C2 
                           => n454, A => n477, ZN => n636);
   U717 : MUX2_X1 port map( A => n637, B => n638, S => DATA1(36), Z => n635);
   U718 : NOR2_X1 port map( A1 => n455, A2 => n639, ZN => n638);
   U719 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(36), Z => n639);
   U720 : NAND2_X1 port map( A1 => DATA2(36), A2 => n481, ZN => n637);
   U721 : AOI22_X1 port map( A1 => N82, A2 => n464, B1 => N343, B2 => n483, ZN 
                           => n634);
   U722 : NAND3_X1 port map( A1 => n640, A2 => n641, A3 => n642, ZN => N599);
   U723 : AOI221_X1 port map( B1 => DATA1(36), B2 => n453, C1 => DATA1(34), C2 
                           => n454, A => n477, ZN => n642);
   U724 : MUX2_X1 port map( A => n643, B => n644, S => DATA1(35), Z => n641);
   U725 : NOR2_X1 port map( A1 => n455, A2 => n645, ZN => n644);
   U726 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(35), Z => n645);
   U727 : NAND2_X1 port map( A1 => DATA2(35), A2 => n481, ZN => n643);
   U728 : AOI22_X1 port map( A1 => N81, A2 => n464, B1 => N342, B2 => n483, ZN 
                           => n640);
   U729 : NAND3_X1 port map( A1 => n646, A2 => n647, A3 => n648, ZN => N598);
   U730 : AOI221_X1 port map( B1 => DATA1(35), B2 => n453, C1 => DATA1(33), C2 
                           => n454, A => n477, ZN => n648);
   U731 : MUX2_X1 port map( A => n649, B => n650, S => DATA1(34), Z => n647);
   U732 : NOR2_X1 port map( A1 => n455, A2 => n651, ZN => n650);
   U733 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(34), Z => n651);
   U734 : NAND2_X1 port map( A1 => DATA2(34), A2 => n481, ZN => n649);
   U735 : AOI22_X1 port map( A1 => N80, A2 => n464, B1 => N341, B2 => n483, ZN 
                           => n646);
   U736 : NAND3_X1 port map( A1 => n652, A2 => n653, A3 => n654, ZN => N597);
   U737 : AOI221_X1 port map( B1 => DATA1(34), B2 => n453, C1 => DATA1(32), C2 
                           => n454, A => n477, ZN => n654);
   U738 : MUX2_X1 port map( A => n655, B => n656, S => DATA1(33), Z => n653);
   U739 : NOR2_X1 port map( A1 => n455, A2 => n657, ZN => n656);
   U740 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(33), Z => n657);
   U741 : NAND2_X1 port map( A1 => DATA2(33), A2 => n481, ZN => n655);
   U742 : AOI22_X1 port map( A1 => N79, A2 => n464, B1 => N340, B2 => n483, ZN 
                           => n652);
   U743 : NAND3_X1 port map( A1 => n658, A2 => n659, A3 => n660, ZN => N596);
   U744 : AOI221_X1 port map( B1 => DATA1(33), B2 => n453, C1 => DATA1(31), C2 
                           => n454, A => n477, ZN => n660);
   U745 : MUX2_X1 port map( A => n661, B => n662, S => DATA1(32), Z => n659);
   U746 : NOR2_X1 port map( A1 => n455, A2 => n663, ZN => n662);
   U747 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(32), Z => n663);
   U748 : NAND2_X1 port map( A1 => DATA2(32), A2 => n481, ZN => n661);
   U749 : AOI22_X1 port map( A1 => N78, A2 => n464, B1 => N339, B2 => n483, ZN 
                           => n658);
   U750 : NAND3_X1 port map( A1 => n664, A2 => n665, A3 => n666, ZN => N595);
   U751 : AOI221_X1 port map( B1 => DATA1(32), B2 => n453, C1 => DATA1(30), C2 
                           => n454, A => n477, ZN => n666);
   U752 : MUX2_X1 port map( A => n667, B => n668, S => DATA1(31), Z => n665);
   U753 : NOR2_X1 port map( A1 => n455, A2 => n669, ZN => n668);
   U754 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(31), Z => n669);
   U755 : NAND2_X1 port map( A1 => DATA2(31), A2 => n481, ZN => n667);
   U756 : AOI22_X1 port map( A1 => N77, A2 => n464, B1 => N338, B2 => n483, ZN 
                           => n664);
   U757 : NAND3_X1 port map( A1 => n670, A2 => n671, A3 => n672, ZN => N594);
   U758 : AOI221_X1 port map( B1 => DATA1(31), B2 => n453, C1 => DATA1(29), C2 
                           => n454, A => n477, ZN => n672);
   U759 : MUX2_X1 port map( A => n673, B => n674, S => DATA1(30), Z => n671);
   U760 : NOR2_X1 port map( A1 => n455, A2 => n675, ZN => n674);
   U761 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(30), Z => n675);
   U762 : NAND2_X1 port map( A1 => DATA2(30), A2 => n481, ZN => n673);
   U763 : AOI22_X1 port map( A1 => N76, A2 => n464, B1 => N337, B2 => n483, ZN 
                           => n670);
   U764 : NAND3_X1 port map( A1 => n676, A2 => n677, A3 => n678, ZN => N593);
   U765 : AOI221_X1 port map( B1 => DATA1(30), B2 => n453, C1 => DATA1(28), C2 
                           => n454, A => n477, ZN => n678);
   U766 : MUX2_X1 port map( A => n679, B => n680, S => DATA1(29), Z => n677);
   U767 : NOR2_X1 port map( A1 => n455, A2 => n681, ZN => n680);
   U768 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(29), Z => n681);
   U769 : NAND2_X1 port map( A1 => DATA2(29), A2 => n481, ZN => n679);
   U770 : AOI22_X1 port map( A1 => N75, A2 => n464, B1 => N336, B2 => n483, ZN 
                           => n676);
   U771 : NAND3_X1 port map( A1 => n682, A2 => n683, A3 => n684, ZN => N592);
   U772 : AOI221_X1 port map( B1 => DATA1(29), B2 => n453, C1 => DATA1(27), C2 
                           => n454, A => n477, ZN => n684);
   U773 : MUX2_X1 port map( A => n685, B => n686, S => DATA1(28), Z => n683);
   U774 : NOR2_X1 port map( A1 => n455, A2 => n687, ZN => n686);
   U775 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(28), Z => n687);
   U776 : NAND2_X1 port map( A1 => DATA2(28), A2 => n481, ZN => n685);
   U777 : AOI22_X1 port map( A1 => N74, A2 => n464, B1 => N335, B2 => n483, ZN 
                           => n682);
   U778 : NAND3_X1 port map( A1 => n688, A2 => n689, A3 => n690, ZN => N591);
   U779 : AOI221_X1 port map( B1 => DATA1(28), B2 => n453, C1 => DATA1(26), C2 
                           => n454, A => n477, ZN => n690);
   U780 : MUX2_X1 port map( A => n691, B => n692, S => DATA1(27), Z => n689);
   U781 : NOR2_X1 port map( A1 => n455, A2 => n693, ZN => n692);
   U782 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(27), Z => n693);
   U783 : NAND2_X1 port map( A1 => DATA2(27), A2 => n481, ZN => n691);
   U784 : AOI22_X1 port map( A1 => N73, A2 => n464, B1 => N334, B2 => n483, ZN 
                           => n688);
   U785 : NAND3_X1 port map( A1 => n694, A2 => n695, A3 => n696, ZN => N590);
   U786 : AOI221_X1 port map( B1 => DATA1(27), B2 => n453, C1 => DATA1(25), C2 
                           => n454, A => n477, ZN => n696);
   U787 : MUX2_X1 port map( A => n697, B => n698, S => DATA1(26), Z => n695);
   U788 : NOR2_X1 port map( A1 => n455, A2 => n699, ZN => n698);
   U789 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(26), Z => n699);
   U790 : NAND2_X1 port map( A1 => DATA2(26), A2 => n481, ZN => n697);
   U791 : AOI22_X1 port map( A1 => N72, A2 => n464, B1 => N333, B2 => n483, ZN 
                           => n694);
   U792 : NAND3_X1 port map( A1 => n700, A2 => n701, A3 => n702, ZN => N589);
   U793 : AOI221_X1 port map( B1 => DATA1(26), B2 => n453, C1 => DATA1(24), C2 
                           => n454, A => n477, ZN => n702);
   U794 : MUX2_X1 port map( A => n703, B => n704, S => DATA1(25), Z => n701);
   U795 : NOR2_X1 port map( A1 => n455, A2 => n705, ZN => n704);
   U796 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(25), Z => n705);
   U797 : NAND2_X1 port map( A1 => DATA2(25), A2 => n481, ZN => n703);
   U798 : AOI22_X1 port map( A1 => N71, A2 => n464, B1 => N332, B2 => n483, ZN 
                           => n700);
   U799 : NAND3_X1 port map( A1 => n706, A2 => n707, A3 => n708, ZN => N588);
   U800 : AOI221_X1 port map( B1 => DATA1(25), B2 => n453, C1 => DATA1(23), C2 
                           => n454, A => n477, ZN => n708);
   U801 : MUX2_X1 port map( A => n709, B => n710, S => DATA1(24), Z => n707);
   U802 : NOR2_X1 port map( A1 => n455, A2 => n711, ZN => n710);
   U803 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(24), Z => n711);
   U804 : NAND2_X1 port map( A1 => DATA2(24), A2 => n481, ZN => n709);
   U805 : AOI22_X1 port map( A1 => N70, A2 => n464, B1 => N331, B2 => n483, ZN 
                           => n706);
   U806 : NAND3_X1 port map( A1 => n712, A2 => n713, A3 => n714, ZN => N587);
   U807 : AOI221_X1 port map( B1 => DATA1(24), B2 => n453, C1 => DATA1(22), C2 
                           => n454, A => n477, ZN => n714);
   U808 : MUX2_X1 port map( A => n715, B => n716, S => DATA1(23), Z => n713);
   U809 : NOR2_X1 port map( A1 => n455, A2 => n717, ZN => n716);
   U810 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(23), Z => n717);
   U811 : NAND2_X1 port map( A1 => DATA2(23), A2 => n481, ZN => n715);
   U812 : AOI22_X1 port map( A1 => N69, A2 => n464, B1 => N330, B2 => n483, ZN 
                           => n712);
   U813 : NAND3_X1 port map( A1 => n718, A2 => n719, A3 => n720, ZN => N586);
   U814 : AOI221_X1 port map( B1 => DATA1(23), B2 => n453, C1 => DATA1(21), C2 
                           => n454, A => n477, ZN => n720);
   U815 : MUX2_X1 port map( A => n721, B => n722, S => DATA1(22), Z => n719);
   U816 : NOR2_X1 port map( A1 => n455, A2 => n723, ZN => n722);
   U817 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(22), Z => n723);
   U818 : NAND2_X1 port map( A1 => DATA2(22), A2 => n481, ZN => n721);
   U819 : AOI22_X1 port map( A1 => N68, A2 => n464, B1 => N329, B2 => n483, ZN 
                           => n718);
   U820 : NAND3_X1 port map( A1 => n724, A2 => n725, A3 => n726, ZN => N585);
   U821 : AOI221_X1 port map( B1 => DATA1(22), B2 => n453, C1 => DATA1(20), C2 
                           => n454, A => n477, ZN => n726);
   U822 : MUX2_X1 port map( A => n727, B => n728, S => DATA1(21), Z => n725);
   U823 : NOR2_X1 port map( A1 => n455, A2 => n729, ZN => n728);
   U824 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(21), Z => n729);
   U825 : NAND2_X1 port map( A1 => DATA2(21), A2 => n481, ZN => n727);
   U826 : AOI22_X1 port map( A1 => N67, A2 => n464, B1 => N328, B2 => n483, ZN 
                           => n724);
   U827 : NAND3_X1 port map( A1 => n730, A2 => n731, A3 => n732, ZN => N584);
   U828 : AOI221_X1 port map( B1 => DATA1(21), B2 => n453, C1 => DATA1(19), C2 
                           => n454, A => n477, ZN => n732);
   U829 : MUX2_X1 port map( A => n733, B => n734, S => DATA1(20), Z => n731);
   U830 : NOR2_X1 port map( A1 => n455, A2 => n735, ZN => n734);
   U831 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(20), Z => n735);
   U832 : NAND2_X1 port map( A1 => DATA2(20), A2 => n481, ZN => n733);
   U833 : AOI22_X1 port map( A1 => N66, A2 => n464, B1 => N327, B2 => n483, ZN 
                           => n730);
   U834 : NAND3_X1 port map( A1 => n736, A2 => n737, A3 => n738, ZN => N583);
   U835 : AOI221_X1 port map( B1 => DATA1(20), B2 => n453, C1 => DATA1(18), C2 
                           => n454, A => n477, ZN => n738);
   U836 : MUX2_X1 port map( A => n739, B => n740, S => DATA1(19), Z => n737);
   U837 : NOR2_X1 port map( A1 => n455, A2 => n741, ZN => n740);
   U838 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(19), Z => n741);
   U839 : NAND2_X1 port map( A1 => DATA2(19), A2 => n481, ZN => n739);
   U840 : AOI22_X1 port map( A1 => N65, A2 => n464, B1 => N326, B2 => n483, ZN 
                           => n736);
   U841 : NAND3_X1 port map( A1 => n742, A2 => n743, A3 => n744, ZN => N582);
   U842 : AOI221_X1 port map( B1 => DATA1(19), B2 => n453, C1 => DATA1(17), C2 
                           => n454, A => n477, ZN => n744);
   U843 : MUX2_X1 port map( A => n745, B => n746, S => DATA1(18), Z => n743);
   U844 : NOR2_X1 port map( A1 => n455, A2 => n747, ZN => n746);
   U845 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(18), Z => n747);
   U846 : NAND2_X1 port map( A1 => DATA2(18), A2 => n481, ZN => n745);
   U847 : AOI22_X1 port map( A1 => N64, A2 => n464, B1 => N325, B2 => n483, ZN 
                           => n742);
   U848 : NAND3_X1 port map( A1 => n748, A2 => n749, A3 => n750, ZN => N581);
   U849 : AOI221_X1 port map( B1 => DATA1(18), B2 => n453, C1 => DATA1(16), C2 
                           => n454, A => n477, ZN => n750);
   U850 : MUX2_X1 port map( A => n751, B => n752, S => DATA1(17), Z => n749);
   U851 : NOR2_X1 port map( A1 => n455, A2 => n753, ZN => n752);
   U852 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(17), Z => n753);
   U853 : NAND2_X1 port map( A1 => DATA2(17), A2 => n481, ZN => n751);
   U854 : AOI22_X1 port map( A1 => N63, A2 => n464, B1 => N324, B2 => n483, ZN 
                           => n748);
   U855 : NAND3_X1 port map( A1 => n754, A2 => n755, A3 => n756, ZN => N580);
   U856 : AOI221_X1 port map( B1 => DATA1(17), B2 => n453, C1 => DATA1(15), C2 
                           => n454, A => n477, ZN => n756);
   U857 : MUX2_X1 port map( A => n757, B => n758, S => DATA1(16), Z => n755);
   U858 : NOR2_X1 port map( A1 => n455, A2 => n759, ZN => n758);
   U859 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(16), Z => n759);
   U860 : NAND2_X1 port map( A1 => DATA2(16), A2 => n481, ZN => n757);
   U861 : AOI22_X1 port map( A1 => N62, A2 => n464, B1 => N323, B2 => n483, ZN 
                           => n754);
   U862 : NAND3_X1 port map( A1 => n760, A2 => n761, A3 => n762, ZN => N579);
   U863 : AOI221_X1 port map( B1 => DATA1(16), B2 => n453, C1 => DATA1(14), C2 
                           => n454, A => n477, ZN => n762);
   U864 : MUX2_X1 port map( A => n763, B => n764, S => DATA1(15), Z => n761);
   U865 : NOR2_X1 port map( A1 => n455, A2 => n765, ZN => n764);
   U866 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(15), Z => n765);
   U867 : NAND2_X1 port map( A1 => DATA2(15), A2 => n481, ZN => n763);
   U868 : AOI22_X1 port map( A1 => N61, A2 => n464, B1 => N322, B2 => n483, ZN 
                           => n760);
   U869 : NAND3_X1 port map( A1 => n766, A2 => n767, A3 => n768, ZN => N578);
   U870 : AOI221_X1 port map( B1 => DATA1(15), B2 => n453, C1 => DATA1(13), C2 
                           => n454, A => n477, ZN => n768);
   U871 : MUX2_X1 port map( A => n769, B => n770, S => DATA1(14), Z => n767);
   U872 : NOR2_X1 port map( A1 => n455, A2 => n771, ZN => n770);
   U873 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(14), Z => n771);
   U874 : NAND2_X1 port map( A1 => DATA2(14), A2 => n481, ZN => n769);
   U875 : AOI22_X1 port map( A1 => N60, A2 => n464, B1 => N321, B2 => n483, ZN 
                           => n766);
   U876 : NAND3_X1 port map( A1 => n772, A2 => n773, A3 => n774, ZN => N577);
   U877 : AOI221_X1 port map( B1 => DATA1(14), B2 => n453, C1 => DATA1(12), C2 
                           => n454, A => n477, ZN => n774);
   U878 : MUX2_X1 port map( A => n775, B => n776, S => DATA1(13), Z => n773);
   U879 : NOR2_X1 port map( A1 => n455, A2 => n777, ZN => n776);
   U880 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(13), Z => n777);
   U881 : NAND2_X1 port map( A1 => DATA2(13), A2 => n481, ZN => n775);
   U882 : AOI22_X1 port map( A1 => N59, A2 => n464, B1 => N320, B2 => n483, ZN 
                           => n772);
   U883 : NAND3_X1 port map( A1 => n778, A2 => n779, A3 => n780, ZN => N576);
   U884 : AOI221_X1 port map( B1 => DATA1(13), B2 => n453, C1 => DATA1(11), C2 
                           => n454, A => n477, ZN => n780);
   U885 : MUX2_X1 port map( A => n781, B => n782, S => DATA1(12), Z => n779);
   U886 : NOR2_X1 port map( A1 => n455, A2 => n783, ZN => n782);
   U887 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(12), Z => n783);
   U888 : NAND2_X1 port map( A1 => DATA2(12), A2 => n481, ZN => n781);
   U889 : AOI22_X1 port map( A1 => N58, A2 => n464, B1 => N319, B2 => n483, ZN 
                           => n778);
   U890 : NAND3_X1 port map( A1 => n784, A2 => n785, A3 => n786, ZN => N575);
   U891 : AOI221_X1 port map( B1 => DATA1(12), B2 => n453, C1 => DATA1(10), C2 
                           => n454, A => n477, ZN => n786);
   U892 : MUX2_X1 port map( A => n787, B => n788, S => DATA1(11), Z => n785);
   U893 : NOR2_X1 port map( A1 => n455, A2 => n789, ZN => n788);
   U894 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(11), Z => n789);
   U895 : NAND2_X1 port map( A1 => DATA2(11), A2 => n481, ZN => n787);
   U896 : AOI22_X1 port map( A1 => N57, A2 => n464, B1 => N318, B2 => n483, ZN 
                           => n784);
   U897 : NAND3_X1 port map( A1 => n790, A2 => n791, A3 => n792, ZN => N574);
   U898 : AOI221_X1 port map( B1 => DATA1(11), B2 => n453, C1 => DATA1(9), C2 
                           => n454, A => n477, ZN => n792);
   U899 : MUX2_X1 port map( A => n793, B => n794, S => DATA1(10), Z => n791);
   U900 : NOR2_X1 port map( A1 => n455, A2 => n795, ZN => n794);
   U901 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(10), Z => n795);
   U902 : NAND2_X1 port map( A1 => DATA2(10), A2 => n481, ZN => n793);
   U903 : AOI22_X1 port map( A1 => N56, A2 => n464, B1 => N317, B2 => n483, ZN 
                           => n790);
   U904 : NAND3_X1 port map( A1 => n796, A2 => n797, A3 => n798, ZN => N573);
   U905 : AOI221_X1 port map( B1 => DATA1(10), B2 => n453, C1 => DATA1(8), C2 
                           => n454, A => n477, ZN => n798);
   U906 : MUX2_X1 port map( A => n799, B => n800, S => DATA1(9), Z => n797);
   U907 : NOR2_X1 port map( A1 => n455, A2 => n801, ZN => n800);
   U908 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(9), Z => n801);
   U909 : NAND2_X1 port map( A1 => DATA2(9), A2 => n481, ZN => n799);
   U910 : AOI22_X1 port map( A1 => N55, A2 => n464, B1 => N316, B2 => n483, ZN 
                           => n796);
   U911 : NAND3_X1 port map( A1 => n802, A2 => n803, A3 => n804, ZN => N572);
   U912 : AOI221_X1 port map( B1 => DATA1(9), B2 => n453, C1 => DATA1(7), C2 =>
                           n454, A => n477, ZN => n804);
   U913 : MUX2_X1 port map( A => n805, B => n806, S => DATA1(8), Z => n803);
   U914 : NOR2_X1 port map( A1 => n455, A2 => n807, ZN => n806);
   U915 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(8), Z => n807);
   U916 : NAND2_X1 port map( A1 => DATA2(8), A2 => n481, ZN => n805);
   U917 : AOI22_X1 port map( A1 => N54, A2 => n464, B1 => N315, B2 => n483, ZN 
                           => n802);
   U918 : NAND3_X1 port map( A1 => n808, A2 => n809, A3 => n810, ZN => N571);
   U919 : AOI221_X1 port map( B1 => DATA1(8), B2 => n453, C1 => DATA1(6), C2 =>
                           n454, A => n477, ZN => n810);
   U920 : MUX2_X1 port map( A => n811, B => n812, S => DATA1(7), Z => n809);
   U921 : NOR2_X1 port map( A1 => n455, A2 => n813, ZN => n812);
   U922 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(7), Z => n813);
   U923 : NAND2_X1 port map( A1 => DATA2(7), A2 => n481, ZN => n811);
   U924 : AOI22_X1 port map( A1 => N53, A2 => n464, B1 => N314, B2 => n483, ZN 
                           => n808);
   U925 : NAND3_X1 port map( A1 => n814, A2 => n815, A3 => n816, ZN => N570);
   U926 : AOI221_X1 port map( B1 => DATA1(7), B2 => n453, C1 => DATA1(5), C2 =>
                           n454, A => n477, ZN => n816);
   U927 : MUX2_X1 port map( A => n817, B => n818, S => DATA1(6), Z => n815);
   U928 : NOR2_X1 port map( A1 => n455, A2 => n819, ZN => n818);
   U929 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(6), Z => n819);
   U930 : NAND2_X1 port map( A1 => DATA2(6), A2 => n481, ZN => n817);
   U931 : AOI22_X1 port map( A1 => N52, A2 => n464, B1 => N313, B2 => n483, ZN 
                           => n814);
   U932 : NAND3_X1 port map( A1 => n820, A2 => n821, A3 => n822, ZN => N569);
   U933 : AOI221_X1 port map( B1 => DATA1(6), B2 => n453, C1 => DATA1(4), C2 =>
                           n454, A => n477, ZN => n822);
   U934 : MUX2_X1 port map( A => n823, B => n824, S => DATA1(5), Z => n821);
   U935 : NOR2_X1 port map( A1 => n455, A2 => n825, ZN => n824);
   U936 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(5), Z => n825);
   U937 : NAND2_X1 port map( A1 => DATA2(5), A2 => n481, ZN => n823);
   U938 : AOI22_X1 port map( A1 => N51, A2 => n464, B1 => N312, B2 => n483, ZN 
                           => n820);
   U939 : NAND3_X1 port map( A1 => n826, A2 => n827, A3 => n828, ZN => N568);
   U940 : AOI221_X1 port map( B1 => DATA1(5), B2 => n453, C1 => DATA1(3), C2 =>
                           n454, A => n477, ZN => n828);
   U941 : MUX2_X1 port map( A => n829, B => n830, S => DATA1(4), Z => n827);
   U942 : NOR2_X1 port map( A1 => n455, A2 => n831, ZN => n830);
   U943 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(4), Z => n831);
   U944 : NAND2_X1 port map( A1 => DATA2(4), A2 => n481, ZN => n829);
   U945 : AOI22_X1 port map( A1 => N50, A2 => n464, B1 => N311, B2 => n483, ZN 
                           => n826);
   U946 : NAND3_X1 port map( A1 => n832, A2 => n833, A3 => n834, ZN => N567);
   U947 : AOI221_X1 port map( B1 => DATA1(4), B2 => n453, C1 => DATA1(2), C2 =>
                           n454, A => n477, ZN => n834);
   U948 : MUX2_X1 port map( A => n835, B => n836, S => DATA1(3), Z => n833);
   U949 : NOR2_X1 port map( A1 => n455, A2 => n837, ZN => n836);
   U950 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(3), Z => n837);
   U951 : NAND2_X1 port map( A1 => DATA2(3), A2 => n481, ZN => n835);
   U952 : AOI22_X1 port map( A1 => N49, A2 => n464, B1 => N310, B2 => n483, ZN 
                           => n832);
   U953 : NAND3_X1 port map( A1 => n838, A2 => n839, A3 => n840, ZN => N566);
   U954 : AOI221_X1 port map( B1 => DATA1(3), B2 => n453, C1 => DATA1(1), C2 =>
                           n454, A => n477, ZN => n840);
   U955 : MUX2_X1 port map( A => n841, B => n842, S => DATA1(2), Z => n839);
   U956 : NOR2_X1 port map( A1 => n455, A2 => n843, ZN => n842);
   U957 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(2), Z => n843);
   U958 : NAND2_X1 port map( A1 => DATA2(2), A2 => n481, ZN => n841);
   U959 : AOI22_X1 port map( A1 => N48, A2 => n464, B1 => N309, B2 => n483, ZN 
                           => n838);
   U960 : NAND3_X1 port map( A1 => n844, A2 => n845, A3 => n846, ZN => N565);
   U961 : AOI221_X1 port map( B1 => DATA1(2), B2 => n453, C1 => n454, C2 => 
                           DATA1(0), A => n477, ZN => n846);
   U962 : MUX2_X1 port map( A => n848, B => n849, S => DATA1(1), Z => n845);
   U963 : NOR2_X1 port map( A1 => n455, A2 => n850, ZN => n849);
   U964 : MUX2_X1 port map( A => n481, B => n482, S => DATA2(1), Z => n850);
   U965 : NAND2_X1 port map( A1 => DATA2(1), A2 => n481, ZN => n848);
   U966 : AOI22_X1 port map( A1 => N47, A2 => n464, B1 => N308, B2 => n483, ZN 
                           => n844);
   U967 : NAND4_X1 port map( A1 => n853, A2 => n854, A3 => n855, A4 => n462, ZN
                           => N564);
   U968 : NAND4_X1 port map( A1 => N110, A2 => n856, A3 => n458, A4 => n857, ZN
                           => n462);
   U969 : NAND3_X1 port map( A1 => FUNC_0_port, A2 => n463, A3 => DATA1(1), ZN 
                           => n855);
   U970 : OAI21_X1 port map( B1 => n468, B2 => n858, A => n859, ZN => n463);
   U971 : NAND2_X1 port map( A1 => N46, A2 => n464, ZN => n854);
   U972 : MUX2_X1 port map( A => n860, B => n861, S => FUNC_2_port, Z => n853);
   U973 : NAND2_X1 port map( A1 => n862, A2 => n468, ZN => n861);
   U974 : MUX2_X1 port map( A => DATA1(0), B => n863, S => DATA2(0), Z => n862)
                           ;
   U975 : NAND2_X1 port map( A1 => DATA1(0), A2 => FUNC_0_port, ZN => n863);
   U976 : AOI21_X1 port map( B1 => N307, B2 => n471, A => n864, ZN => n860);
   U977 : MUX2_X1 port map( A => n865, B => n866, S => FUNC_1_port, Z => n864);
   U978 : AND3_X1 port map( A1 => DATA2(0), A2 => FUNC_0_port, A3 => DATA1(0), 
                           ZN => n866);
   U979 : AND3_X1 port map( A1 => DATA1(63), A2 => n458, A3 => FUNC_3_port, ZN 
                           => n865);
   U980 : INV_X1 port map( A => FUNC_0_port, ZN => n458);
   U981 : NAND3_X1 port map( A1 => n468, A2 => n857, A3 => FUNC_2_port, ZN => 
                           n852);
   U982 : NOR2_X1 port map( A1 => n483, A2 => n856, ZN => n867);
   U983 : NOR2_X1 port map( A1 => n468, A2 => FUNC_0_port, ZN => n471);
   U984 : NAND4_X1 port map( A1 => FUNC_1_port, A2 => FUNC_0_port, A3 => n858, 
                           A4 => n857, ZN => n851);
   U985 : AND2_X1 port map( A1 => n859, A2 => n868, ZN => n847);
   U986 : NAND3_X1 port map( A1 => FUNC_1_port, A2 => n857, A3 => FUNC_2_port, 
                           ZN => n868);
   U987 : INV_X1 port map( A => FUNC_3_port, ZN => n857);
   U988 : NAND2_X1 port map( A1 => FUNC_3_port, A2 => n856, ZN => n859);
   U989 : INV_X1 port map( A => n457, ZN => n856);
   U990 : NAND2_X1 port map( A1 => n468, A2 => n858, ZN => n457);
   U991 : INV_X1 port map( A => FUNC_2_port, ZN => n858);
   U992 : INV_X1 port map( A => FUNC_1_port, ZN => n468);

end SYN_BEHAVIOR_1;
