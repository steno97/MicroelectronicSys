
module windRF_M8_N8_F2_NBIT64 ( CLK, RESET, ENABLE, CALL, RETRN, FILL, SPILL, 
        BUSin, BUSout, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, 
        OUT2 );
  input [63:0] BUSin;
  output [63:0] BUSout;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, CALL, RETRN, RD1, RD2, WR;
  output FILL, SPILL;
  wire   \i[3] , \i[2] , \i[1] , N659, N660, N661, N688, N689, N690, N811,
         N812, N813, N929, N930, N931, N932, N6270, N6271, N6272, N6273, N6395,
         N6396, N6397, N6398, \U3/U193/Z_1 , \U3/U193/Z_2 , \U3/U193/Z_3 ,
         \U3/U193/Z_4 , \U3/U194/Z_1 , \U3/U194/Z_2 , \U3/U194/Z_3 ,
         \U3/U194/Z_4 , \U3/U195/Z_1 , \U3/U195/Z_2 , \U3/U195/Z_3 ,
         \U3/U195/Z_4 , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n2683, n2695, n2696, n2697, n2698, n2699,
         n2700, n2706, n2707, n2709, n2710, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, \add_146/carry[4] , \add_146/carry[3] ,
         \add_146/carry[2] , n12791, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n23853, n25394, \r510/n3 , \r510/carry[5] ,
         \r510/carry[4] , \r510/carry[3] , \r510/carry[2] , \r504/n3 ,
         \r504/carry[5] , \r504/carry[4] , \r504/carry[3] , \r504/carry[2] ,
         \r498/n1 , \r498/carry[5] , \r498/carry[4] , \r498/carry[3] ,
         \r498/carry[2] , \add_136/carry[2] , \add_136/carry[3] ,
         \add_136/carry[4] , n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n27870,
         n27871, n27872, n27874, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
         n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
         n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
         n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
         n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28840, n28841, n28842, n28843, n28844, n28845,
         n28846, n28847, n28848, n28849, n28850, n29043, n29044, n29045,
         n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
         n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061,
         n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069,
         n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
         n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085,
         n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
         n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
         n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109,
         n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117,
         n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
         n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
         n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
         n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149,
         n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157,
         n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
         n29166, n29167, n29168, n29169, n29170, n29363, n29364, n29365,
         n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373,
         n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381,
         n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389,
         n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397,
         n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405,
         n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
         n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
         n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
         n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
         n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
         n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453,
         n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461,
         n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469,
         n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
         n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
         n29486, n29487, n29488, n29489, n29490, n29683, n29684, n29685,
         n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693,
         n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
         n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709,
         n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
         n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
         n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733,
         n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
         n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749,
         n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757,
         n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765,
         n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
         n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781,
         n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
         n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797,
         n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805,
         n29806, n29807, n29808, n29809, n29810, n30003, n30004, n30005,
         n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013,
         n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021,
         n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029,
         n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037,
         n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045,
         n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053,
         n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
         n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069,
         n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077,
         n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085,
         n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093,
         n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101,
         n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109,
         n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117,
         n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125,
         n30126, n30127, n30128, n30129, n30130, n30458, n30459, n30460,
         n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468,
         n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476,
         n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
         n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492,
         n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
         n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
         n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516,
         n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
         n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
         n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
         n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548,
         n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
         n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564,
         n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572,
         n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580,
         n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588,
         n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
         n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604,
         n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612,
         n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620,
         n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
         n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636,
         n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644,
         n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652,
         n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660,
         n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
         n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676,
         n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684,
         n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692,
         n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
         n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708,
         n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716,
         n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724,
         n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732,
         n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740,
         n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
         n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756,
         n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764,
         n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
         n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780,
         n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
         n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796,
         n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804,
         n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812,
         n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820,
         n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828,
         n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836,
         n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
         n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852,
         n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860,
         n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868,
         n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876,
         n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884,
         n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892,
         n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900,
         n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908,
         n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
         n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924,
         n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
         n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940,
         n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948,
         n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956,
         n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964,
         n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972,
         n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980,
         n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
         n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996,
         n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
         n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012,
         n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020,
         n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028,
         n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
         n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
         n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052,
         n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
         n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068,
         n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
         n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
         n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
         n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
         n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
         n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
         n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124,
         n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
         n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140,
         n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
         n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
         n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164,
         n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
         n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
         n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188,
         n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196,
         n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
         n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212,
         n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
         n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
         n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236,
         n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244,
         n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
         n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260,
         n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
         n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
         n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284,
         n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
         n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
         n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308,
         n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
         n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324,
         n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332,
         n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340,
         n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
         n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
         n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
         n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
         n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380,
         n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
         n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
         n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428,
         n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
         n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
         n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452,
         n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
         n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
         n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476,
         n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484,
         n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
         n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500,
         n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
         n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516,
         n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524,
         n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
         n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
         n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548,
         n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
         n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
         n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
         n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
         n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
         n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596,
         n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
         n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
         n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
         n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
         n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
         n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644,
         n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
         n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
         n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668,
         n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
         n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
         n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
         n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
         n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
         n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
         n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740,
         n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
         n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
         n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764,
         n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
         n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
         n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
         n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
         n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
         n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
         n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
         n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
         n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
         n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
         n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
         n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
         n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
         n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
         n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
         n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908,
         n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
         n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
         n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
         n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
         n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
         n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
         n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
         n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
         n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980,
         n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
         n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
         n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
         n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
         n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
         n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
         n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
         n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052,
         n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
         n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
         n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
         n32077, n32079, n32080, n32081, n32082, n32083, n32084, n32085,
         n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
         n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101,
         n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109,
         n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117,
         n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125,
         n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133,
         n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141,
         n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149,
         n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157,
         n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165,
         n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173,
         n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181,
         n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189,
         n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197,
         n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205,
         n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213,
         n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221,
         n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229,
         n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237,
         n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32246,
         n32247, n32248, n32249, n32251, n32253, n32254, n32255, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32384, n32444, n32456, n32457, n32458, n32459, n32460,
         n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
         n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
         n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484,
         n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946,
         n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
         n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
         n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
         n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
         n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
         n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994,
         n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
         n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
         n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018,
         n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33087, n33088, n33089, n33090,
         n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
         n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
         n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
         n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122,
         n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
         n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33139,
         n33195, n33196, n33197, n33199, n33207, n33208, n33209, n33210,
         n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
         n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
         n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234,
         n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
         n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
         n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258,
         n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266,
         n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
         n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282,
         n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
         n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
         n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
         n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
         n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
         n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
         n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
         n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
         n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354,
         n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
         n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
         n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378,
         n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
         n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410,
         n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
         n33419, n33420, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155,
         n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
         n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
         n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
         n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
         n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203,
         n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211,
         n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
         n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
         n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
         n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
         n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419,
         n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
         n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443,
         n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
         n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
         n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467,
         n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
         n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
         n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491,
         n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
         n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
         n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515,
         n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
         n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
         n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539,
         n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
         n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
         n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563,
         n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
         n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587,
         n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
         n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
         n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
         n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
         n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
         n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635,
         n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
         n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
         n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659,
         n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
         n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
         n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
         n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731,
         n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
         n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
         n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
         n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
         n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
         n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
         n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
         n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
         n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
         n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
         n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
         n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827,
         n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
         n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
         n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851,
         n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
         n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
         n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
         n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
         n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
         n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899,
         n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
         n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
         n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923,
         n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931,
         n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
         n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
         n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
         n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003,
         n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
         n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
         n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
         n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
         n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
         n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
         n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
         n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075,
         n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
         n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
         n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115,
         n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
         n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
         n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
         n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147,
         n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
         n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
         n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
         n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
         n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187,
         n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
         n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
         n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
         n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219,
         n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
         n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
         n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259,
         n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
         n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
         n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
         n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291,
         n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
         n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
         n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331,
         n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
         n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
         n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363,
         n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
         n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379,
         n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
         n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
         n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403,
         n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
         n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
         n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435,
         n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
         n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451,
         n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
         n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
         n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
         n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
         n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499,
         n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
         n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
         n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
         n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
         n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
         n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595,
         n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
         n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
         n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619,
         n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
         n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
         n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643,
         n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
         n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
         n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667,
         n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
         n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
         n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
         n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
         n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
         n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715,
         n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
         n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
         n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739,
         n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
         n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
         n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787,
         n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
         n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
         n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811,
         n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
         n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
         n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835,
         n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
         n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
         n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883,
         n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
         n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
         n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
         n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931,
         n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
         n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
         n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955,
         n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
         n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
         n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
         n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011,
         n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
         n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027,
         n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
         n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
         n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083,
         n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
         n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099,
         n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
         n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
         n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
         n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
         n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
         n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155,
         n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
         n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171,
         n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195,
         n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
         n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
         n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
         n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227,
         n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
         n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243,
         n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
         n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
         n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267,
         n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
         n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299,
         n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
         n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
         n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
         n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
         n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339,
         n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
         n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
         n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363,
         n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371,
         n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
         n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
         n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
         n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
         n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411,
         n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
         n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
         n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
         n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
         n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483,
         n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
         n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507,
         n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515,
         n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
         n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
         n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
         n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
         n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
         n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
         n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579,
         n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
         n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
         n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
         n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627,
         n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
         n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
         n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
         n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
         n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
         n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
         n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
         n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
         n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
         n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
         n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
         n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
         n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
         n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
         n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
         n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
         n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
         n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
         n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
         n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
         n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
         n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
         n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
         n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
         n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867,
         n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875,
         n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
         n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891,
         n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
         n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
         n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
         n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
         n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811,
         n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819,
         n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
         n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835,
         n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
         n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851,
         n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859,
         n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
         n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875,
         n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883,
         n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891,
         n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
         n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907,
         n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
         n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
         n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931,
         n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939,
         n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947,
         n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955,
         n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963,
         n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
         n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979,
         n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
         n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
         n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003,
         n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
         n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019,
         n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027,
         n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035,
         n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
         n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051,
         n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
         n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067,
         n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075,
         n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
         n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091,
         n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099,
         n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107,
         n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
         n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123,
         n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
         n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139,
         n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147,
         n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
         n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163,
         n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
         n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
         n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
         n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195,
         n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
         n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211,
         n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219,
         n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227,
         n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235,
         n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243,
         n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
         n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
         n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267,
         n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
         n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283,
         n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291,
         n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299,
         n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307,
         n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
         n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
         n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
         n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339,
         n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
         n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
         n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363,
         n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371,
         n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379,
         n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387,
         n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395,
         n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
         n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411,
         n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
         n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427,
         n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435,
         n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
         n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451,
         n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459,
         n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467,
         n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
         n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483,
         n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
         n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
         n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
         n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
         n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523,
         n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531,
         n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
         n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
         n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555,
         n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
         n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
         n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579,
         n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
         n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595,
         n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
         n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
         n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
         n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
         n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
         n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
         n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651,
         n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659,
         n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667,
         n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675,
         n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683,
         n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
         n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699,
         n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
         n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715,
         n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
         n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731,
         n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739,
         n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747,
         n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755,
         n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
         n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771,
         n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
         n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
         n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795,
         n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803,
         n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811,
         n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
         n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827,
         n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
         n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843,
         n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
         n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859,
         n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867,
         n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
         n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883,
         n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891,
         n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899,
         n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
         n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915,
         n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
         n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931,
         n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
         n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947,
         n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955,
         n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963,
         n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971,
         n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
         n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987,
         n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
         n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
         n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011,
         n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019,
         n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027,
         n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035,
         n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043,
         n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
         n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059,
         n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
         n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075,
         n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083,
         n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091,
         n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
         n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107,
         n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115,
         n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
         n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131,
         n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
         n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147,
         n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155,
         n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163,
         n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171,
         n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179,
         n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187,
         n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
         n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203,
         n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
         n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219,
         n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227,
         n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235,
         n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243,
         n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251,
         n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259,
         n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
         n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275,
         n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
         n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291,
         n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299,
         n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307,
         n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315,
         n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323,
         n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331,
         n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
         n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347,
         n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
         n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
         n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371,
         n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379,
         n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387,
         n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395,
         n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403,
         n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
         n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419,
         n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
         n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
         n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443,
         n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451,
         n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459,
         n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467,
         n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
         n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
         n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
         n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
         n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
         n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515,
         n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
         n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
         n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
         n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
         n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
         n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
         n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
         n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
         n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
         n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
         n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
         n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
         n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
         n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
         n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
         n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
         n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
         n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
         n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
         n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675,
         n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
         n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
         n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
         n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731,
         n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
         n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
         n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755,
         n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
         n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
         n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779,
         n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
         n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
         n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803,
         n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
         n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819,
         n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
         n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835,
         n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
         n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851,
         n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
         n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
         n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875,
         n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
         n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891,
         n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
         n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
         n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923,
         n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
         n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
         n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
         n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
         n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963,
         n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971,
         n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
         n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
         n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995,
         n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
         n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
         n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019,
         n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
         n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035,
         n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043,
         n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
         n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
         n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091,
         n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
         n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
         n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
         n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
         n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163,
         n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
         n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179,
         n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
         n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
         n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
         n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211,
         n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
         n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
         n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235,
         n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
         n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
         n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259,
         n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267,
         n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
         n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283,
         n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
         n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
         n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307,
         n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
         n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339,
         n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
         n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355,
         n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
         n41364, n41365, n41366, n41367, n41368, n41369, n41370;

  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n7459), .CK(CLK), .QN(n30481) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n7460), .CK(CLK), .QN(n30482) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n7461), .CK(CLK), .QN(n30483) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n7462), .CK(CLK), .QN(n30484) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n7463), .CK(CLK), .QN(n30485) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n7464), .CK(CLK), .QN(n30486) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n7465), .CK(CLK), .QN(n30487) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n7466), .CK(CLK), .QN(n30488) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n7467), .CK(CLK), .QN(n30489) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n7468), .CK(CLK), .QN(n30490) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n7469), .CK(CLK), .QN(n30491) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n7470), .CK(CLK), .QN(n30492) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n7471), .CK(CLK), .QN(n30493) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n7472), .CK(CLK), .QN(n30494) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n7473), .CK(CLK), .QN(n30495) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n7474), .CK(CLK), .QN(n30496) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n7475), .CK(CLK), .QN(n30497) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n7476), .CK(CLK), .QN(n30498) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n7477), .CK(CLK), .QN(n30499) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n7478), .CK(CLK), .QN(n30500) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n7479), .CK(CLK), .QN(n30501) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n7480), .CK(CLK), .QN(n30502) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n7481), .CK(CLK), .QN(n30503) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n7482), .CK(CLK), .QN(n30504) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n7483), .CK(CLK), .QN(n30505) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n7484), .CK(CLK), .QN(n30506) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n7485), .CK(CLK), .QN(n30507) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n7486), .CK(CLK), .QN(n30508) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n7487), .CK(CLK), .QN(n30509) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n7488), .CK(CLK), .QN(n30510) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n7489), .CK(CLK), .QN(n30511) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n7490), .CK(CLK), .QN(n30512) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n7491), .CK(CLK), .QN(n30513) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n7492), .CK(CLK), .QN(n30514) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n7493), .CK(CLK), .QN(n30515) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n7494), .CK(CLK), .QN(n30516) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n7495), .CK(CLK), .QN(n30517) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n7496), .CK(CLK), .QN(n30518) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n7497), .CK(CLK), .QN(n30519) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n7498), .CK(CLK), .QN(n30520) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n7499), .CK(CLK), .QN(n30521) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n7500), .CK(CLK), .QN(n30522) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n7501), .CK(CLK), .QN(n30523) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n7502), .CK(CLK), .QN(n30524) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n7503), .CK(CLK), .QN(n30525) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n7504), .CK(CLK), .QN(n30526) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n7505), .CK(CLK), .QN(n30527) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n7506), .CK(CLK), .QN(n30528) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n7507), .CK(CLK), .QN(n30529) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n7508), .CK(CLK), .QN(n30530) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n7509), .CK(CLK), .QN(n30531) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n7510), .CK(CLK), .QN(n30532) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n7511), .CK(CLK), .QN(n30533) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n7512), .CK(CLK), .QN(n30534) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n7513), .CK(CLK), .QN(n30535) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n7514), .CK(CLK), .QN(n30536) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n7515), .CK(CLK), .QN(n30537) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n7516), .CK(CLK), .QN(n30538) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n7517), .CK(CLK), .QN(n30539) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n7518), .CK(CLK), .QN(n30540) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n7523), .CK(CLK), .QN(n30545) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n7524), .CK(CLK), .QN(n30546) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n7525), .CK(CLK), .QN(n30547) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n7527), .CK(CLK), .QN(n30549) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n7547), .CK(CLK), .QN(n30569) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n7548), .CK(CLK), .QN(n30570) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n7549), .CK(CLK), .QN(n30571) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n7550), .CK(CLK), .QN(n30572) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n7551), .CK(CLK), .QN(n30573) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n7552), .CK(CLK), .QN(n30574) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n7553), .CK(CLK), .QN(n30575) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n7554), .CK(CLK), .QN(n30576) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n7555), .CK(CLK), .QN(n30577) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n7556), .CK(CLK), .QN(n30578) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n7557), .CK(CLK), .QN(n30579) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n7558), .CK(CLK), .QN(n30580) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n7559), .CK(CLK), .QN(n30581) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n7560), .CK(CLK), .QN(n30582) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n7561), .CK(CLK), .QN(n30583) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n7562), .CK(CLK), .QN(n30584) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n7563), .CK(CLK), .QN(n30585) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n7564), .CK(CLK), .QN(n30586) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n7565), .CK(CLK), .QN(n30587) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n7566), .CK(CLK), .QN(n30588) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n7567), .CK(CLK), .QN(n30589) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n7568), .CK(CLK), .QN(n30590) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n7569), .CK(CLK), .QN(n30591) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n7570), .CK(CLK), .QN(n30592) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n7571), .CK(CLK), .QN(n30593) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n7572), .CK(CLK), .QN(n30594) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n7573), .CK(CLK), .QN(n30595) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n7574), .CK(CLK), .QN(n30596) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n7575), .CK(CLK), .QN(n30597) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n7576), .CK(CLK), .QN(n30598) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n7577), .CK(CLK), .QN(n30599) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n7578), .CK(CLK), .QN(n30600) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n7579), .CK(CLK), .QN(n30601) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n7580), .CK(CLK), .QN(n30602) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n7581), .CK(CLK), .QN(n30603) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n7582), .CK(CLK), .QN(n30604) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n7587), .CK(CLK), .QN(n30609) );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n7588), .CK(CLK), .QN(n30610) );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n7589), .CK(CLK), .QN(n30611) );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n7590), .CK(CLK), .QN(n30612) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n7591), .CK(CLK), .QN(n30613) );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n7592), .CK(CLK), .QN(n30614) );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n7593), .CK(CLK), .QN(n30615) );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n7594), .CK(CLK), .QN(n30616) );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n7595), .CK(CLK), .QN(n30617) );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n7596), .CK(CLK), .QN(n30618) );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n7597), .CK(CLK), .QN(n30619) );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n7598), .CK(CLK), .QN(n30620) );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n7599), .CK(CLK), .QN(n30621) );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n7600), .CK(CLK), .QN(n30622) );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n7601), .CK(CLK), .QN(n30623) );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n7602), .CK(CLK), .QN(n30624) );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n7603), .CK(CLK), .QN(n30625) );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n7604), .CK(CLK), .QN(n30626) );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n7605), .CK(CLK), .QN(n30627) );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n7606), .CK(CLK), .QN(n30628) );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n7607), .CK(CLK), .QN(n30629) );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n7608), .CK(CLK), .QN(n30630) );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n7609), .CK(CLK), .QN(n30631) );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n7610), .CK(CLK), .QN(n30632) );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n7611), .CK(CLK), .QN(n30633) );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n7612), .CK(CLK), .QN(n30634) );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n7613), .CK(CLK), .QN(n30635) );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n7614), .CK(CLK), .QN(n30636) );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n7615), .CK(CLK), .QN(n30637) );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n7616), .CK(CLK), .QN(n30638) );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n7617), .CK(CLK), .QN(n30639) );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n7618), .CK(CLK), .QN(n30640) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n7619), .CK(CLK), .QN(n30641) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n7620), .CK(CLK), .QN(n30642) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n7621), .CK(CLK), .QN(n30643) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n7622), .CK(CLK), .QN(n30644) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n7623), .CK(CLK), .QN(n30645) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n7624), .CK(CLK), .QN(n30646) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n7625), .CK(CLK), .QN(n30647) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n7626), .CK(CLK), .QN(n30648) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n7627), .CK(CLK), .QN(n30649) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n7628), .CK(CLK), .QN(n30650) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n7629), .CK(CLK), .QN(n30651) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n7630), .CK(CLK), .QN(n30652) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n7631), .CK(CLK), .QN(n30653) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n7632), .CK(CLK), .QN(n30654) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n7633), .CK(CLK), .QN(n30655) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n7634), .CK(CLK), .QN(n30656) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n7635), .CK(CLK), .QN(n30657) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n7636), .CK(CLK), .QN(n30658) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n7637), .CK(CLK), .QN(n30659) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n7638), .CK(CLK), .QN(n30660) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n7639), .CK(CLK), .QN(n30661) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n7640), .CK(CLK), .QN(n30662) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n7641), .CK(CLK), .QN(n30663) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n7642), .CK(CLK), .QN(n30664) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n7643), .CK(CLK), .QN(n30665) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n7644), .CK(CLK), .QN(n30666) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n7645), .CK(CLK), .QN(n30667) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n7646), .CK(CLK), .QN(n30668) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n7779), .CK(CLK), .QN(n30673) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n7780), .CK(CLK), .QN(n30674) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n7781), .CK(CLK), .QN(n30675) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n7782), .CK(CLK), .QN(n30676) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n7783), .CK(CLK), .QN(n30677) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n7784), .CK(CLK), .QN(n30678) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n7785), .CK(CLK), .QN(n30679) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n7786), .CK(CLK), .QN(n30680) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n7787), .CK(CLK), .QN(n30681) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n7788), .CK(CLK), .QN(n30682) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n7789), .CK(CLK), .QN(n30683) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n7790), .CK(CLK), .QN(n30684) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n7791), .CK(CLK), .QN(n30685) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n7792), .CK(CLK), .QN(n30686) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n7793), .CK(CLK), .QN(n30687) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n7794), .CK(CLK), .QN(n30688) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n7795), .CK(CLK), .QN(n30689) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n7796), .CK(CLK), .QN(n30690) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n7797), .CK(CLK), .QN(n30691) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n7798), .CK(CLK), .QN(n30692) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n7799), .CK(CLK), .QN(n30693) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n7800), .CK(CLK), .QN(n30694) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n7801), .CK(CLK), .QN(n30695) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n7802), .CK(CLK), .QN(n30696) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n7803), .CK(CLK), .QN(n30697) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n7804), .CK(CLK), .QN(n30698) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n7805), .CK(CLK), .QN(n30699) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n7806), .CK(CLK), .QN(n30700) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n7807), .CK(CLK), .QN(n30701) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n7808), .CK(CLK), .QN(n30702) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n7809), .CK(CLK), .QN(n30703) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n7810), .CK(CLK), .QN(n30704) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n7811), .CK(CLK), .QN(n30705) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n7812), .CK(CLK), .QN(n30706) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n7813), .CK(CLK), .QN(n30707) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n7814), .CK(CLK), .QN(n30708) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n7815), .CK(CLK), .QN(n30709) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n7816), .CK(CLK), .QN(n30710) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n7817), .CK(CLK), .QN(n30711) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n7818), .CK(CLK), .QN(n30712) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n7819), .CK(CLK), .QN(n30713) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n7820), .CK(CLK), .QN(n30714) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n7821), .CK(CLK), .QN(n30715) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n7822), .CK(CLK), .QN(n30716) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n7823), .CK(CLK), .QN(n30717) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n7824), .CK(CLK), .QN(n30718) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n7825), .CK(CLK), .QN(n30719) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n7826), .CK(CLK), .QN(n30720) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n7827), .CK(CLK), .QN(n30721) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n7828), .CK(CLK), .QN(n30722) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n7829), .CK(CLK), .QN(n30723) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n7830), .CK(CLK), .QN(n30724) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n7831), .CK(CLK), .QN(n30725) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n7832), .CK(CLK), .QN(n30726) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n7833), .CK(CLK), .QN(n30727) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n7834), .CK(CLK), .QN(n30728) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n7835), .CK(CLK), .QN(n30729) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n7836), .CK(CLK), .QN(n30730) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n7837), .CK(CLK), .QN(n30731) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n7838), .CK(CLK), .QN(n30732) );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n7843), .CK(CLK), .QN(n30737) );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n7844), .CK(CLK), .QN(n30738) );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n7845), .CK(CLK), .QN(n30739) );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n7846), .CK(CLK), .QN(n30740) );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n7847), .CK(CLK), .QN(n30741) );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n7848), .CK(CLK), .QN(n30742) );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n7849), .CK(CLK), .QN(n30743) );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n7850), .CK(CLK), .QN(n30744) );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n7851), .CK(CLK), .QN(n30745) );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n7852), .CK(CLK), .QN(n30746) );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n7853), .CK(CLK), .QN(n30747) );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n7854), .CK(CLK), .QN(n30748) );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n7855), .CK(CLK), .QN(n30749) );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n7856), .CK(CLK), .QN(n30750) );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n7857), .CK(CLK), .QN(n30751) );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n7858), .CK(CLK), .QN(n30752) );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n7859), .CK(CLK), .QN(n30753) );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n7860), .CK(CLK), .QN(n30754) );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n7861), .CK(CLK), .QN(n30755) );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n7862), .CK(CLK), .QN(n30756) );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n7863), .CK(CLK), .QN(n30757) );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n7864), .CK(CLK), .QN(n30758) );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n7865), .CK(CLK), .QN(n30759) );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n7866), .CK(CLK), .QN(n30760) );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n7867), .CK(CLK), .QN(n30761) );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n7868), .CK(CLK), .QN(n30762) );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n7869), .CK(CLK), .QN(n30763) );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n7870), .CK(CLK), .QN(n30764) );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n7871), .CK(CLK), .QN(n30765) );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n7872), .CK(CLK), .QN(n30766) );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n7873), .CK(CLK), .QN(n30767) );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n7874), .CK(CLK), .QN(n30768) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n7875), .CK(CLK), .QN(n30769) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n7876), .CK(CLK), .QN(n30770) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n7877), .CK(CLK), .QN(n30771) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n7878), .CK(CLK), .QN(n30772) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n7879), .CK(CLK), .QN(n30773) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n7880), .CK(CLK), .QN(n30774) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n7881), .CK(CLK), .QN(n30775) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n7882), .CK(CLK), .QN(n30776) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n7883), .CK(CLK), .QN(n30777) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n7884), .CK(CLK), .QN(n30778) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n7885), .CK(CLK), .QN(n30779) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n7886), .CK(CLK), .QN(n30780) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n7887), .CK(CLK), .QN(n30781) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n7888), .CK(CLK), .QN(n30782) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n7889), .CK(CLK), .QN(n30783) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n7890), .CK(CLK), .QN(n30784) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n7891), .CK(CLK), .QN(n30785) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n7892), .CK(CLK), .QN(n30786) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n7893), .CK(CLK), .QN(n30787) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n7894), .CK(CLK), .QN(n30788) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n7895), .CK(CLK), .QN(n30789) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n7896), .CK(CLK), .QN(n30790) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n7897), .CK(CLK), .QN(n30791) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n7898), .CK(CLK), .QN(n30792) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n7899), .CK(CLK), .QN(n30793) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n7900), .CK(CLK), .QN(n30794) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n7901), .CK(CLK), .QN(n30795) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n7902), .CK(CLK), .QN(n30796) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n7907), .CK(CLK), .QN(n30801) );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n7908), .CK(CLK), .QN(n30802) );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n7909), .CK(CLK), .QN(n30803) );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n7910), .CK(CLK), .QN(n30804) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n7911), .CK(CLK), .QN(n30805) );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n7912), .CK(CLK), .QN(n30806) );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n7913), .CK(CLK), .QN(n30807) );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n7914), .CK(CLK), .QN(n30808) );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n7915), .CK(CLK), .QN(n30809) );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n7916), .CK(CLK), .QN(n30810) );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n7917), .CK(CLK), .QN(n30811) );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n7918), .CK(CLK), .QN(n30812) );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n7919), .CK(CLK), .QN(n30813) );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n7920), .CK(CLK), .QN(n30814) );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n7921), .CK(CLK), .QN(n30815) );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n7922), .CK(CLK), .QN(n30816) );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n7923), .CK(CLK), .QN(n30817) );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n7924), .CK(CLK), .QN(n30818) );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n7925), .CK(CLK), .QN(n30819) );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n7926), .CK(CLK), .QN(n30820) );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n7927), .CK(CLK), .QN(n30821) );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n7928), .CK(CLK), .QN(n30822) );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n7929), .CK(CLK), .QN(n30823) );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n7930), .CK(CLK), .QN(n30824) );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n7931), .CK(CLK), .QN(n30825) );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n7932), .CK(CLK), .QN(n30826) );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n7933), .CK(CLK), .QN(n30827) );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n7934), .CK(CLK), .QN(n30828) );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n7935), .CK(CLK), .QN(n30829) );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n7936), .CK(CLK), .QN(n30830) );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n7937), .CK(CLK), .QN(n30831) );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n7938), .CK(CLK), .QN(n30832) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n7939), .CK(CLK), .QN(n30833) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n7940), .CK(CLK), .QN(n30834) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n7941), .CK(CLK), .QN(n30835) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n7942), .CK(CLK), .QN(n30836) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n7943), .CK(CLK), .QN(n30837) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n7944), .CK(CLK), .QN(n30838) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n7945), .CK(CLK), .QN(n30839) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n7946), .CK(CLK), .QN(n30840) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n7947), .CK(CLK), .QN(n30841) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n7948), .CK(CLK), .QN(n30842) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n7949), .CK(CLK), .QN(n30843) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n7950), .CK(CLK), .QN(n30844) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n7951), .CK(CLK), .QN(n30845) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n7952), .CK(CLK), .QN(n30846) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n7953), .CK(CLK), .QN(n30847) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n7954), .CK(CLK), .QN(n30848) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n7955), .CK(CLK), .QN(n30849) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n7956), .CK(CLK), .QN(n30850) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n7957), .CK(CLK), .QN(n30851) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n7958), .CK(CLK), .QN(n30852) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n7959), .CK(CLK), .QN(n30853) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n7960), .CK(CLK), .QN(n30854) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n7961), .CK(CLK), .QN(n30855) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n7962), .CK(CLK), .QN(n30856) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n7963), .CK(CLK), .QN(n30857) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n7964), .CK(CLK), .QN(n30858) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n7965), .CK(CLK), .QN(n30859) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n7966), .CK(CLK), .QN(n30860) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n8099), .CK(CLK), .QN(n30865) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n8100), .CK(CLK), .QN(n30866) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n8101), .CK(CLK), .QN(n30867) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n8102), .CK(CLK), .QN(n30868) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n8103), .CK(CLK), .QN(n30869) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n8104), .CK(CLK), .QN(n30870) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n8105), .CK(CLK), .QN(n30871) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n8106), .CK(CLK), .QN(n30872) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n8107), .CK(CLK), .QN(n30873) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n8108), .CK(CLK), .QN(n30874) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n8109), .CK(CLK), .QN(n30875) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n8110), .CK(CLK), .QN(n30876) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n8111), .CK(CLK), .QN(n30877) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n8112), .CK(CLK), .QN(n30878) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n8113), .CK(CLK), .QN(n30879) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n8114), .CK(CLK), .QN(n30880) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n8115), .CK(CLK), .QN(n30881) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n8116), .CK(CLK), .QN(n30882) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n8117), .CK(CLK), .QN(n30883) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n8118), .CK(CLK), .QN(n30884) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n8119), .CK(CLK), .QN(n30885) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n8120), .CK(CLK), .QN(n30886) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n8121), .CK(CLK), .QN(n30887) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n8122), .CK(CLK), .QN(n30888) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n8123), .CK(CLK), .QN(n30889) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n8124), .CK(CLK), .QN(n30890) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n8125), .CK(CLK), .QN(n30891) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n8126), .CK(CLK), .QN(n30892) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n8127), .CK(CLK), .QN(n30893) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n8128), .CK(CLK), .QN(n30894) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n8129), .CK(CLK), .QN(n30895) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n8130), .CK(CLK), .QN(n30896) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n8131), .CK(CLK), .QN(n30897) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n8132), .CK(CLK), .QN(n30898) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n8133), .CK(CLK), .QN(n30899) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n8134), .CK(CLK), .QN(n30900) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n8135), .CK(CLK), .QN(n30901) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n8136), .CK(CLK), .QN(n30902) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n8137), .CK(CLK), .QN(n30903) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n8138), .CK(CLK), .QN(n30904) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n8139), .CK(CLK), .QN(n30905) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n8140), .CK(CLK), .QN(n30906) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n8141), .CK(CLK), .QN(n30907) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n8142), .CK(CLK), .QN(n30908) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n8143), .CK(CLK), .QN(n30909) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n8144), .CK(CLK), .QN(n30910) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n8145), .CK(CLK), .QN(n30911) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n8146), .CK(CLK), .QN(n30912) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n8147), .CK(CLK), .QN(n30913) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n8148), .CK(CLK), .QN(n30914) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n8149), .CK(CLK), .QN(n30915) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n8150), .CK(CLK), .QN(n30916) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n8151), .CK(CLK), .QN(n30917) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n8152), .CK(CLK), .QN(n30918) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n8153), .CK(CLK), .QN(n30919) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n8154), .CK(CLK), .QN(n30920) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n8155), .CK(CLK), .QN(n30921) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n8156), .CK(CLK), .QN(n30922) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n8157), .CK(CLK), .QN(n30923) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n8158), .CK(CLK), .QN(n30924) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n8159), .CK(CLK), .QN(n30925) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n8160), .CK(CLK), .QN(n30926) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n8161), .CK(CLK), .QN(n30927) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n8162), .CK(CLK), .QN(n30928) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n8163), .CK(CLK), .QN(n30929) );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n8164), .CK(CLK), .QN(n30930) );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n8165), .CK(CLK), .QN(n30931) );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n8166), .CK(CLK), .QN(n30932) );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n8167), .CK(CLK), .QN(n30933) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n8168), .CK(CLK), .QN(n30934) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n8169), .CK(CLK), .QN(n30935) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n8170), .CK(CLK), .QN(n30936) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n8171), .CK(CLK), .QN(n30937) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n8172), .CK(CLK), .QN(n30938) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n8173), .CK(CLK), .QN(n30939) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n8174), .CK(CLK), .QN(n30940) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n8175), .CK(CLK), .QN(n30941) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n8176), .CK(CLK), .QN(n30942) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n8177), .CK(CLK), .QN(n30943) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n8178), .CK(CLK), .QN(n30944) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n8179), .CK(CLK), .QN(n30945) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n8180), .CK(CLK), .QN(n30946) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n8181), .CK(CLK), .QN(n30947) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n8182), .CK(CLK), .QN(n30948) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n8183), .CK(CLK), .QN(n30949) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n8184), .CK(CLK), .QN(n30950) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n8185), .CK(CLK), .QN(n30951) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n8186), .CK(CLK), .QN(n30952) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n8187), .CK(CLK), .QN(n30953) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n8188), .CK(CLK), .QN(n30954) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n8189), .CK(CLK), .QN(n30955) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n8190), .CK(CLK), .QN(n30956) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n8191), .CK(CLK), .QN(n30957) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n8192), .CK(CLK), .QN(n30958) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n8193), .CK(CLK), .QN(n30959) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n8194), .CK(CLK), .QN(n30960) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n8195), .CK(CLK), .QN(n30961) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n8196), .CK(CLK), .QN(n30962) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n8197), .CK(CLK), .QN(n30963) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n8198), .CK(CLK), .QN(n30964) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n8199), .CK(CLK), .QN(n30965) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n8200), .CK(CLK), .QN(n30966) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n8201), .CK(CLK), .QN(n30967) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n8202), .CK(CLK), .QN(n30968) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n8203), .CK(CLK), .QN(n30969) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n8204), .CK(CLK), .QN(n30970) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n8205), .CK(CLK), .QN(n30971) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n8206), .CK(CLK), .QN(n30972) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n8207), .CK(CLK), .QN(n30973) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n8208), .CK(CLK), .QN(n30974) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n8209), .CK(CLK), .QN(n30975) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n8210), .CK(CLK), .QN(n30976) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n8211), .CK(CLK), .QN(n30977) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n8212), .CK(CLK), .QN(n30978) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n8213), .CK(CLK), .QN(n30979) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n8214), .CK(CLK), .QN(n30980) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n8215), .CK(CLK), .QN(n30981) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n8216), .CK(CLK), .QN(n30982) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n8217), .CK(CLK), .QN(n30983) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n8218), .CK(CLK), .QN(n30984) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n8219), .CK(CLK), .QN(n30985) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n8220), .CK(CLK), .QN(n30986) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n8221), .CK(CLK), .QN(n30987) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n8222), .CK(CLK), .QN(n30988) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n8223), .CK(CLK), .QN(n30989) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n8224), .CK(CLK), .QN(n30990) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n8225), .CK(CLK), .QN(n30991) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n8226), .CK(CLK), .QN(n30992) );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n8227), .CK(CLK), .QN(n30993) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n8228), .CK(CLK), .QN(n30994) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n8229), .CK(CLK), .QN(n30995) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n8230), .CK(CLK), .QN(n30996) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n8231), .CK(CLK), .QN(n30997) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n8232), .CK(CLK), .QN(n30998) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n8233), .CK(CLK), .QN(n30999) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n8234), .CK(CLK), .QN(n31000) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n8235), .CK(CLK), .QN(n31001) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n8236), .CK(CLK), .QN(n31002) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n8237), .CK(CLK), .QN(n31003) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n8238), .CK(CLK), .QN(n31004) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n8239), .CK(CLK), .QN(n31005) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n8240), .CK(CLK), .QN(n31006) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n8241), .CK(CLK), .QN(n31007) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n8242), .CK(CLK), .QN(n31008) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n8243), .CK(CLK), .QN(n31009) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n8244), .CK(CLK), .QN(n31010) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n8245), .CK(CLK), .QN(n31011) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n8246), .CK(CLK), .QN(n31012) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n8247), .CK(CLK), .QN(n31013) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n8248), .CK(CLK), .QN(n31014) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n8249), .CK(CLK), .QN(n31015) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n8250), .CK(CLK), .QN(n31016) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n8251), .CK(CLK), .QN(n31017) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n8252), .CK(CLK), .QN(n31018) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n8253), .CK(CLK), .QN(n31019) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n8254), .CK(CLK), .QN(n31020) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n8255), .CK(CLK), .QN(n31021) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n8256), .CK(CLK), .QN(n31022) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n8257), .CK(CLK), .QN(n31023) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n8258), .CK(CLK), .QN(n31024) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n8259), .CK(CLK), .QN(n31025) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n8260), .CK(CLK), .QN(n31026) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n8261), .CK(CLK), .QN(n31027) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n8262), .CK(CLK), .QN(n31028) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n8263), .CK(CLK), .QN(n31029) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n8264), .CK(CLK), .QN(n31030) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n8265), .CK(CLK), .QN(n31031) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n8266), .CK(CLK), .QN(n31032) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n8267), .CK(CLK), .QN(n31033) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n8268), .CK(CLK), .QN(n31034) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n8269), .CK(CLK), .QN(n31035) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n8270), .CK(CLK), .QN(n31036) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n8271), .CK(CLK), .QN(n31037) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n8272), .CK(CLK), .QN(n31038) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n8273), .CK(CLK), .QN(n31039) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n8274), .CK(CLK), .QN(n31040) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n8275), .CK(CLK), .QN(n31041) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n8276), .CK(CLK), .QN(n31042) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n8277), .CK(CLK), .QN(n31043) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n8278), .CK(CLK), .QN(n31044) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n8279), .CK(CLK), .QN(n31045) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n8280), .CK(CLK), .QN(n31046) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n8281), .CK(CLK), .QN(n31047) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n8282), .CK(CLK), .QN(n31048) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n8283), .CK(CLK), .QN(n31049) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n8284), .CK(CLK), .QN(n31050) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n8285), .CK(CLK), .QN(n31051) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n8286), .CK(CLK), .QN(n31052) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n8287), .CK(CLK), .QN(n31053) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n8288), .CK(CLK), .QN(n31054) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n8289), .CK(CLK), .QN(n31055) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n8290), .CK(CLK), .QN(n31056) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n8419), .CK(CLK), .QN(n31175) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n8420), .CK(CLK), .QN(n31176) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n8421), .CK(CLK), .QN(n31177) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n8422), .CK(CLK), .QN(n31178) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n8423), .CK(CLK), .QN(n31179) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n8424), .CK(CLK), .QN(n31180) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n8425), .CK(CLK), .QN(n31181) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n8426), .CK(CLK), .QN(n31182) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n8427), .CK(CLK), .QN(n31183) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n8428), .CK(CLK), .QN(n31184) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n8429), .CK(CLK), .QN(n31185) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n8430), .CK(CLK), .QN(n31186) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n8431), .CK(CLK), .QN(n31187) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n8432), .CK(CLK), .QN(n31188) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n8433), .CK(CLK), .QN(n31189) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n8434), .CK(CLK), .QN(n31190) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n8435), .CK(CLK), .QN(n31191) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n8436), .CK(CLK), .QN(n31192) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n8437), .CK(CLK), .QN(n31193) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n8438), .CK(CLK), .QN(n31194) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n8439), .CK(CLK), .QN(n31195) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n8440), .CK(CLK), .QN(n31196) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n8441), .CK(CLK), .QN(n31197) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n8442), .CK(CLK), .QN(n31198) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n8443), .CK(CLK), .QN(n31199) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n8444), .CK(CLK), .QN(n31200) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n8445), .CK(CLK), .QN(n31201) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n8446), .CK(CLK), .QN(n31202) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n8447), .CK(CLK), .QN(n31203) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n8448), .CK(CLK), .QN(n31204) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n8449), .CK(CLK), .QN(n31205) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n8450), .CK(CLK), .QN(n31206) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n8451), .CK(CLK), .QN(n31207) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n8452), .CK(CLK), .QN(n31208) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n8453), .CK(CLK), .QN(n31209) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n8454), .CK(CLK), .QN(n31210) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n8455), .CK(CLK), .QN(n31211) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n8456), .CK(CLK), .QN(n31212) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n8457), .CK(CLK), .QN(n31213) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n8458), .CK(CLK), .QN(n31214) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n8459), .CK(CLK), .QN(n31215) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n8460), .CK(CLK), .QN(n31216) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n8461), .CK(CLK), .QN(n31217) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n8462), .CK(CLK), .QN(n31218) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n8463), .CK(CLK), .QN(n31219) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n8464), .CK(CLK), .QN(n31220) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n8465), .CK(CLK), .QN(n31221) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n8466), .CK(CLK), .QN(n31222) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n8467), .CK(CLK), .QN(n31223) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n8468), .CK(CLK), .QN(n31224) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n8469), .CK(CLK), .QN(n31225) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n8470), .CK(CLK), .QN(n31226) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n8471), .CK(CLK), .QN(n31227) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n8472), .CK(CLK), .QN(n31228) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n8473), .CK(CLK), .QN(n31229) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n8474), .CK(CLK), .QN(n31230) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n8475), .CK(CLK), .QN(n31231) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n8476), .CK(CLK), .QN(n31232) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n8477), .CK(CLK), .QN(n31233) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n8478), .CK(CLK), .QN(n31234) );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n8483), .CK(CLK), .QN(n31239) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n8484), .CK(CLK), .QN(n31240) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n8485), .CK(CLK), .QN(n31241) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n8486), .CK(CLK), .QN(n31242) );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n8487), .CK(CLK), .QN(n31243) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n8488), .CK(CLK), .QN(n31244) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n8489), .CK(CLK), .QN(n31245) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n8490), .CK(CLK), .QN(n31246) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n8491), .CK(CLK), .QN(n31247) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n8492), .CK(CLK), .QN(n31248) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n8493), .CK(CLK), .QN(n31249) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n8494), .CK(CLK), .QN(n31250) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n8495), .CK(CLK), .QN(n31251) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n8496), .CK(CLK), .QN(n31252) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n8497), .CK(CLK), .QN(n31253) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n8498), .CK(CLK), .QN(n31254) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n8499), .CK(CLK), .QN(n31255) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n8500), .CK(CLK), .QN(n31256) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n8501), .CK(CLK), .QN(n31257) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n8502), .CK(CLK), .QN(n31258) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n8503), .CK(CLK), .QN(n31259) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n8504), .CK(CLK), .QN(n31260) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n8505), .CK(CLK), .QN(n31261) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n8506), .CK(CLK), .QN(n31262) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n8507), .CK(CLK), .QN(n31263) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n8508), .CK(CLK), .QN(n31264) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n8509), .CK(CLK), .QN(n31265) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n8510), .CK(CLK), .QN(n31266) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n8511), .CK(CLK), .QN(n31267) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n8512), .CK(CLK), .QN(n31268) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n8513), .CK(CLK), .QN(n31269) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n8514), .CK(CLK), .QN(n31270) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n8515), .CK(CLK), .QN(n31271) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n8516), .CK(CLK), .QN(n31272) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n8517), .CK(CLK), .QN(n31273) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n8518), .CK(CLK), .QN(n31274) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n8519), .CK(CLK), .QN(n31275) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n8520), .CK(CLK), .QN(n31276) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n8521), .CK(CLK), .QN(n31277) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n8522), .CK(CLK), .QN(n31278) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n8523), .CK(CLK), .QN(n31279) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n8524), .CK(CLK), .QN(n31280) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n8525), .CK(CLK), .QN(n31281) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n8526), .CK(CLK), .QN(n31282) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n8527), .CK(CLK), .QN(n31283) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n8528), .CK(CLK), .QN(n31284) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n8529), .CK(CLK), .QN(n31285) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n8530), .CK(CLK), .QN(n31286) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n8531), .CK(CLK), .QN(n31287) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n8532), .CK(CLK), .QN(n31288) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n8533), .CK(CLK), .QN(n31289) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n8534), .CK(CLK), .QN(n31290) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n8535), .CK(CLK), .QN(n31291) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n8536), .CK(CLK), .QN(n31292) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n8537), .CK(CLK), .QN(n31293) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n8538), .CK(CLK), .QN(n31294) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n8539), .CK(CLK), .QN(n31295) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n8540), .CK(CLK), .QN(n31296) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n8541), .CK(CLK), .QN(n31297) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n8542), .CK(CLK), .QN(n31298) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n8547), .CK(CLK), .QN(n31303) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n8548), .CK(CLK), .QN(n31304) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n8549), .CK(CLK), .QN(n31305) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n8550), .CK(CLK), .QN(n31306) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n8551), .CK(CLK), .QN(n31307) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n8552), .CK(CLK), .QN(n31308) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n8553), .CK(CLK), .QN(n31309) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n8554), .CK(CLK), .QN(n31310) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n8555), .CK(CLK), .QN(n31311) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n8556), .CK(CLK), .QN(n31312) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n8557), .CK(CLK), .QN(n31313) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n8558), .CK(CLK), .QN(n31314) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n8559), .CK(CLK), .QN(n31315) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n8560), .CK(CLK), .QN(n31316) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n8561), .CK(CLK), .QN(n31317) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n8562), .CK(CLK), .QN(n31318) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n8563), .CK(CLK), .QN(n31319) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n8564), .CK(CLK), .QN(n31320) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n8565), .CK(CLK), .QN(n31321) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n8566), .CK(CLK), .QN(n31322) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n8567), .CK(CLK), .QN(n31323) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n8568), .CK(CLK), .QN(n31324) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n8569), .CK(CLK), .QN(n31325) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n8570), .CK(CLK), .QN(n31326) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n8571), .CK(CLK), .QN(n31327) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n8572), .CK(CLK), .QN(n31328) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n8573), .CK(CLK), .QN(n31329) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n8574), .CK(CLK), .QN(n31330) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n8575), .CK(CLK), .QN(n31331) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n8576), .CK(CLK), .QN(n31332) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n8577), .CK(CLK), .QN(n31333) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n8578), .CK(CLK), .QN(n31334) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n8579), .CK(CLK), .QN(n31335) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n8580), .CK(CLK), .QN(n31336) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n8581), .CK(CLK), .QN(n31337) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n8582), .CK(CLK), .QN(n31338) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n8583), .CK(CLK), .QN(n31339) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n8584), .CK(CLK), .QN(n31340) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n8585), .CK(CLK), .QN(n31341) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n8586), .CK(CLK), .QN(n31342) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n8587), .CK(CLK), .QN(n31343) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n8588), .CK(CLK), .QN(n31344) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n8589), .CK(CLK), .QN(n31345) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n8590), .CK(CLK), .QN(n31346) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n8591), .CK(CLK), .QN(n31347) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n8592), .CK(CLK), .QN(n31348) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n8593), .CK(CLK), .QN(n31349) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n8594), .CK(CLK), .QN(n31350) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n8595), .CK(CLK), .QN(n31351) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n8596), .CK(CLK), .QN(n31352) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n8597), .CK(CLK), .QN(n31353) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n8598), .CK(CLK), .QN(n31354) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n8599), .CK(CLK), .QN(n31355) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n8600), .CK(CLK), .QN(n31356) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n8601), .CK(CLK), .QN(n31357) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n8602), .CK(CLK), .QN(n31358) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n8603), .CK(CLK), .QN(n31359) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n8604), .CK(CLK), .QN(n31360) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n8605), .CK(CLK), .QN(n31361) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n8606), .CK(CLK), .QN(n31362) );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n8739), .CK(CLK), .QN(n31367) );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n8740), .CK(CLK), .QN(n31368) );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n8741), .CK(CLK), .QN(n31369) );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n8742), .CK(CLK), .QN(n31370) );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n8743), .CK(CLK), .QN(n31371) );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n8744), .CK(CLK), .QN(n31372) );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n8745), .CK(CLK), .QN(n31373) );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n8746), .CK(CLK), .QN(n31374) );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n8747), .CK(CLK), .QN(n31375) );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n8748), .CK(CLK), .QN(n31376) );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n8749), .CK(CLK), .QN(n31377) );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n8750), .CK(CLK), .QN(n31378) );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n8751), .CK(CLK), .QN(n31379) );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n8752), .CK(CLK), .QN(n31380) );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n8753), .CK(CLK), .QN(n31381) );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n8754), .CK(CLK), .QN(n31382) );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n8755), .CK(CLK), .QN(n31383) );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n8756), .CK(CLK), .QN(n31384) );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n8757), .CK(CLK), .QN(n31385) );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n8758), .CK(CLK), .QN(n31386) );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n8759), .CK(CLK), .QN(n31387) );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n8760), .CK(CLK), .QN(n31388) );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n8761), .CK(CLK), .QN(n31389) );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n8762), .CK(CLK), .QN(n31390) );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n8763), .CK(CLK), .QN(n31391) );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n8764), .CK(CLK), .QN(n31392) );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n8765), .CK(CLK), .QN(n31393) );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n8766), .CK(CLK), .QN(n31394) );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n8767), .CK(CLK), .QN(n31395) );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n8768), .CK(CLK), .QN(n31396) );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n8769), .CK(CLK), .QN(n31397) );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n8770), .CK(CLK), .QN(n31398) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n8771), .CK(CLK), .QN(n31399) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n8772), .CK(CLK), .QN(n31400) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n8773), .CK(CLK), .QN(n31401) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n8774), .CK(CLK), .QN(n31402) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n8775), .CK(CLK), .QN(n31403) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n8776), .CK(CLK), .QN(n31404) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n8777), .CK(CLK), .QN(n31405) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n8778), .CK(CLK), .QN(n31406) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n8779), .CK(CLK), .QN(n31407) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n8780), .CK(CLK), .QN(n31408) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n8781), .CK(CLK), .QN(n31409) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n8782), .CK(CLK), .QN(n31410) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n8783), .CK(CLK), .QN(n31411) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n8784), .CK(CLK), .QN(n31412) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n8785), .CK(CLK), .QN(n31413) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n8786), .CK(CLK), .QN(n31414) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n8787), .CK(CLK), .QN(n31415) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n8788), .CK(CLK), .QN(n31416) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n8789), .CK(CLK), .QN(n31417) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n8790), .CK(CLK), .QN(n31418) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n8791), .CK(CLK), .QN(n31419) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n8792), .CK(CLK), .QN(n31420) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n8793), .CK(CLK), .QN(n31421) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n8794), .CK(CLK), .QN(n31422) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n8795), .CK(CLK), .QN(n31423) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n8796), .CK(CLK), .QN(n31424) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n8797), .CK(CLK), .QN(n31425) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n8798), .CK(CLK), .QN(n31426) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n8799), .CK(CLK), .QN(n31427) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n8800), .CK(CLK), .QN(n31428) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n8801), .CK(CLK), .QN(n31429) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n8802), .CK(CLK), .QN(n31430) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n8803), .CK(CLK), .QN(n31431) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n8804), .CK(CLK), .QN(n31432) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n8805), .CK(CLK), .QN(n31433) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n8806), .CK(CLK), .QN(n31434) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n8807), .CK(CLK), .QN(n31435) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n8808), .CK(CLK), .QN(n31436) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n8809), .CK(CLK), .QN(n31437) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n8810), .CK(CLK), .QN(n31438) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n8811), .CK(CLK), .QN(n31439) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n8812), .CK(CLK), .QN(n31440) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n8813), .CK(CLK), .QN(n31441) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n8814), .CK(CLK), .QN(n31442) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n8815), .CK(CLK), .QN(n31443) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n8816), .CK(CLK), .QN(n31444) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n8817), .CK(CLK), .QN(n31445) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n8818), .CK(CLK), .QN(n31446) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n8819), .CK(CLK), .QN(n31447) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n8820), .CK(CLK), .QN(n31448) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n8821), .CK(CLK), .QN(n31449) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n8822), .CK(CLK), .QN(n31450) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n8823), .CK(CLK), .QN(n31451) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n8824), .CK(CLK), .QN(n31452) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n8825), .CK(CLK), .QN(n31453) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n8826), .CK(CLK), .QN(n31454) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n8827), .CK(CLK), .QN(n31455) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n8828), .CK(CLK), .QN(n31456) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n8829), .CK(CLK), .QN(n31457) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n8830), .CK(CLK), .QN(n31458) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n8831), .CK(CLK), .QN(n31459) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n8832), .CK(CLK), .QN(n31460) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n8833), .CK(CLK), .QN(n31461) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n8834), .CK(CLK), .QN(n31462) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n8835), .CK(CLK), .QN(n31463) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n8836), .CK(CLK), .QN(n31464) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n8837), .CK(CLK), .QN(n31465) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n8838), .CK(CLK), .QN(n31466) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n8839), .CK(CLK), .QN(n31467) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n8840), .CK(CLK), .QN(n31468) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n8841), .CK(CLK), .QN(n31469) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n8842), .CK(CLK), .QN(n31470) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n8843), .CK(CLK), .QN(n31471) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n8844), .CK(CLK), .QN(n31472) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n8845), .CK(CLK), .QN(n31473) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n8846), .CK(CLK), .QN(n31474) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n8847), .CK(CLK), .QN(n31475) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n8848), .CK(CLK), .QN(n31476) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n8849), .CK(CLK), .QN(n31477) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n8850), .CK(CLK), .QN(n31478) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n8851), .CK(CLK), .QN(n31479) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n8852), .CK(CLK), .QN(n31480) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n8853), .CK(CLK), .QN(n31481) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n8854), .CK(CLK), .QN(n31482) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n8855), .CK(CLK), .QN(n31483) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n8856), .CK(CLK), .QN(n31484) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n8857), .CK(CLK), .QN(n31485) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n8858), .CK(CLK), .QN(n31486) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n8859), .CK(CLK), .QN(n31487) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n8860), .CK(CLK), .QN(n31488) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n8861), .CK(CLK), .QN(n31489) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n8862), .CK(CLK), .QN(n31490) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n8863), .CK(CLK), .QN(n31491) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n8864), .CK(CLK), .QN(n31492) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n8865), .CK(CLK), .QN(n31493) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n8866), .CK(CLK), .QN(n31494) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n8867), .CK(CLK), .QN(n31495) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n8868), .CK(CLK), .QN(n31496) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n8869), .CK(CLK), .QN(n31497) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n8870), .CK(CLK), .QN(n31498) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n8871), .CK(CLK), .QN(n31499) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n8872), .CK(CLK), .QN(n31500) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n8873), .CK(CLK), .QN(n31501) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n8874), .CK(CLK), .QN(n31502) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n8875), .CK(CLK), .QN(n31503) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n8876), .CK(CLK), .QN(n31504) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n8877), .CK(CLK), .QN(n31505) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n8878), .CK(CLK), .QN(n31506) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n8879), .CK(CLK), .QN(n31507) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n8880), .CK(CLK), .QN(n31508) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n8881), .CK(CLK), .QN(n31509) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n8882), .CK(CLK), .QN(n31510) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n8883), .CK(CLK), .QN(n31511) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n8884), .CK(CLK), .QN(n31512) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n8885), .CK(CLK), .QN(n31513) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n8886), .CK(CLK), .QN(n31514) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n8887), .CK(CLK), .QN(n31515) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n8888), .CK(CLK), .QN(n31516) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n8889), .CK(CLK), .QN(n31517) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n8890), .CK(CLK), .QN(n31518) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n8891), .CK(CLK), .QN(n31519) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n8892), .CK(CLK), .QN(n31520) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n8893), .CK(CLK), .QN(n31521) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n8894), .CK(CLK), .QN(n31522) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n8895), .CK(CLK), .QN(n31523) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n8896), .CK(CLK), .QN(n31524) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n8897), .CK(CLK), .QN(n31525) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n8898), .CK(CLK), .QN(n31526) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n8899), .CK(CLK), .QN(n31527) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n8900), .CK(CLK), .QN(n31528) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n8901), .CK(CLK), .QN(n31529) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n8902), .CK(CLK), .QN(n31530) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n8903), .CK(CLK), .QN(n31531) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n8904), .CK(CLK), .QN(n31532) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n8905), .CK(CLK), .QN(n31533) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n8906), .CK(CLK), .QN(n31534) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n8907), .CK(CLK), .QN(n31535) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n8908), .CK(CLK), .QN(n31536) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n8909), .CK(CLK), .QN(n31537) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n8910), .CK(CLK), .QN(n31538) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n8911), .CK(CLK), .QN(n31539) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n8912), .CK(CLK), .QN(n31540) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n8913), .CK(CLK), .QN(n31541) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n8914), .CK(CLK), .QN(n31542) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n8915), .CK(CLK), .QN(n31543) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n8916), .CK(CLK), .QN(n31544) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n8917), .CK(CLK), .QN(n31545) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n8918), .CK(CLK), .QN(n31546) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n8919), .CK(CLK), .QN(n31547) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n8920), .CK(CLK), .QN(n31548) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n8921), .CK(CLK), .QN(n31549) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n8922), .CK(CLK), .QN(n31550) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n8923), .CK(CLK), .QN(n31551) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n8924), .CK(CLK), .QN(n31552) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n8925), .CK(CLK), .QN(n31553) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n8926), .CK(CLK), .QN(n31554) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n8927), .CK(CLK), .QN(n31555) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n8928), .CK(CLK), .QN(n31556) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n8929), .CK(CLK), .QN(n31557) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n8930), .CK(CLK), .QN(n31558) );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n9059), .CK(CLK), .QN(n31559) );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n9060), .CK(CLK), .QN(n31560) );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n9061), .CK(CLK), .QN(n31561) );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n9062), .CK(CLK), .QN(n31562) );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n9063), .CK(CLK), .QN(n31563) );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n9064), .CK(CLK), .QN(n31564) );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n9065), .CK(CLK), .QN(n31565) );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n9066), .CK(CLK), .QN(n31566) );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n9067), .CK(CLK), .QN(n31567) );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n9068), .CK(CLK), .QN(n31568) );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n9069), .CK(CLK), .QN(n31569) );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n9070), .CK(CLK), .QN(n31570) );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n9071), .CK(CLK), .QN(n31571) );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n9072), .CK(CLK), .QN(n31572) );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n9073), .CK(CLK), .QN(n31573) );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n9074), .CK(CLK), .QN(n31574) );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n9075), .CK(CLK), .QN(n31575) );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n9076), .CK(CLK), .QN(n31576) );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n9077), .CK(CLK), .QN(n31577) );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n9078), .CK(CLK), .QN(n31578) );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n9079), .CK(CLK), .QN(n31579) );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n9080), .CK(CLK), .QN(n31580) );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n9081), .CK(CLK), .QN(n31581) );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n9082), .CK(CLK), .QN(n31582) );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n9083), .CK(CLK), .QN(n31583) );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n9084), .CK(CLK), .QN(n31584) );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n9085), .CK(CLK), .QN(n31585) );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n9086), .CK(CLK), .QN(n31586) );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n9087), .CK(CLK), .QN(n31587) );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n9088), .CK(CLK), .QN(n31588) );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n9089), .CK(CLK), .QN(n31589) );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n9090), .CK(CLK), .QN(n31590) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n9091), .CK(CLK), .QN(n31591) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n9092), .CK(CLK), .QN(n31592) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n9093), .CK(CLK), .QN(n31593) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n9094), .CK(CLK), .QN(n31594) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n9095), .CK(CLK), .QN(n31595) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n9096), .CK(CLK), .QN(n31596) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n9097), .CK(CLK), .QN(n31597) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n9098), .CK(CLK), .QN(n31598) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n9099), .CK(CLK), .QN(n31599) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n9100), .CK(CLK), .QN(n31600) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n9101), .CK(CLK), .QN(n31601) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n9102), .CK(CLK), .QN(n31602) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n9103), .CK(CLK), .QN(n31603) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n9104), .CK(CLK), .QN(n31604) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n9105), .CK(CLK), .QN(n31605) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n9106), .CK(CLK), .QN(n31606) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n9107), .CK(CLK), .QN(n31607) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n9108), .CK(CLK), .QN(n31608) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n9109), .CK(CLK), .QN(n31609) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n9110), .CK(CLK), .QN(n31610) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n9111), .CK(CLK), .QN(n31611) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n9112), .CK(CLK), .QN(n31612) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n9113), .CK(CLK), .QN(n31613) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n9114), .CK(CLK), .QN(n31614) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n9115), .CK(CLK), .QN(n31615) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n9116), .CK(CLK), .QN(n31616) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n9117), .CK(CLK), .QN(n31617) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n9118), .CK(CLK), .QN(n31618) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n9119), .CK(CLK), .QN(n31619) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n9120), .CK(CLK), .QN(n31620) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n9121), .CK(CLK), .QN(n31621) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n9122), .CK(CLK), .QN(n31622) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n9123), .CK(CLK), .QN(n31623) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n9124), .CK(CLK), .QN(n31624) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n9125), .CK(CLK), .QN(n31625) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n9126), .CK(CLK), .QN(n31626) );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n9127), .CK(CLK), .QN(n31627) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n9128), .CK(CLK), .QN(n31628) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n9129), .CK(CLK), .QN(n31629) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n9130), .CK(CLK), .QN(n31630) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n9131), .CK(CLK), .QN(n31631) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n9132), .CK(CLK), .QN(n31632) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n9133), .CK(CLK), .QN(n31633) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n9134), .CK(CLK), .QN(n31634) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n9135), .CK(CLK), .QN(n31635) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n9136), .CK(CLK), .QN(n31636) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n9137), .CK(CLK), .QN(n31637) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n9138), .CK(CLK), .QN(n31638) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n9139), .CK(CLK), .QN(n31639) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n9140), .CK(CLK), .QN(n31640) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n9141), .CK(CLK), .QN(n31641) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n9142), .CK(CLK), .QN(n31642) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n9143), .CK(CLK), .QN(n31643) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n9144), .CK(CLK), .QN(n31644) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n9145), .CK(CLK), .QN(n31645) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n9146), .CK(CLK), .QN(n31646) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n9147), .CK(CLK), .QN(n31647) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n9148), .CK(CLK), .QN(n31648) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n9149), .CK(CLK), .QN(n31649) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n9150), .CK(CLK), .QN(n31650) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n9151), .CK(CLK), .QN(n31651) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n9152), .CK(CLK), .QN(n31652) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n9153), .CK(CLK), .QN(n31653) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n9154), .CK(CLK), .QN(n31654) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n9155), .CK(CLK), .QN(n31655) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n9156), .CK(CLK), .QN(n31656) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n9157), .CK(CLK), .QN(n31657) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n9158), .CK(CLK), .QN(n31658) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n9159), .CK(CLK), .QN(n31659) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n9160), .CK(CLK), .QN(n31660) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n9161), .CK(CLK), .QN(n31661) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n9162), .CK(CLK), .QN(n31662) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n9163), .CK(CLK), .QN(n31663) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n9164), .CK(CLK), .QN(n31664) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n9165), .CK(CLK), .QN(n31665) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n9166), .CK(CLK), .QN(n31666) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n9167), .CK(CLK), .QN(n31667) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n9168), .CK(CLK), .QN(n31668) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n9169), .CK(CLK), .QN(n31669) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n9170), .CK(CLK), .QN(n31670) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n9171), .CK(CLK), .QN(n31671) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n9172), .CK(CLK), .QN(n31672) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n9173), .CK(CLK), .QN(n31673) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n9174), .CK(CLK), .QN(n31674) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n9175), .CK(CLK), .QN(n31675) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n9176), .CK(CLK), .QN(n31676) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n9177), .CK(CLK), .QN(n31677) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n9178), .CK(CLK), .QN(n31678) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n9179), .CK(CLK), .QN(n31679) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n9180), .CK(CLK), .QN(n31680) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n9181), .CK(CLK), .QN(n31681) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n9182), .CK(CLK), .QN(n31682) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n9183), .CK(CLK), .QN(n31683) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n9184), .CK(CLK), .QN(n31684) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n9185), .CK(CLK), .QN(n31685) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n9186), .CK(CLK), .QN(n31686) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n9187), .CK(CLK), .QN(n31687) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n9188), .CK(CLK), .QN(n31688) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n9189), .CK(CLK), .QN(n31689) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n9190), .CK(CLK), .QN(n31690) );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n9191), .CK(CLK), .QN(n31691) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n9192), .CK(CLK), .QN(n31692) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n9193), .CK(CLK), .QN(n31693) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n9194), .CK(CLK), .QN(n31694) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n9195), .CK(CLK), .QN(n31695) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n9196), .CK(CLK), .QN(n31696) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n9197), .CK(CLK), .QN(n31697) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n9198), .CK(CLK), .QN(n31698) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n9199), .CK(CLK), .QN(n31699) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n9200), .CK(CLK), .QN(n31700) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n9201), .CK(CLK), .QN(n31701) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n9202), .CK(CLK), .QN(n31702) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n9203), .CK(CLK), .QN(n31703) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n9204), .CK(CLK), .QN(n31704) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n9205), .CK(CLK), .QN(n31705) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n9206), .CK(CLK), .QN(n31706) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n9207), .CK(CLK), .QN(n31707) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n9208), .CK(CLK), .QN(n31708) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n9209), .CK(CLK), .QN(n31709) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n9210), .CK(CLK), .QN(n31710) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n9211), .CK(CLK), .QN(n31711) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n9212), .CK(CLK), .QN(n31712) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n9213), .CK(CLK), .QN(n31713) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n9214), .CK(CLK), .QN(n31714) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n9215), .CK(CLK), .QN(n31715) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n9216), .CK(CLK), .QN(n31716) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n9217), .CK(CLK), .QN(n31717) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n9218), .CK(CLK), .QN(n31718) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n9219), .CK(CLK), .QN(n31719) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n9220), .CK(CLK), .QN(n31720) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n9221), .CK(CLK), .QN(n31721) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n9222), .CK(CLK), .QN(n31722) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n9223), .CK(CLK), .QN(n31723) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n9224), .CK(CLK), .QN(n31724) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n9225), .CK(CLK), .QN(n31725) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n9226), .CK(CLK), .QN(n31726) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n9227), .CK(CLK), .QN(n31727) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n9228), .CK(CLK), .QN(n31728) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n9229), .CK(CLK), .QN(n31729) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n9230), .CK(CLK), .QN(n31730) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n9231), .CK(CLK), .QN(n31731) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n9232), .CK(CLK), .QN(n31732) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n9233), .CK(CLK), .QN(n31733) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n9234), .CK(CLK), .QN(n31734) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n9235), .CK(CLK), .QN(n31735) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n9236), .CK(CLK), .QN(n31736) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n9237), .CK(CLK), .QN(n31737) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n9238), .CK(CLK), .QN(n31738) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n9239), .CK(CLK), .QN(n31739) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n9240), .CK(CLK), .QN(n31740) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n9241), .CK(CLK), .QN(n31741) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n9242), .CK(CLK), .QN(n31742) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n9243), .CK(CLK), .QN(n31743) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n9244), .CK(CLK), .QN(n31744) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n9245), .CK(CLK), .QN(n31745) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n9246), .CK(CLK), .QN(n31746) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n9247), .CK(CLK), .QN(n31747) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n9248), .CK(CLK), .QN(n31748) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n9249), .CK(CLK), .QN(n31749) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n9250), .CK(CLK), .QN(n31750) );
  DFF_X1 \REGISTERS_reg[32][63]  ( .D(n9379), .CK(CLK), .QN(n31751) );
  DFF_X1 \REGISTERS_reg[32][62]  ( .D(n9380), .CK(CLK), .QN(n31752) );
  DFF_X1 \REGISTERS_reg[32][61]  ( .D(n9381), .CK(CLK), .QN(n31753) );
  DFF_X1 \REGISTERS_reg[32][60]  ( .D(n9382), .CK(CLK), .QN(n31754) );
  DFF_X1 \REGISTERS_reg[32][59]  ( .D(n9383), .CK(CLK), .QN(n31755) );
  DFF_X1 \REGISTERS_reg[32][58]  ( .D(n9384), .CK(CLK), .QN(n31756) );
  DFF_X1 \REGISTERS_reg[32][57]  ( .D(n9385), .CK(CLK), .QN(n31757) );
  DFF_X1 \REGISTERS_reg[32][56]  ( .D(n9386), .CK(CLK), .QN(n31758) );
  DFF_X1 \REGISTERS_reg[32][55]  ( .D(n9387), .CK(CLK), .QN(n31759) );
  DFF_X1 \REGISTERS_reg[32][54]  ( .D(n9388), .CK(CLK), .QN(n31760) );
  DFF_X1 \REGISTERS_reg[32][53]  ( .D(n9389), .CK(CLK), .QN(n31761) );
  DFF_X1 \REGISTERS_reg[32][52]  ( .D(n9390), .CK(CLK), .QN(n31762) );
  DFF_X1 \REGISTERS_reg[32][51]  ( .D(n9391), .CK(CLK), .QN(n31763) );
  DFF_X1 \REGISTERS_reg[32][50]  ( .D(n9392), .CK(CLK), .QN(n31764) );
  DFF_X1 \REGISTERS_reg[32][49]  ( .D(n9393), .CK(CLK), .QN(n31765) );
  DFF_X1 \REGISTERS_reg[32][48]  ( .D(n9394), .CK(CLK), .QN(n31766) );
  DFF_X1 \REGISTERS_reg[32][47]  ( .D(n9395), .CK(CLK), .QN(n31767) );
  DFF_X1 \REGISTERS_reg[32][46]  ( .D(n9396), .CK(CLK), .QN(n31768) );
  DFF_X1 \REGISTERS_reg[32][45]  ( .D(n9397), .CK(CLK), .QN(n31769) );
  DFF_X1 \REGISTERS_reg[32][44]  ( .D(n9398), .CK(CLK), .QN(n31770) );
  DFF_X1 \REGISTERS_reg[32][43]  ( .D(n9399), .CK(CLK), .QN(n31771) );
  DFF_X1 \REGISTERS_reg[32][42]  ( .D(n9400), .CK(CLK), .QN(n31772) );
  DFF_X1 \REGISTERS_reg[32][41]  ( .D(n9401), .CK(CLK), .QN(n31773) );
  DFF_X1 \REGISTERS_reg[32][40]  ( .D(n9402), .CK(CLK), .QN(n31774) );
  DFF_X1 \REGISTERS_reg[32][39]  ( .D(n9403), .CK(CLK), .QN(n31775) );
  DFF_X1 \REGISTERS_reg[32][38]  ( .D(n9404), .CK(CLK), .QN(n31776) );
  DFF_X1 \REGISTERS_reg[32][37]  ( .D(n9405), .CK(CLK), .QN(n31777) );
  DFF_X1 \REGISTERS_reg[32][36]  ( .D(n9406), .CK(CLK), .QN(n31778) );
  DFF_X1 \REGISTERS_reg[32][35]  ( .D(n9407), .CK(CLK), .QN(n31779) );
  DFF_X1 \REGISTERS_reg[32][34]  ( .D(n9408), .CK(CLK), .QN(n31780) );
  DFF_X1 \REGISTERS_reg[32][33]  ( .D(n9409), .CK(CLK), .QN(n31781) );
  DFF_X1 \REGISTERS_reg[32][32]  ( .D(n9410), .CK(CLK), .QN(n31782) );
  DFF_X1 \REGISTERS_reg[32][31]  ( .D(n9411), .CK(CLK), .QN(n31783) );
  DFF_X1 \REGISTERS_reg[32][30]  ( .D(n9412), .CK(CLK), .QN(n31784) );
  DFF_X1 \REGISTERS_reg[32][29]  ( .D(n9413), .CK(CLK), .QN(n31785) );
  DFF_X1 \REGISTERS_reg[32][28]  ( .D(n9414), .CK(CLK), .QN(n31786) );
  DFF_X1 \REGISTERS_reg[32][27]  ( .D(n9415), .CK(CLK), .QN(n31787) );
  DFF_X1 \REGISTERS_reg[32][26]  ( .D(n9416), .CK(CLK), .QN(n31788) );
  DFF_X1 \REGISTERS_reg[32][25]  ( .D(n9417), .CK(CLK), .QN(n31789) );
  DFF_X1 \REGISTERS_reg[32][24]  ( .D(n9418), .CK(CLK), .QN(n31790) );
  DFF_X1 \REGISTERS_reg[32][23]  ( .D(n9419), .CK(CLK), .QN(n31791) );
  DFF_X1 \REGISTERS_reg[32][22]  ( .D(n9420), .CK(CLK), .QN(n31792) );
  DFF_X1 \REGISTERS_reg[32][21]  ( .D(n9421), .CK(CLK), .QN(n31793) );
  DFF_X1 \REGISTERS_reg[32][20]  ( .D(n9422), .CK(CLK), .QN(n31794) );
  DFF_X1 \REGISTERS_reg[32][19]  ( .D(n9423), .CK(CLK), .QN(n31795) );
  DFF_X1 \REGISTERS_reg[32][18]  ( .D(n9424), .CK(CLK), .QN(n31796) );
  DFF_X1 \REGISTERS_reg[32][17]  ( .D(n9425), .CK(CLK), .QN(n31797) );
  DFF_X1 \REGISTERS_reg[32][16]  ( .D(n9426), .CK(CLK), .QN(n31798) );
  DFF_X1 \REGISTERS_reg[32][15]  ( .D(n9427), .CK(CLK), .QN(n31799) );
  DFF_X1 \REGISTERS_reg[32][14]  ( .D(n9428), .CK(CLK), .QN(n31800) );
  DFF_X1 \REGISTERS_reg[32][13]  ( .D(n9429), .CK(CLK), .QN(n31801) );
  DFF_X1 \REGISTERS_reg[32][12]  ( .D(n9430), .CK(CLK), .QN(n31802) );
  DFF_X1 \REGISTERS_reg[32][11]  ( .D(n9431), .CK(CLK), .QN(n31803) );
  DFF_X1 \REGISTERS_reg[32][10]  ( .D(n9432), .CK(CLK), .QN(n31804) );
  DFF_X1 \REGISTERS_reg[32][9]  ( .D(n9433), .CK(CLK), .QN(n31805) );
  DFF_X1 \REGISTERS_reg[32][8]  ( .D(n9434), .CK(CLK), .QN(n31806) );
  DFF_X1 \REGISTERS_reg[32][7]  ( .D(n9435), .CK(CLK), .QN(n31807) );
  DFF_X1 \REGISTERS_reg[32][6]  ( .D(n9436), .CK(CLK), .QN(n31808) );
  DFF_X1 \REGISTERS_reg[32][5]  ( .D(n9437), .CK(CLK), .QN(n31809) );
  DFF_X1 \REGISTERS_reg[32][4]  ( .D(n9438), .CK(CLK), .QN(n31810) );
  DFF_X1 \REGISTERS_reg[33][63]  ( .D(n9443), .CK(CLK), .QN(n31811) );
  DFF_X1 \REGISTERS_reg[33][62]  ( .D(n9444), .CK(CLK), .QN(n31812) );
  DFF_X1 \REGISTERS_reg[33][61]  ( .D(n9445), .CK(CLK), .QN(n31813) );
  DFF_X1 \REGISTERS_reg[33][60]  ( .D(n9446), .CK(CLK), .QN(n31814) );
  DFF_X1 \REGISTERS_reg[33][59]  ( .D(n9447), .CK(CLK), .QN(n31815) );
  DFF_X1 \REGISTERS_reg[33][58]  ( .D(n9448), .CK(CLK), .QN(n31816) );
  DFF_X1 \REGISTERS_reg[33][57]  ( .D(n9449), .CK(CLK), .QN(n31817) );
  DFF_X1 \REGISTERS_reg[33][56]  ( .D(n9450), .CK(CLK), .QN(n31818) );
  DFF_X1 \REGISTERS_reg[33][55]  ( .D(n9451), .CK(CLK), .QN(n31819) );
  DFF_X1 \REGISTERS_reg[33][54]  ( .D(n9452), .CK(CLK), .QN(n31820) );
  DFF_X1 \REGISTERS_reg[33][53]  ( .D(n9453), .CK(CLK), .QN(n31821) );
  DFF_X1 \REGISTERS_reg[33][52]  ( .D(n9454), .CK(CLK), .QN(n31822) );
  DFF_X1 \REGISTERS_reg[33][51]  ( .D(n9455), .CK(CLK), .QN(n31823) );
  DFF_X1 \REGISTERS_reg[33][50]  ( .D(n9456), .CK(CLK), .QN(n31824) );
  DFF_X1 \REGISTERS_reg[33][49]  ( .D(n9457), .CK(CLK), .QN(n31825) );
  DFF_X1 \REGISTERS_reg[33][48]  ( .D(n9458), .CK(CLK), .QN(n31826) );
  DFF_X1 \REGISTERS_reg[33][47]  ( .D(n9459), .CK(CLK), .QN(n31827) );
  DFF_X1 \REGISTERS_reg[33][46]  ( .D(n9460), .CK(CLK), .QN(n31828) );
  DFF_X1 \REGISTERS_reg[33][45]  ( .D(n9461), .CK(CLK), .QN(n31829) );
  DFF_X1 \REGISTERS_reg[33][44]  ( .D(n9462), .CK(CLK), .QN(n31830) );
  DFF_X1 \REGISTERS_reg[33][43]  ( .D(n9463), .CK(CLK), .QN(n31831) );
  DFF_X1 \REGISTERS_reg[33][42]  ( .D(n9464), .CK(CLK), .QN(n31832) );
  DFF_X1 \REGISTERS_reg[33][41]  ( .D(n9465), .CK(CLK), .QN(n31833) );
  DFF_X1 \REGISTERS_reg[33][40]  ( .D(n9466), .CK(CLK), .QN(n31834) );
  DFF_X1 \REGISTERS_reg[33][39]  ( .D(n9467), .CK(CLK), .QN(n31835) );
  DFF_X1 \REGISTERS_reg[33][38]  ( .D(n9468), .CK(CLK), .QN(n31836) );
  DFF_X1 \REGISTERS_reg[33][37]  ( .D(n9469), .CK(CLK), .QN(n31837) );
  DFF_X1 \REGISTERS_reg[33][36]  ( .D(n9470), .CK(CLK), .QN(n31838) );
  DFF_X1 \REGISTERS_reg[33][35]  ( .D(n9471), .CK(CLK), .QN(n31839) );
  DFF_X1 \REGISTERS_reg[33][34]  ( .D(n9472), .CK(CLK), .QN(n31840) );
  DFF_X1 \REGISTERS_reg[33][33]  ( .D(n9473), .CK(CLK), .QN(n31841) );
  DFF_X1 \REGISTERS_reg[33][32]  ( .D(n9474), .CK(CLK), .QN(n31842) );
  DFF_X1 \REGISTERS_reg[33][31]  ( .D(n9475), .CK(CLK), .QN(n31843) );
  DFF_X1 \REGISTERS_reg[33][30]  ( .D(n9476), .CK(CLK), .QN(n31844) );
  DFF_X1 \REGISTERS_reg[33][29]  ( .D(n9477), .CK(CLK), .QN(n31845) );
  DFF_X1 \REGISTERS_reg[33][28]  ( .D(n9478), .CK(CLK), .QN(n31846) );
  DFF_X1 \REGISTERS_reg[33][27]  ( .D(n9479), .CK(CLK), .QN(n31847) );
  DFF_X1 \REGISTERS_reg[33][26]  ( .D(n9480), .CK(CLK), .QN(n31848) );
  DFF_X1 \REGISTERS_reg[33][25]  ( .D(n9481), .CK(CLK), .QN(n31849) );
  DFF_X1 \REGISTERS_reg[33][24]  ( .D(n9482), .CK(CLK), .QN(n31850) );
  DFF_X1 \REGISTERS_reg[33][23]  ( .D(n9483), .CK(CLK), .QN(n31851) );
  DFF_X1 \REGISTERS_reg[33][22]  ( .D(n9484), .CK(CLK), .QN(n31852) );
  DFF_X1 \REGISTERS_reg[33][21]  ( .D(n9485), .CK(CLK), .QN(n31853) );
  DFF_X1 \REGISTERS_reg[33][20]  ( .D(n9486), .CK(CLK), .QN(n31854) );
  DFF_X1 \REGISTERS_reg[33][19]  ( .D(n9487), .CK(CLK), .QN(n31855) );
  DFF_X1 \REGISTERS_reg[33][18]  ( .D(n9488), .CK(CLK), .QN(n31856) );
  DFF_X1 \REGISTERS_reg[33][17]  ( .D(n9489), .CK(CLK), .QN(n31857) );
  DFF_X1 \REGISTERS_reg[33][16]  ( .D(n9490), .CK(CLK), .QN(n31858) );
  DFF_X1 \REGISTERS_reg[33][15]  ( .D(n9491), .CK(CLK), .QN(n31859) );
  DFF_X1 \REGISTERS_reg[33][14]  ( .D(n9492), .CK(CLK), .QN(n31860) );
  DFF_X1 \REGISTERS_reg[33][13]  ( .D(n9493), .CK(CLK), .QN(n31861) );
  DFF_X1 \REGISTERS_reg[33][12]  ( .D(n9494), .CK(CLK), .QN(n31862) );
  DFF_X1 \REGISTERS_reg[33][11]  ( .D(n9495), .CK(CLK), .QN(n31863) );
  DFF_X1 \REGISTERS_reg[33][10]  ( .D(n9496), .CK(CLK), .QN(n31864) );
  DFF_X1 \REGISTERS_reg[33][9]  ( .D(n9497), .CK(CLK), .QN(n31865) );
  DFF_X1 \REGISTERS_reg[33][8]  ( .D(n9498), .CK(CLK), .QN(n31866) );
  DFF_X1 \REGISTERS_reg[33][7]  ( .D(n9499), .CK(CLK), .QN(n31867) );
  DFF_X1 \REGISTERS_reg[33][6]  ( .D(n9500), .CK(CLK), .QN(n31868) );
  DFF_X1 \REGISTERS_reg[33][5]  ( .D(n9501), .CK(CLK), .QN(n31869) );
  DFF_X1 \REGISTERS_reg[33][4]  ( .D(n9502), .CK(CLK), .QN(n31870) );
  DFF_X1 \REGISTERS_reg[34][63]  ( .D(n9507), .CK(CLK), .QN(n31871) );
  DFF_X1 \REGISTERS_reg[34][62]  ( .D(n9508), .CK(CLK), .QN(n31872) );
  DFF_X1 \REGISTERS_reg[34][61]  ( .D(n9509), .CK(CLK), .QN(n31873) );
  DFF_X1 \REGISTERS_reg[34][60]  ( .D(n9510), .CK(CLK), .QN(n31874) );
  DFF_X1 \REGISTERS_reg[34][59]  ( .D(n9511), .CK(CLK), .QN(n31875) );
  DFF_X1 \REGISTERS_reg[34][58]  ( .D(n9512), .CK(CLK), .QN(n31876) );
  DFF_X1 \REGISTERS_reg[34][57]  ( .D(n9513), .CK(CLK), .QN(n31877) );
  DFF_X1 \REGISTERS_reg[34][56]  ( .D(n9514), .CK(CLK), .QN(n31878) );
  DFF_X1 \REGISTERS_reg[34][55]  ( .D(n9515), .CK(CLK), .QN(n31879) );
  DFF_X1 \REGISTERS_reg[34][54]  ( .D(n9516), .CK(CLK), .QN(n31880) );
  DFF_X1 \REGISTERS_reg[34][53]  ( .D(n9517), .CK(CLK), .QN(n31881) );
  DFF_X1 \REGISTERS_reg[34][52]  ( .D(n9518), .CK(CLK), .QN(n31882) );
  DFF_X1 \REGISTERS_reg[34][51]  ( .D(n9519), .CK(CLK), .QN(n31883) );
  DFF_X1 \REGISTERS_reg[34][50]  ( .D(n9520), .CK(CLK), .QN(n31884) );
  DFF_X1 \REGISTERS_reg[34][49]  ( .D(n9521), .CK(CLK), .QN(n31885) );
  DFF_X1 \REGISTERS_reg[34][48]  ( .D(n9522), .CK(CLK), .QN(n31886) );
  DFF_X1 \REGISTERS_reg[34][47]  ( .D(n9523), .CK(CLK), .QN(n31887) );
  DFF_X1 \REGISTERS_reg[34][46]  ( .D(n9524), .CK(CLK), .QN(n31888) );
  DFF_X1 \REGISTERS_reg[34][45]  ( .D(n9525), .CK(CLK), .QN(n31889) );
  DFF_X1 \REGISTERS_reg[34][44]  ( .D(n9526), .CK(CLK), .QN(n31890) );
  DFF_X1 \REGISTERS_reg[34][43]  ( .D(n9527), .CK(CLK), .QN(n31891) );
  DFF_X1 \REGISTERS_reg[34][42]  ( .D(n9528), .CK(CLK), .QN(n31892) );
  DFF_X1 \REGISTERS_reg[34][41]  ( .D(n9529), .CK(CLK), .QN(n31893) );
  DFF_X1 \REGISTERS_reg[34][40]  ( .D(n9530), .CK(CLK), .QN(n31894) );
  DFF_X1 \REGISTERS_reg[34][39]  ( .D(n9531), .CK(CLK), .QN(n31895) );
  DFF_X1 \REGISTERS_reg[34][38]  ( .D(n9532), .CK(CLK), .QN(n31896) );
  DFF_X1 \REGISTERS_reg[34][37]  ( .D(n9533), .CK(CLK), .QN(n31897) );
  DFF_X1 \REGISTERS_reg[34][36]  ( .D(n9534), .CK(CLK), .QN(n31898) );
  DFF_X1 \REGISTERS_reg[34][35]  ( .D(n9535), .CK(CLK), .QN(n31899) );
  DFF_X1 \REGISTERS_reg[34][34]  ( .D(n9536), .CK(CLK), .QN(n31900) );
  DFF_X1 \REGISTERS_reg[34][33]  ( .D(n9537), .CK(CLK), .QN(n31901) );
  DFF_X1 \REGISTERS_reg[34][32]  ( .D(n9538), .CK(CLK), .QN(n31902) );
  DFF_X1 \REGISTERS_reg[34][31]  ( .D(n9539), .CK(CLK), .QN(n31903) );
  DFF_X1 \REGISTERS_reg[34][30]  ( .D(n9540), .CK(CLK), .QN(n31904) );
  DFF_X1 \REGISTERS_reg[34][29]  ( .D(n9541), .CK(CLK), .QN(n31905) );
  DFF_X1 \REGISTERS_reg[34][28]  ( .D(n9542), .CK(CLK), .QN(n31906) );
  DFF_X1 \REGISTERS_reg[34][27]  ( .D(n9543), .CK(CLK), .QN(n31907) );
  DFF_X1 \REGISTERS_reg[34][26]  ( .D(n9544), .CK(CLK), .QN(n31908) );
  DFF_X1 \REGISTERS_reg[34][25]  ( .D(n9545), .CK(CLK), .QN(n31909) );
  DFF_X1 \REGISTERS_reg[34][24]  ( .D(n9546), .CK(CLK), .QN(n31910) );
  DFF_X1 \REGISTERS_reg[34][23]  ( .D(n9547), .CK(CLK), .QN(n31911) );
  DFF_X1 \REGISTERS_reg[34][22]  ( .D(n9548), .CK(CLK), .QN(n31912) );
  DFF_X1 \REGISTERS_reg[34][21]  ( .D(n9549), .CK(CLK), .QN(n31913) );
  DFF_X1 \REGISTERS_reg[34][20]  ( .D(n9550), .CK(CLK), .QN(n31914) );
  DFF_X1 \REGISTERS_reg[34][19]  ( .D(n9551), .CK(CLK), .QN(n31915) );
  DFF_X1 \REGISTERS_reg[34][18]  ( .D(n9552), .CK(CLK), .QN(n31916) );
  DFF_X1 \REGISTERS_reg[34][17]  ( .D(n9553), .CK(CLK), .QN(n31917) );
  DFF_X1 \REGISTERS_reg[34][16]  ( .D(n9554), .CK(CLK), .QN(n31918) );
  DFF_X1 \REGISTERS_reg[34][15]  ( .D(n9555), .CK(CLK), .QN(n31919) );
  DFF_X1 \REGISTERS_reg[34][14]  ( .D(n9556), .CK(CLK), .QN(n31920) );
  DFF_X1 \REGISTERS_reg[34][13]  ( .D(n9557), .CK(CLK), .QN(n31921) );
  DFF_X1 \REGISTERS_reg[34][12]  ( .D(n9558), .CK(CLK), .QN(n31922) );
  DFF_X1 \REGISTERS_reg[34][11]  ( .D(n9559), .CK(CLK), .QN(n31923) );
  DFF_X1 \REGISTERS_reg[34][10]  ( .D(n9560), .CK(CLK), .QN(n31924) );
  DFF_X1 \REGISTERS_reg[34][9]  ( .D(n9561), .CK(CLK), .QN(n31925) );
  DFF_X1 \REGISTERS_reg[34][8]  ( .D(n9562), .CK(CLK), .QN(n31926) );
  DFF_X1 \REGISTERS_reg[34][7]  ( .D(n9563), .CK(CLK), .QN(n31927) );
  DFF_X1 \REGISTERS_reg[34][6]  ( .D(n9564), .CK(CLK), .QN(n31928) );
  DFF_X1 \REGISTERS_reg[34][5]  ( .D(n9565), .CK(CLK), .QN(n31929) );
  DFF_X1 \REGISTERS_reg[34][4]  ( .D(n9566), .CK(CLK), .QN(n31930) );
  DFF_X1 \REGISTERS_reg[37][63]  ( .D(n9699), .CK(CLK), .QN(n31931) );
  DFF_X1 \REGISTERS_reg[37][62]  ( .D(n9700), .CK(CLK), .QN(n31932) );
  DFF_X1 \REGISTERS_reg[37][61]  ( .D(n9701), .CK(CLK), .QN(n31933) );
  DFF_X1 \REGISTERS_reg[37][60]  ( .D(n9702), .CK(CLK), .QN(n31934) );
  DFF_X1 \REGISTERS_reg[37][59]  ( .D(n9703), .CK(CLK), .QN(n31935) );
  DFF_X1 \REGISTERS_reg[37][58]  ( .D(n9704), .CK(CLK), .QN(n31936) );
  DFF_X1 \REGISTERS_reg[37][57]  ( .D(n9705), .CK(CLK), .QN(n31937) );
  DFF_X1 \REGISTERS_reg[37][56]  ( .D(n9706), .CK(CLK), .QN(n31938) );
  DFF_X1 \REGISTERS_reg[37][55]  ( .D(n9707), .CK(CLK), .QN(n31939) );
  DFF_X1 \REGISTERS_reg[37][54]  ( .D(n9708), .CK(CLK), .QN(n31940) );
  DFF_X1 \REGISTERS_reg[37][53]  ( .D(n9709), .CK(CLK), .QN(n31941) );
  DFF_X1 \REGISTERS_reg[37][52]  ( .D(n9710), .CK(CLK), .QN(n31942) );
  DFF_X1 \REGISTERS_reg[37][51]  ( .D(n9711), .CK(CLK), .QN(n31943) );
  DFF_X1 \REGISTERS_reg[37][50]  ( .D(n9712), .CK(CLK), .QN(n31944) );
  DFF_X1 \REGISTERS_reg[37][49]  ( .D(n9713), .CK(CLK), .QN(n31945) );
  DFF_X1 \REGISTERS_reg[37][48]  ( .D(n9714), .CK(CLK), .QN(n31946) );
  DFF_X1 \REGISTERS_reg[37][47]  ( .D(n9715), .CK(CLK), .QN(n31947) );
  DFF_X1 \REGISTERS_reg[37][46]  ( .D(n9716), .CK(CLK), .QN(n31948) );
  DFF_X1 \REGISTERS_reg[37][45]  ( .D(n9717), .CK(CLK), .QN(n31949) );
  DFF_X1 \REGISTERS_reg[37][44]  ( .D(n9718), .CK(CLK), .QN(n31950) );
  DFF_X1 \REGISTERS_reg[37][43]  ( .D(n9719), .CK(CLK), .QN(n31951) );
  DFF_X1 \REGISTERS_reg[37][42]  ( .D(n9720), .CK(CLK), .QN(n31952) );
  DFF_X1 \REGISTERS_reg[37][41]  ( .D(n9721), .CK(CLK), .QN(n31953) );
  DFF_X1 \REGISTERS_reg[37][40]  ( .D(n9722), .CK(CLK), .QN(n31954) );
  DFF_X1 \REGISTERS_reg[37][39]  ( .D(n9723), .CK(CLK), .QN(n31955) );
  DFF_X1 \REGISTERS_reg[37][38]  ( .D(n9724), .CK(CLK), .QN(n31956) );
  DFF_X1 \REGISTERS_reg[37][37]  ( .D(n9725), .CK(CLK), .QN(n31957) );
  DFF_X1 \REGISTERS_reg[37][36]  ( .D(n9726), .CK(CLK), .QN(n31958) );
  DFF_X1 \REGISTERS_reg[37][35]  ( .D(n9727), .CK(CLK), .QN(n31959) );
  DFF_X1 \REGISTERS_reg[37][34]  ( .D(n9728), .CK(CLK), .QN(n31960) );
  DFF_X1 \REGISTERS_reg[37][33]  ( .D(n9729), .CK(CLK), .QN(n31961) );
  DFF_X1 \REGISTERS_reg[37][32]  ( .D(n9730), .CK(CLK), .QN(n31962) );
  DFF_X1 \REGISTERS_reg[37][31]  ( .D(n9731), .CK(CLK), .QN(n31963) );
  DFF_X1 \REGISTERS_reg[37][30]  ( .D(n9732), .CK(CLK), .QN(n31964) );
  DFF_X1 \REGISTERS_reg[37][29]  ( .D(n9733), .CK(CLK), .QN(n31965) );
  DFF_X1 \REGISTERS_reg[37][28]  ( .D(n9734), .CK(CLK), .QN(n31966) );
  DFF_X1 \REGISTERS_reg[37][27]  ( .D(n9735), .CK(CLK), .QN(n31967) );
  DFF_X1 \REGISTERS_reg[37][26]  ( .D(n9736), .CK(CLK), .QN(n31968) );
  DFF_X1 \REGISTERS_reg[37][25]  ( .D(n9737), .CK(CLK), .QN(n31969) );
  DFF_X1 \REGISTERS_reg[37][24]  ( .D(n9738), .CK(CLK), .QN(n31970) );
  DFF_X1 \REGISTERS_reg[37][23]  ( .D(n9739), .CK(CLK), .QN(n31971) );
  DFF_X1 \REGISTERS_reg[37][22]  ( .D(n9740), .CK(CLK), .QN(n31972) );
  DFF_X1 \REGISTERS_reg[37][21]  ( .D(n9741), .CK(CLK), .QN(n31973) );
  DFF_X1 \REGISTERS_reg[37][20]  ( .D(n9742), .CK(CLK), .QN(n31974) );
  DFF_X1 \REGISTERS_reg[37][19]  ( .D(n9743), .CK(CLK), .QN(n31975) );
  DFF_X1 \REGISTERS_reg[37][18]  ( .D(n9744), .CK(CLK), .QN(n31976) );
  DFF_X1 \REGISTERS_reg[37][17]  ( .D(n9745), .CK(CLK), .QN(n31977) );
  DFF_X1 \REGISTERS_reg[37][16]  ( .D(n9746), .CK(CLK), .QN(n31978) );
  DFF_X1 \REGISTERS_reg[37][15]  ( .D(n9747), .CK(CLK), .QN(n31979) );
  DFF_X1 \REGISTERS_reg[37][14]  ( .D(n9748), .CK(CLK), .QN(n31980) );
  DFF_X1 \REGISTERS_reg[37][13]  ( .D(n9749), .CK(CLK), .QN(n31981) );
  DFF_X1 \REGISTERS_reg[37][12]  ( .D(n9750), .CK(CLK), .QN(n31982) );
  DFF_X1 \REGISTERS_reg[37][11]  ( .D(n9751), .CK(CLK), .QN(n31983) );
  DFF_X1 \REGISTERS_reg[37][10]  ( .D(n9752), .CK(CLK), .QN(n31984) );
  DFF_X1 \REGISTERS_reg[37][9]  ( .D(n9753), .CK(CLK), .QN(n31985) );
  DFF_X1 \REGISTERS_reg[37][8]  ( .D(n9754), .CK(CLK), .QN(n31986) );
  DFF_X1 \REGISTERS_reg[37][7]  ( .D(n9755), .CK(CLK), .QN(n31987) );
  DFF_X1 \REGISTERS_reg[37][6]  ( .D(n9756), .CK(CLK), .QN(n31988) );
  DFF_X1 \REGISTERS_reg[37][5]  ( .D(n9757), .CK(CLK), .QN(n31989) );
  DFF_X1 \REGISTERS_reg[37][4]  ( .D(n9758), .CK(CLK), .QN(n31990) );
  DFF_X1 \REGISTERS_reg[38][63]  ( .D(n9763), .CK(CLK), .QN(n31991) );
  DFF_X1 \REGISTERS_reg[38][62]  ( .D(n9764), .CK(CLK), .QN(n31992) );
  DFF_X1 \REGISTERS_reg[38][61]  ( .D(n9765), .CK(CLK), .QN(n31993) );
  DFF_X1 \REGISTERS_reg[38][60]  ( .D(n9766), .CK(CLK), .QN(n31994) );
  DFF_X1 \REGISTERS_reg[38][59]  ( .D(n9767), .CK(CLK), .QN(n31995) );
  DFF_X1 \REGISTERS_reg[38][58]  ( .D(n9768), .CK(CLK), .QN(n31996) );
  DFF_X1 \REGISTERS_reg[38][57]  ( .D(n9769), .CK(CLK), .QN(n31997) );
  DFF_X1 \REGISTERS_reg[38][56]  ( .D(n9770), .CK(CLK), .QN(n31998) );
  DFF_X1 \REGISTERS_reg[38][55]  ( .D(n9771), .CK(CLK), .QN(n31999) );
  DFF_X1 \REGISTERS_reg[38][54]  ( .D(n9772), .CK(CLK), .QN(n32000) );
  DFF_X1 \REGISTERS_reg[38][53]  ( .D(n9773), .CK(CLK), .QN(n32001) );
  DFF_X1 \REGISTERS_reg[38][52]  ( .D(n9774), .CK(CLK), .QN(n32002) );
  DFF_X1 \REGISTERS_reg[38][51]  ( .D(n9775), .CK(CLK), .QN(n32003) );
  DFF_X1 \REGISTERS_reg[38][50]  ( .D(n9776), .CK(CLK), .QN(n32004) );
  DFF_X1 \REGISTERS_reg[38][49]  ( .D(n9777), .CK(CLK), .QN(n32005) );
  DFF_X1 \REGISTERS_reg[38][48]  ( .D(n9778), .CK(CLK), .QN(n32006) );
  DFF_X1 \REGISTERS_reg[38][47]  ( .D(n9779), .CK(CLK), .QN(n32007) );
  DFF_X1 \REGISTERS_reg[38][46]  ( .D(n9780), .CK(CLK), .QN(n32008) );
  DFF_X1 \REGISTERS_reg[38][45]  ( .D(n9781), .CK(CLK), .QN(n32009) );
  DFF_X1 \REGISTERS_reg[38][44]  ( .D(n9782), .CK(CLK), .QN(n32010) );
  DFF_X1 \REGISTERS_reg[38][43]  ( .D(n9783), .CK(CLK), .QN(n32011) );
  DFF_X1 \REGISTERS_reg[38][42]  ( .D(n9784), .CK(CLK), .QN(n32012) );
  DFF_X1 \REGISTERS_reg[38][41]  ( .D(n9785), .CK(CLK), .QN(n32013) );
  DFF_X1 \REGISTERS_reg[38][40]  ( .D(n9786), .CK(CLK), .QN(n32014) );
  DFF_X1 \REGISTERS_reg[38][39]  ( .D(n9787), .CK(CLK), .QN(n32015) );
  DFF_X1 \REGISTERS_reg[38][38]  ( .D(n9788), .CK(CLK), .QN(n32016) );
  DFF_X1 \REGISTERS_reg[38][37]  ( .D(n9789), .CK(CLK), .QN(n32017) );
  DFF_X1 \REGISTERS_reg[38][36]  ( .D(n9790), .CK(CLK), .QN(n32018) );
  DFF_X1 \REGISTERS_reg[38][35]  ( .D(n9791), .CK(CLK), .QN(n32019) );
  DFF_X1 \REGISTERS_reg[38][34]  ( .D(n9792), .CK(CLK), .QN(n32020) );
  DFF_X1 \REGISTERS_reg[38][33]  ( .D(n9793), .CK(CLK), .QN(n32021) );
  DFF_X1 \REGISTERS_reg[38][32]  ( .D(n9794), .CK(CLK), .QN(n32022) );
  DFF_X1 \REGISTERS_reg[38][31]  ( .D(n9795), .CK(CLK), .QN(n32023) );
  DFF_X1 \REGISTERS_reg[38][30]  ( .D(n9796), .CK(CLK), .QN(n32024) );
  DFF_X1 \REGISTERS_reg[38][29]  ( .D(n9797), .CK(CLK), .QN(n32025) );
  DFF_X1 \REGISTERS_reg[38][28]  ( .D(n9798), .CK(CLK), .QN(n32026) );
  DFF_X1 \REGISTERS_reg[38][27]  ( .D(n9799), .CK(CLK), .QN(n32027) );
  DFF_X1 \REGISTERS_reg[38][26]  ( .D(n9800), .CK(CLK), .QN(n32028) );
  DFF_X1 \REGISTERS_reg[38][25]  ( .D(n9801), .CK(CLK), .QN(n32029) );
  DFF_X1 \REGISTERS_reg[38][24]  ( .D(n9802), .CK(CLK), .QN(n32030) );
  DFF_X1 \REGISTERS_reg[38][23]  ( .D(n9803), .CK(CLK), .QN(n32031) );
  DFF_X1 \REGISTERS_reg[38][22]  ( .D(n9804), .CK(CLK), .QN(n32032) );
  DFF_X1 \REGISTERS_reg[38][21]  ( .D(n9805), .CK(CLK), .QN(n32033) );
  DFF_X1 \REGISTERS_reg[38][20]  ( .D(n9806), .CK(CLK), .QN(n32034) );
  DFF_X1 \REGISTERS_reg[38][19]  ( .D(n9807), .CK(CLK), .QN(n32035) );
  DFF_X1 \REGISTERS_reg[38][18]  ( .D(n9808), .CK(CLK), .QN(n32036) );
  DFF_X1 \REGISTERS_reg[38][17]  ( .D(n9809), .CK(CLK), .QN(n32037) );
  DFF_X1 \REGISTERS_reg[38][16]  ( .D(n9810), .CK(CLK), .QN(n32038) );
  DFF_X1 \REGISTERS_reg[38][15]  ( .D(n9811), .CK(CLK), .QN(n32039) );
  DFF_X1 \REGISTERS_reg[38][14]  ( .D(n9812), .CK(CLK), .QN(n32040) );
  DFF_X1 \REGISTERS_reg[38][13]  ( .D(n9813), .CK(CLK), .QN(n32041) );
  DFF_X1 \REGISTERS_reg[38][12]  ( .D(n9814), .CK(CLK), .QN(n32042) );
  DFF_X1 \REGISTERS_reg[38][11]  ( .D(n9815), .CK(CLK), .QN(n32043) );
  DFF_X1 \REGISTERS_reg[38][10]  ( .D(n9816), .CK(CLK), .QN(n32044) );
  DFF_X1 \REGISTERS_reg[38][9]  ( .D(n9817), .CK(CLK), .QN(n32045) );
  DFF_X1 \REGISTERS_reg[38][8]  ( .D(n9818), .CK(CLK), .QN(n32046) );
  DFF_X1 \REGISTERS_reg[38][7]  ( .D(n9819), .CK(CLK), .QN(n32047) );
  DFF_X1 \REGISTERS_reg[38][6]  ( .D(n9820), .CK(CLK), .QN(n32048) );
  DFF_X1 \REGISTERS_reg[38][5]  ( .D(n9821), .CK(CLK), .QN(n32049) );
  DFF_X1 \REGISTERS_reg[38][4]  ( .D(n9822), .CK(CLK), .QN(n32050) );
  DFF_X1 \REGISTERS_reg[39][63]  ( .D(n9827), .CK(CLK), .QN(n32051) );
  DFF_X1 \OUT2_reg[63]  ( .D(n7203), .CK(CLK), .Q(OUT2[63]), .QN(n16942) );
  DFF_X1 \OUT1_reg[63]  ( .D(n7267), .CK(CLK), .Q(OUT1[63]), .QN(n17006) );
  DFF_X1 \REGISTERS_reg[39][62]  ( .D(n9828), .CK(CLK), .QN(n32052) );
  DFF_X1 \OUT2_reg[62]  ( .D(n7204), .CK(CLK), .Q(OUT2[62]), .QN(n16943) );
  DFF_X1 \OUT1_reg[62]  ( .D(n7268), .CK(CLK), .Q(OUT1[62]), .QN(n17007) );
  DFF_X1 \REGISTERS_reg[39][61]  ( .D(n9829), .CK(CLK), .QN(n32053) );
  DFF_X1 \OUT2_reg[61]  ( .D(n7205), .CK(CLK), .Q(OUT2[61]), .QN(n16944) );
  DFF_X1 \OUT1_reg[61]  ( .D(n7269), .CK(CLK), .Q(OUT1[61]), .QN(n17008) );
  DFF_X1 \OUT2_reg[60]  ( .D(n7206), .CK(CLK), .Q(OUT2[60]), .QN(n16945) );
  DFF_X1 \OUT1_reg[60]  ( .D(n7270), .CK(CLK), .Q(OUT1[60]), .QN(n17009) );
  DFF_X1 \REGISTERS_reg[39][59]  ( .D(n9831), .CK(CLK), .QN(n32054) );
  DFF_X1 \OUT2_reg[59]  ( .D(n7207), .CK(CLK), .Q(OUT2[59]), .QN(n16946) );
  DFF_X1 \OUT1_reg[59]  ( .D(n7271), .CK(CLK), .Q(OUT1[59]), .QN(n17010) );
  DFF_X1 \OUT2_reg[58]  ( .D(n7208), .CK(CLK), .Q(OUT2[58]), .QN(n16947) );
  DFF_X1 \OUT1_reg[58]  ( .D(n7272), .CK(CLK), .Q(OUT1[58]), .QN(n17011) );
  DFF_X1 \OUT2_reg[57]  ( .D(n7209), .CK(CLK), .Q(OUT2[57]), .QN(n16948) );
  DFF_X1 \OUT1_reg[57]  ( .D(n7273), .CK(CLK), .Q(OUT1[57]), .QN(n17012) );
  DFF_X1 \OUT2_reg[56]  ( .D(n7210), .CK(CLK), .Q(OUT2[56]), .QN(n16949) );
  DFF_X1 \OUT1_reg[56]  ( .D(n7274), .CK(CLK), .Q(OUT1[56]), .QN(n17013) );
  DFF_X1 \OUT2_reg[55]  ( .D(n7211), .CK(CLK), .Q(OUT2[55]), .QN(n16950) );
  DFF_X1 \OUT1_reg[55]  ( .D(n7275), .CK(CLK), .Q(OUT1[55]), .QN(n17014) );
  DFF_X1 \OUT2_reg[54]  ( .D(n7212), .CK(CLK), .Q(OUT2[54]), .QN(n16951) );
  DFF_X1 \OUT1_reg[54]  ( .D(n7276), .CK(CLK), .Q(OUT1[54]), .QN(n17015) );
  DFF_X1 \OUT2_reg[53]  ( .D(n7213), .CK(CLK), .Q(OUT2[53]), .QN(n16952) );
  DFF_X1 \OUT1_reg[53]  ( .D(n7277), .CK(CLK), .Q(OUT1[53]), .QN(n17016) );
  DFF_X1 \OUT2_reg[52]  ( .D(n7214), .CK(CLK), .Q(OUT2[52]), .QN(n16953) );
  DFF_X1 \OUT1_reg[52]  ( .D(n7278), .CK(CLK), .Q(OUT1[52]), .QN(n17017) );
  DFF_X1 \OUT2_reg[51]  ( .D(n7215), .CK(CLK), .Q(OUT2[51]), .QN(n16954) );
  DFF_X1 \OUT1_reg[51]  ( .D(n7279), .CK(CLK), .Q(OUT1[51]), .QN(n17018) );
  DFF_X1 \OUT2_reg[50]  ( .D(n7216), .CK(CLK), .Q(OUT2[50]), .QN(n16955) );
  DFF_X1 \OUT1_reg[50]  ( .D(n7280), .CK(CLK), .Q(OUT1[50]), .QN(n17019) );
  DFF_X1 \OUT2_reg[49]  ( .D(n7217), .CK(CLK), .Q(OUT2[49]), .QN(n16956) );
  DFF_X1 \OUT1_reg[49]  ( .D(n7281), .CK(CLK), .Q(OUT1[49]), .QN(n17020) );
  DFF_X1 \OUT2_reg[48]  ( .D(n7218), .CK(CLK), .Q(OUT2[48]), .QN(n16957) );
  DFF_X1 \OUT1_reg[48]  ( .D(n7282), .CK(CLK), .Q(OUT1[48]), .QN(n17021) );
  DFF_X1 \OUT2_reg[47]  ( .D(n7219), .CK(CLK), .Q(OUT2[47]), .QN(n16958) );
  DFF_X1 \OUT1_reg[47]  ( .D(n7283), .CK(CLK), .Q(OUT1[47]), .QN(n17022) );
  DFF_X1 \OUT2_reg[46]  ( .D(n7220), .CK(CLK), .Q(OUT2[46]), .QN(n16959) );
  DFF_X1 \OUT1_reg[46]  ( .D(n7284), .CK(CLK), .Q(OUT1[46]), .QN(n17023) );
  DFF_X1 \OUT2_reg[45]  ( .D(n7221), .CK(CLK), .Q(OUT2[45]), .QN(n16960) );
  DFF_X1 \OUT1_reg[45]  ( .D(n7285), .CK(CLK), .Q(OUT1[45]), .QN(n17024) );
  DFF_X1 \OUT2_reg[44]  ( .D(n7222), .CK(CLK), .Q(OUT2[44]), .QN(n16961) );
  DFF_X1 \OUT1_reg[44]  ( .D(n7286), .CK(CLK), .Q(OUT1[44]), .QN(n17025) );
  DFF_X1 \OUT2_reg[43]  ( .D(n7223), .CK(CLK), .Q(OUT2[43]), .QN(n16962) );
  DFF_X1 \OUT1_reg[43]  ( .D(n7287), .CK(CLK), .Q(OUT1[43]), .QN(n17026) );
  DFF_X1 \OUT2_reg[42]  ( .D(n7224), .CK(CLK), .Q(OUT2[42]), .QN(n16963) );
  DFF_X1 \OUT1_reg[42]  ( .D(n7288), .CK(CLK), .Q(OUT1[42]), .QN(n17027) );
  DFF_X1 \OUT2_reg[41]  ( .D(n7225), .CK(CLK), .Q(OUT2[41]), .QN(n16964) );
  DFF_X1 \OUT1_reg[41]  ( .D(n7289), .CK(CLK), .Q(OUT1[41]), .QN(n17028) );
  DFF_X1 \OUT2_reg[40]  ( .D(n7226), .CK(CLK), .Q(OUT2[40]), .QN(n16965) );
  DFF_X1 \OUT1_reg[40]  ( .D(n7290), .CK(CLK), .Q(OUT1[40]), .QN(n17029) );
  DFF_X1 \OUT2_reg[39]  ( .D(n7227), .CK(CLK), .Q(OUT2[39]), .QN(n16966) );
  DFF_X1 \OUT1_reg[39]  ( .D(n7291), .CK(CLK), .Q(OUT1[39]), .QN(n17030) );
  DFF_X1 \OUT2_reg[38]  ( .D(n7228), .CK(CLK), .Q(OUT2[38]), .QN(n16967) );
  DFF_X1 \OUT1_reg[38]  ( .D(n7292), .CK(CLK), .Q(OUT1[38]), .QN(n17031) );
  DFF_X1 \OUT2_reg[37]  ( .D(n7229), .CK(CLK), .Q(OUT2[37]), .QN(n16968) );
  DFF_X1 \OUT1_reg[37]  ( .D(n7293), .CK(CLK), .Q(OUT1[37]), .QN(n17032) );
  DFF_X1 \OUT2_reg[36]  ( .D(n7230), .CK(CLK), .Q(OUT2[36]), .QN(n16969) );
  DFF_X1 \OUT1_reg[36]  ( .D(n7294), .CK(CLK), .Q(OUT1[36]), .QN(n17033) );
  DFF_X1 \OUT2_reg[35]  ( .D(n7231), .CK(CLK), .Q(OUT2[35]), .QN(n16970) );
  DFF_X1 \OUT1_reg[35]  ( .D(n7295), .CK(CLK), .Q(OUT1[35]), .QN(n17034) );
  DFF_X1 \OUT2_reg[34]  ( .D(n7232), .CK(CLK), .Q(OUT2[34]), .QN(n16971) );
  DFF_X1 \OUT1_reg[34]  ( .D(n7296), .CK(CLK), .Q(OUT1[34]), .QN(n17035) );
  DFF_X1 \OUT2_reg[33]  ( .D(n7233), .CK(CLK), .Q(OUT2[33]), .QN(n16972) );
  DFF_X1 \OUT1_reg[33]  ( .D(n7297), .CK(CLK), .Q(OUT1[33]), .QN(n17036) );
  DFF_X1 \OUT2_reg[32]  ( .D(n7234), .CK(CLK), .Q(OUT2[32]), .QN(n16973) );
  DFF_X1 \OUT1_reg[32]  ( .D(n7298), .CK(CLK), .Q(OUT1[32]), .QN(n17037) );
  DFF_X1 \OUT2_reg[31]  ( .D(n7235), .CK(CLK), .Q(OUT2[31]), .QN(n16974) );
  DFF_X1 \OUT1_reg[31]  ( .D(n7299), .CK(CLK), .Q(OUT1[31]), .QN(n17038) );
  DFF_X1 \OUT2_reg[30]  ( .D(n7236), .CK(CLK), .Q(OUT2[30]), .QN(n16975) );
  DFF_X1 \OUT1_reg[30]  ( .D(n7300), .CK(CLK), .Q(OUT1[30]), .QN(n17039) );
  DFF_X1 \OUT2_reg[29]  ( .D(n7237), .CK(CLK), .Q(OUT2[29]), .QN(n16976) );
  DFF_X1 \OUT1_reg[29]  ( .D(n7301), .CK(CLK), .Q(OUT1[29]), .QN(n17040) );
  DFF_X1 \OUT2_reg[28]  ( .D(n7238), .CK(CLK), .Q(OUT2[28]), .QN(n16977) );
  DFF_X1 \OUT1_reg[28]  ( .D(n7302), .CK(CLK), .Q(OUT1[28]), .QN(n17041) );
  DFF_X1 \OUT2_reg[27]  ( .D(n7239), .CK(CLK), .Q(OUT2[27]), .QN(n16978) );
  DFF_X1 \OUT1_reg[27]  ( .D(n7303), .CK(CLK), .Q(OUT1[27]), .QN(n17042) );
  DFF_X1 \OUT2_reg[26]  ( .D(n7240), .CK(CLK), .Q(OUT2[26]), .QN(n16979) );
  DFF_X1 \OUT1_reg[26]  ( .D(n7304), .CK(CLK), .Q(OUT1[26]), .QN(n17043) );
  DFF_X1 \OUT2_reg[25]  ( .D(n7241), .CK(CLK), .Q(OUT2[25]), .QN(n16980) );
  DFF_X1 \OUT1_reg[25]  ( .D(n7305), .CK(CLK), .Q(OUT1[25]), .QN(n17044) );
  DFF_X1 \OUT2_reg[24]  ( .D(n7242), .CK(CLK), .Q(OUT2[24]), .QN(n16981) );
  DFF_X1 \OUT1_reg[24]  ( .D(n7306), .CK(CLK), .Q(OUT1[24]), .QN(n17045) );
  DFF_X1 \REGISTERS_reg[39][23]  ( .D(n9867), .CK(CLK), .QN(n32055) );
  DFF_X1 \OUT2_reg[23]  ( .D(n7243), .CK(CLK), .Q(OUT2[23]), .QN(n16982) );
  DFF_X1 \OUT1_reg[23]  ( .D(n7307), .CK(CLK), .Q(OUT1[23]), .QN(n17046) );
  DFF_X1 \REGISTERS_reg[39][22]  ( .D(n9868), .CK(CLK), .QN(n32056) );
  DFF_X1 \OUT2_reg[22]  ( .D(n7244), .CK(CLK), .Q(OUT2[22]), .QN(n16983) );
  DFF_X1 \OUT1_reg[22]  ( .D(n7308), .CK(CLK), .Q(OUT1[22]), .QN(n17047) );
  DFF_X1 \REGISTERS_reg[39][21]  ( .D(n9869), .CK(CLK), .QN(n32057) );
  DFF_X1 \OUT2_reg[21]  ( .D(n7245), .CK(CLK), .Q(OUT2[21]), .QN(n16984) );
  DFF_X1 \OUT1_reg[21]  ( .D(n7309), .CK(CLK), .Q(OUT1[21]), .QN(n17048) );
  DFF_X1 \REGISTERS_reg[39][20]  ( .D(n9870), .CK(CLK), .QN(n32058) );
  DFF_X1 \OUT2_reg[20]  ( .D(n7246), .CK(CLK), .Q(OUT2[20]), .QN(n16985) );
  DFF_X1 \OUT1_reg[20]  ( .D(n7310), .CK(CLK), .Q(OUT1[20]), .QN(n17049) );
  DFF_X1 \REGISTERS_reg[39][19]  ( .D(n9871), .CK(CLK), .QN(n32059) );
  DFF_X1 \OUT2_reg[19]  ( .D(n7247), .CK(CLK), .Q(OUT2[19]), .QN(n16986) );
  DFF_X1 \OUT1_reg[19]  ( .D(n7311), .CK(CLK), .Q(OUT1[19]), .QN(n17050) );
  DFF_X1 \REGISTERS_reg[39][18]  ( .D(n9872), .CK(CLK), .QN(n32060) );
  DFF_X1 \OUT2_reg[18]  ( .D(n7248), .CK(CLK), .Q(OUT2[18]), .QN(n16987) );
  DFF_X1 \OUT1_reg[18]  ( .D(n7312), .CK(CLK), .Q(OUT1[18]), .QN(n17051) );
  DFF_X1 \REGISTERS_reg[39][17]  ( .D(n9873), .CK(CLK), .QN(n32061) );
  DFF_X1 \OUT2_reg[17]  ( .D(n7249), .CK(CLK), .Q(OUT2[17]), .QN(n16988) );
  DFF_X1 \OUT1_reg[17]  ( .D(n7313), .CK(CLK), .Q(OUT1[17]), .QN(n17052) );
  DFF_X1 \REGISTERS_reg[39][16]  ( .D(n9874), .CK(CLK), .QN(n32062) );
  DFF_X1 \OUT2_reg[16]  ( .D(n7250), .CK(CLK), .Q(OUT2[16]), .QN(n16989) );
  DFF_X1 \OUT1_reg[16]  ( .D(n7314), .CK(CLK), .Q(OUT1[16]), .QN(n17053) );
  DFF_X1 \REGISTERS_reg[39][15]  ( .D(n9875), .CK(CLK), .QN(n32063) );
  DFF_X1 \OUT2_reg[15]  ( .D(n7251), .CK(CLK), .Q(OUT2[15]), .QN(n16990) );
  DFF_X1 \OUT1_reg[15]  ( .D(n7315), .CK(CLK), .Q(OUT1[15]), .QN(n17054) );
  DFF_X1 \REGISTERS_reg[39][14]  ( .D(n9876), .CK(CLK), .QN(n32064) );
  DFF_X1 \OUT2_reg[14]  ( .D(n7252), .CK(CLK), .Q(OUT2[14]), .QN(n16991) );
  DFF_X1 \OUT1_reg[14]  ( .D(n7316), .CK(CLK), .Q(OUT1[14]), .QN(n17055) );
  DFF_X1 \REGISTERS_reg[39][13]  ( .D(n9877), .CK(CLK), .QN(n32065) );
  DFF_X1 \OUT2_reg[13]  ( .D(n7253), .CK(CLK), .Q(OUT2[13]), .QN(n16992) );
  DFF_X1 \OUT1_reg[13]  ( .D(n7317), .CK(CLK), .Q(OUT1[13]), .QN(n17056) );
  DFF_X1 \REGISTERS_reg[39][12]  ( .D(n9878), .CK(CLK), .QN(n32066) );
  DFF_X1 \OUT2_reg[12]  ( .D(n7254), .CK(CLK), .Q(OUT2[12]), .QN(n16993) );
  DFF_X1 \OUT1_reg[12]  ( .D(n7318), .CK(CLK), .Q(OUT1[12]), .QN(n17057) );
  DFF_X1 \REGISTERS_reg[39][11]  ( .D(n9879), .CK(CLK), .QN(n32067) );
  DFF_X1 \OUT2_reg[11]  ( .D(n7255), .CK(CLK), .Q(OUT2[11]), .QN(n16994) );
  DFF_X1 \OUT1_reg[11]  ( .D(n7319), .CK(CLK), .Q(OUT1[11]), .QN(n17058) );
  DFF_X1 \REGISTERS_reg[39][10]  ( .D(n9880), .CK(CLK), .QN(n32068) );
  DFF_X1 \OUT2_reg[10]  ( .D(n7256), .CK(CLK), .Q(OUT2[10]), .QN(n16995) );
  DFF_X1 \OUT1_reg[10]  ( .D(n7320), .CK(CLK), .Q(OUT1[10]), .QN(n17059) );
  DFF_X1 \REGISTERS_reg[39][9]  ( .D(n9881), .CK(CLK), .QN(n32069) );
  DFF_X1 \OUT2_reg[9]  ( .D(n7257), .CK(CLK), .Q(OUT2[9]), .QN(n16996) );
  DFF_X1 \OUT1_reg[9]  ( .D(n7321), .CK(CLK), .Q(OUT1[9]), .QN(n17060) );
  DFF_X1 \REGISTERS_reg[39][8]  ( .D(n9882), .CK(CLK), .QN(n32070) );
  DFF_X1 \OUT2_reg[8]  ( .D(n7258), .CK(CLK), .Q(OUT2[8]), .QN(n16997) );
  DFF_X1 \OUT1_reg[8]  ( .D(n7322), .CK(CLK), .Q(OUT1[8]), .QN(n17061) );
  DFF_X1 \REGISTERS_reg[39][7]  ( .D(n9883), .CK(CLK), .QN(n32071) );
  DFF_X1 \OUT2_reg[7]  ( .D(n7259), .CK(CLK), .Q(OUT2[7]), .QN(n16998) );
  DFF_X1 \OUT1_reg[7]  ( .D(n7323), .CK(CLK), .Q(OUT1[7]), .QN(n17062) );
  DFF_X1 \REGISTERS_reg[39][6]  ( .D(n9884), .CK(CLK), .QN(n32072) );
  DFF_X1 \OUT2_reg[6]  ( .D(n7260), .CK(CLK), .Q(OUT2[6]), .QN(n16999) );
  DFF_X1 \OUT1_reg[6]  ( .D(n7324), .CK(CLK), .Q(OUT1[6]), .QN(n17063) );
  DFF_X1 \REGISTERS_reg[39][5]  ( .D(n9885), .CK(CLK), .QN(n32073) );
  DFF_X1 \OUT2_reg[5]  ( .D(n7261), .CK(CLK), .Q(OUT2[5]), .QN(n17000) );
  DFF_X1 \OUT1_reg[5]  ( .D(n7325), .CK(CLK), .Q(OUT1[5]), .QN(n17064) );
  DFF_X1 \REGISTERS_reg[39][4]  ( .D(n9886), .CK(CLK), .QN(n32074) );
  DFF_X1 \OUT2_reg[4]  ( .D(n7262), .CK(CLK), .Q(OUT2[4]), .QN(n17001) );
  DFF_X1 \OUT1_reg[4]  ( .D(n7326), .CK(CLK), .Q(OUT1[4]), .QN(n17065) );
  DFF_X1 \OUT2_reg[3]  ( .D(n7263), .CK(CLK), .Q(OUT2[3]), .QN(n17002) );
  DFF_X1 \OUT1_reg[3]  ( .D(n7327), .CK(CLK), .Q(OUT1[3]), .QN(n17066) );
  DFF_X1 \OUT2_reg[2]  ( .D(n7264), .CK(CLK), .Q(OUT2[2]), .QN(n17003) );
  DFF_X1 \OUT1_reg[2]  ( .D(n7328), .CK(CLK), .Q(OUT1[2]), .QN(n17067) );
  DFF_X1 \OUT2_reg[1]  ( .D(n7265), .CK(CLK), .Q(OUT2[1]), .QN(n17004) );
  DFF_X1 \OUT1_reg[1]  ( .D(n7329), .CK(CLK), .Q(OUT1[1]), .QN(n17068) );
  DFF_X1 \OUT2_reg[0]  ( .D(n7266), .CK(CLK), .Q(OUT2[0]), .QN(n17005) );
  DFF_X1 \OUT1_reg[0]  ( .D(n7330), .CK(CLK), .Q(OUT1[0]), .QN(n17069) );
  DFF_X1 \BUSout_reg[59]  ( .D(n7197), .CK(CLK), .Q(BUSout[59]), .QN(n16937)
         );
  DFF_X1 \BUSout_reg[58]  ( .D(n7196), .CK(CLK), .Q(BUSout[58]), .QN(n16936)
         );
  DFF_X1 \BUSout_reg[57]  ( .D(n7195), .CK(CLK), .Q(BUSout[57]), .QN(n16935)
         );
  DFF_X1 \BUSout_reg[56]  ( .D(n7194), .CK(CLK), .Q(BUSout[56]), .QN(n16934)
         );
  DFF_X1 \BUSout_reg[55]  ( .D(n7193), .CK(CLK), .Q(BUSout[55]), .QN(n16933)
         );
  DFF_X1 \BUSout_reg[54]  ( .D(n7192), .CK(CLK), .Q(BUSout[54]), .QN(n16932)
         );
  DFF_X1 \BUSout_reg[0]  ( .D(n7138), .CK(CLK), .Q(BUSout[0]), .QN(n16878) );
  FA_X1 \add_146/U1_1  ( .A(N659), .B(\i[1] ), .CI(n12791), .CO(
        \add_146/carry[2] ), .S(N811) );
  FA_X1 \add_146/U1_2  ( .A(N660), .B(\i[2] ), .CI(\add_146/carry[2] ), .CO(
        \add_146/carry[3] ), .S(N812) );
  FA_X1 \add_146/U1_3  ( .A(N661), .B(\i[3] ), .CI(\add_146/carry[3] ), .CO(
        \add_146/carry[4] ), .S(N813) );
  FA_X1 \r510/U1_1  ( .A(\U3/U195/Z_1 ), .B(ADD_RD2[1]), .CI(\r510/n3 ), .CO(
        \r510/carry[2] ), .S(N6395) );
  FA_X1 \r510/U1_2  ( .A(\U3/U195/Z_2 ), .B(ADD_RD2[2]), .CI(\r510/carry[2] ), 
        .CO(\r510/carry[3] ), .S(N6396) );
  FA_X1 \r510/U1_3  ( .A(\U3/U195/Z_3 ), .B(ADD_RD2[3]), .CI(\r510/carry[3] ), 
        .CO(\r510/carry[4] ), .S(N6397) );
  FA_X1 \r510/U1_4  ( .A(\U3/U195/Z_4 ), .B(ADD_RD2[4]), .CI(\r510/carry[4] ), 
        .CO(\r510/carry[5] ), .S(N6398) );
  FA_X1 \r504/U1_1  ( .A(\U3/U194/Z_1 ), .B(ADD_RD1[1]), .CI(\r504/n3 ), .CO(
        \r504/carry[2] ), .S(N6270) );
  FA_X1 \r504/U1_2  ( .A(\U3/U194/Z_2 ), .B(ADD_RD1[2]), .CI(\r504/carry[2] ), 
        .CO(\r504/carry[3] ), .S(N6271) );
  FA_X1 \r504/U1_3  ( .A(\U3/U194/Z_3 ), .B(ADD_RD1[3]), .CI(\r504/carry[3] ), 
        .CO(\r504/carry[4] ), .S(N6272) );
  FA_X1 \r504/U1_4  ( .A(\U3/U194/Z_4 ), .B(ADD_RD1[4]), .CI(\r504/carry[4] ), 
        .CO(\r504/carry[5] ), .S(N6273) );
  FA_X1 \r498/U1_1  ( .A(\U3/U193/Z_1 ), .B(ADD_WR[1]), .CI(\r498/n1 ), .CO(
        \r498/carry[2] ), .S(N929) );
  FA_X1 \r498/U1_2  ( .A(\U3/U193/Z_2 ), .B(ADD_WR[2]), .CI(\r498/carry[2] ), 
        .CO(\r498/carry[3] ), .S(N930) );
  FA_X1 \r498/U1_3  ( .A(\U3/U193/Z_3 ), .B(ADD_WR[3]), .CI(\r498/carry[3] ), 
        .CO(\r498/carry[4] ), .S(N931) );
  FA_X1 \r498/U1_4  ( .A(\U3/U193/Z_4 ), .B(ADD_WR[4]), .CI(\r498/carry[4] ), 
        .CO(\r498/carry[5] ), .S(N932) );
  FA_X1 \add_136/U1_1  ( .A(N659), .B(\i[1] ), .CI(n12791), .CO(
        \add_136/carry[2] ), .S(N688) );
  FA_X1 \add_136/U1_2  ( .A(N660), .B(\i[2] ), .CI(\add_136/carry[2] ), .CO(
        \add_136/carry[3] ), .S(N689) );
  FA_X1 \add_136/U1_3  ( .A(N661), .B(\i[3] ), .CI(\add_136/carry[3] ), .CO(
        \add_136/carry[4] ), .S(N690) );
  DFF_X1 \REGISTERS_reg[39][3]  ( .D(n9887), .CK(CLK), .QN(n32262) );
  DFF_X1 \REGISTERS_reg[39][2]  ( .D(n9888), .CK(CLK), .QN(n32263) );
  DFF_X1 \REGISTERS_reg[39][1]  ( .D(n9889), .CK(CLK), .QN(n32264) );
  DFF_X1 \REGISTERS_reg[39][0]  ( .D(n9890), .CK(CLK), .QN(n32265) );
  DFF_X1 \REGISTERS_reg[33][3]  ( .D(n9503), .CK(CLK), .QN(n32266) );
  DFF_X1 \REGISTERS_reg[33][2]  ( .D(n9504), .CK(CLK), .QN(n32267) );
  DFF_X1 \REGISTERS_reg[33][1]  ( .D(n9505), .CK(CLK), .QN(n32268) );
  DFF_X1 \REGISTERS_reg[33][0]  ( .D(n9506), .CK(CLK), .QN(n32269) );
  DFF_X1 \REGISTERS_reg[34][3]  ( .D(n9567), .CK(CLK), .QN(n32270) );
  DFF_X1 \REGISTERS_reg[34][2]  ( .D(n9568), .CK(CLK), .QN(n32271) );
  DFF_X1 \REGISTERS_reg[34][1]  ( .D(n9569), .CK(CLK), .QN(n32272) );
  DFF_X1 \REGISTERS_reg[34][0]  ( .D(n9570), .CK(CLK), .QN(n32273) );
  DFF_X1 \REGISTERS_reg[32][3]  ( .D(n9439), .CK(CLK), .QN(n32274) );
  DFF_X1 \REGISTERS_reg[32][2]  ( .D(n9440), .CK(CLK), .QN(n32275) );
  DFF_X1 \REGISTERS_reg[32][1]  ( .D(n9441), .CK(CLK), .QN(n32276) );
  DFF_X1 \REGISTERS_reg[32][0]  ( .D(n9442), .CK(CLK), .QN(n32277) );
  DFF_X1 \REGISTERS_reg[38][3]  ( .D(n9823), .CK(CLK), .QN(n32278) );
  DFF_X1 \REGISTERS_reg[38][2]  ( .D(n9824), .CK(CLK), .QN(n32279) );
  DFF_X1 \REGISTERS_reg[38][1]  ( .D(n9825), .CK(CLK), .QN(n32280) );
  DFF_X1 \REGISTERS_reg[38][0]  ( .D(n9826), .CK(CLK), .QN(n32281) );
  DFF_X1 \REGISTERS_reg[37][3]  ( .D(n9759), .CK(CLK), .QN(n32282) );
  DFF_X1 \REGISTERS_reg[37][2]  ( .D(n9760), .CK(CLK), .QN(n32283) );
  DFF_X1 \REGISTERS_reg[37][1]  ( .D(n9761), .CK(CLK), .QN(n32284) );
  DFF_X1 \REGISTERS_reg[37][0]  ( .D(n9762), .CK(CLK), .QN(n32285) );
  DFF_X1 \REGISTERS_reg[39][60]  ( .D(n9830), .CK(CLK), .QN(n32286) );
  DFF_X1 \REGISTERS_reg[39][58]  ( .D(n9832), .CK(CLK), .QN(n32287) );
  DFF_X1 \REGISTERS_reg[39][57]  ( .D(n9833), .CK(CLK), .QN(n32288) );
  DFF_X1 \REGISTERS_reg[39][56]  ( .D(n9834), .CK(CLK), .QN(n32289) );
  DFF_X1 \REGISTERS_reg[39][55]  ( .D(n9835), .CK(CLK), .QN(n32290) );
  DFF_X1 \REGISTERS_reg[39][54]  ( .D(n9836), .CK(CLK), .QN(n32291) );
  DFF_X1 \REGISTERS_reg[39][53]  ( .D(n9837), .CK(CLK), .QN(n32292) );
  DFF_X1 \REGISTERS_reg[39][52]  ( .D(n9838), .CK(CLK), .QN(n32293) );
  DFF_X1 \REGISTERS_reg[39][51]  ( .D(n9839), .CK(CLK), .QN(n32294) );
  DFF_X1 \REGISTERS_reg[39][50]  ( .D(n9840), .CK(CLK), .QN(n32295) );
  DFF_X1 \REGISTERS_reg[39][49]  ( .D(n9841), .CK(CLK), .QN(n32296) );
  DFF_X1 \REGISTERS_reg[39][48]  ( .D(n9842), .CK(CLK), .QN(n32297) );
  DFF_X1 \REGISTERS_reg[39][47]  ( .D(n9843), .CK(CLK), .QN(n32298) );
  DFF_X1 \REGISTERS_reg[39][46]  ( .D(n9844), .CK(CLK), .QN(n32299) );
  DFF_X1 \REGISTERS_reg[39][45]  ( .D(n9845), .CK(CLK), .QN(n32300) );
  DFF_X1 \REGISTERS_reg[39][44]  ( .D(n9846), .CK(CLK), .QN(n32301) );
  DFF_X1 \REGISTERS_reg[39][43]  ( .D(n9847), .CK(CLK), .QN(n32302) );
  DFF_X1 \REGISTERS_reg[39][42]  ( .D(n9848), .CK(CLK), .QN(n32303) );
  DFF_X1 \REGISTERS_reg[39][41]  ( .D(n9849), .CK(CLK), .QN(n32304) );
  DFF_X1 \REGISTERS_reg[39][40]  ( .D(n9850), .CK(CLK), .QN(n32305) );
  DFF_X1 \REGISTERS_reg[39][39]  ( .D(n9851), .CK(CLK), .QN(n32306) );
  DFF_X1 \REGISTERS_reg[39][38]  ( .D(n9852), .CK(CLK), .QN(n32307) );
  DFF_X1 \REGISTERS_reg[39][37]  ( .D(n9853), .CK(CLK), .QN(n32308) );
  DFF_X1 \REGISTERS_reg[39][36]  ( .D(n9854), .CK(CLK), .QN(n32309) );
  DFF_X1 \REGISTERS_reg[39][35]  ( .D(n9855), .CK(CLK), .QN(n32310) );
  DFF_X1 \REGISTERS_reg[39][34]  ( .D(n9856), .CK(CLK), .QN(n32311) );
  DFF_X1 \REGISTERS_reg[39][33]  ( .D(n9857), .CK(CLK), .QN(n32312) );
  DFF_X1 \REGISTERS_reg[39][32]  ( .D(n9858), .CK(CLK), .QN(n32313) );
  DFF_X1 \REGISTERS_reg[39][31]  ( .D(n9859), .CK(CLK), .QN(n32314) );
  DFF_X1 \REGISTERS_reg[39][30]  ( .D(n9860), .CK(CLK), .QN(n32315) );
  DFF_X1 \REGISTERS_reg[39][29]  ( .D(n9861), .CK(CLK), .QN(n32316) );
  DFF_X1 \REGISTERS_reg[39][28]  ( .D(n9862), .CK(CLK), .QN(n32317) );
  DFF_X1 \REGISTERS_reg[39][27]  ( .D(n9863), .CK(CLK), .QN(n32318) );
  DFF_X1 \REGISTERS_reg[39][26]  ( .D(n9864), .CK(CLK), .QN(n32319) );
  DFF_X1 \REGISTERS_reg[39][25]  ( .D(n9865), .CK(CLK), .QN(n32320) );
  DFF_X1 \REGISTERS_reg[39][24]  ( .D(n9866), .CK(CLK), .QN(n32321) );
  DFF_X1 \REGISTERS_reg[35][3]  ( .D(n9631), .CK(CLK), .Q(n30063), .QN(n39046)
         );
  DFF_X1 \REGISTERS_reg[35][2]  ( .D(n9632), .CK(CLK), .Q(n30064), .QN(n39045)
         );
  DFF_X1 \REGISTERS_reg[35][1]  ( .D(n9633), .CK(CLK), .Q(n30065), .QN(n39044)
         );
  DFF_X1 \REGISTERS_reg[35][0]  ( .D(n9634), .CK(CLK), .Q(n30066), .QN(n39043)
         );
  DFF_X1 \REGISTERS_reg[36][3]  ( .D(n9695), .CK(CLK), .Q(n30127), .QN(n38923)
         );
  DFF_X1 \REGISTERS_reg[36][2]  ( .D(n9696), .CK(CLK), .Q(n30128), .QN(n38922)
         );
  DFF_X1 \REGISTERS_reg[36][1]  ( .D(n9697), .CK(CLK), .Q(n30129), .QN(n38921)
         );
  DFF_X1 \REGISTERS_reg[36][0]  ( .D(n9698), .CK(CLK), .Q(n30130), .QN(n38920)
         );
  DFF_X1 \REGISTERS_reg[35][51]  ( .D(n9583), .CK(CLK), .Q(n30015), .QN(n39042) );
  DFF_X1 \REGISTERS_reg[35][50]  ( .D(n9584), .CK(CLK), .Q(n30016), .QN(n39041) );
  DFF_X1 \REGISTERS_reg[35][49]  ( .D(n9585), .CK(CLK), .Q(n30017), .QN(n39040) );
  DFF_X1 \REGISTERS_reg[35][48]  ( .D(n9586), .CK(CLK), .Q(n30018), .QN(n39039) );
  DFF_X1 \REGISTERS_reg[35][47]  ( .D(n9587), .CK(CLK), .Q(n30019), .QN(n39038) );
  DFF_X1 \REGISTERS_reg[35][46]  ( .D(n9588), .CK(CLK), .Q(n30020), .QN(n39037) );
  DFF_X1 \REGISTERS_reg[35][45]  ( .D(n9589), .CK(CLK), .Q(n30021), .QN(n39036) );
  DFF_X1 \REGISTERS_reg[35][44]  ( .D(n9590), .CK(CLK), .Q(n30022), .QN(n39035) );
  DFF_X1 \REGISTERS_reg[35][43]  ( .D(n9591), .CK(CLK), .Q(n30023), .QN(n39034) );
  DFF_X1 \REGISTERS_reg[35][42]  ( .D(n9592), .CK(CLK), .Q(n30024), .QN(n39033) );
  DFF_X1 \REGISTERS_reg[35][41]  ( .D(n9593), .CK(CLK), .Q(n30025), .QN(n39032) );
  DFF_X1 \REGISTERS_reg[35][40]  ( .D(n9594), .CK(CLK), .Q(n30026), .QN(n39031) );
  DFF_X1 \REGISTERS_reg[35][39]  ( .D(n9595), .CK(CLK), .Q(n30027), .QN(n39030) );
  DFF_X1 \REGISTERS_reg[35][38]  ( .D(n9596), .CK(CLK), .Q(n30028), .QN(n39029) );
  DFF_X1 \REGISTERS_reg[35][37]  ( .D(n9597), .CK(CLK), .Q(n30029), .QN(n39028) );
  DFF_X1 \REGISTERS_reg[35][36]  ( .D(n9598), .CK(CLK), .Q(n30030), .QN(n39027) );
  DFF_X1 \REGISTERS_reg[35][35]  ( .D(n9599), .CK(CLK), .Q(n30031), .QN(n39026) );
  DFF_X1 \REGISTERS_reg[35][34]  ( .D(n9600), .CK(CLK), .Q(n30032), .QN(n39025) );
  DFF_X1 \REGISTERS_reg[35][33]  ( .D(n9601), .CK(CLK), .Q(n30033), .QN(n39024) );
  DFF_X1 \REGISTERS_reg[35][32]  ( .D(n9602), .CK(CLK), .Q(n30034), .QN(n39023) );
  DFF_X1 \REGISTERS_reg[35][31]  ( .D(n9603), .CK(CLK), .Q(n30035), .QN(n39022) );
  DFF_X1 \REGISTERS_reg[35][30]  ( .D(n9604), .CK(CLK), .Q(n30036), .QN(n39021) );
  DFF_X1 \REGISTERS_reg[35][29]  ( .D(n9605), .CK(CLK), .Q(n30037), .QN(n39020) );
  DFF_X1 \REGISTERS_reg[35][28]  ( .D(n9606), .CK(CLK), .Q(n30038), .QN(n39019) );
  DFF_X1 \REGISTERS_reg[35][27]  ( .D(n9607), .CK(CLK), .Q(n30039), .QN(n39018) );
  DFF_X1 \REGISTERS_reg[35][26]  ( .D(n9608), .CK(CLK), .Q(n30040), .QN(n39017) );
  DFF_X1 \REGISTERS_reg[35][25]  ( .D(n9609), .CK(CLK), .Q(n30041), .QN(n39016) );
  DFF_X1 \REGISTERS_reg[35][24]  ( .D(n9610), .CK(CLK), .Q(n30042), .QN(n39015) );
  DFF_X1 \REGISTERS_reg[35][23]  ( .D(n9611), .CK(CLK), .Q(n30043), .QN(n39014) );
  DFF_X1 \REGISTERS_reg[35][22]  ( .D(n9612), .CK(CLK), .Q(n30044), .QN(n39013) );
  DFF_X1 \REGISTERS_reg[35][21]  ( .D(n9613), .CK(CLK), .Q(n30045), .QN(n39012) );
  DFF_X1 \REGISTERS_reg[35][20]  ( .D(n9614), .CK(CLK), .Q(n30046), .QN(n39011) );
  DFF_X1 \REGISTERS_reg[35][19]  ( .D(n9615), .CK(CLK), .Q(n30047), .QN(n39010) );
  DFF_X1 \REGISTERS_reg[35][18]  ( .D(n9616), .CK(CLK), .Q(n30048), .QN(n39009) );
  DFF_X1 \REGISTERS_reg[35][17]  ( .D(n9617), .CK(CLK), .Q(n30049), .QN(n39008) );
  DFF_X1 \REGISTERS_reg[35][16]  ( .D(n9618), .CK(CLK), .Q(n30050), .QN(n39007) );
  DFF_X1 \REGISTERS_reg[35][15]  ( .D(n9619), .CK(CLK), .Q(n30051), .QN(n39006) );
  DFF_X1 \REGISTERS_reg[35][14]  ( .D(n9620), .CK(CLK), .Q(n30052), .QN(n39005) );
  DFF_X1 \REGISTERS_reg[35][13]  ( .D(n9621), .CK(CLK), .Q(n30053), .QN(n39004) );
  DFF_X1 \REGISTERS_reg[35][12]  ( .D(n9622), .CK(CLK), .Q(n30054), .QN(n39003) );
  DFF_X1 \REGISTERS_reg[35][11]  ( .D(n9623), .CK(CLK), .Q(n30055), .QN(n39002) );
  DFF_X1 \REGISTERS_reg[35][10]  ( .D(n9624), .CK(CLK), .Q(n30056), .QN(n39001) );
  DFF_X1 \REGISTERS_reg[35][9]  ( .D(n9625), .CK(CLK), .Q(n30057), .QN(n39000)
         );
  DFF_X1 \REGISTERS_reg[35][8]  ( .D(n9626), .CK(CLK), .Q(n30058), .QN(n38999)
         );
  DFF_X1 \REGISTERS_reg[35][7]  ( .D(n9627), .CK(CLK), .Q(n30059), .QN(n38998)
         );
  DFF_X1 \REGISTERS_reg[35][6]  ( .D(n9628), .CK(CLK), .Q(n30060), .QN(n38997)
         );
  DFF_X1 \REGISTERS_reg[35][5]  ( .D(n9629), .CK(CLK), .Q(n30061), .QN(n38996)
         );
  DFF_X1 \REGISTERS_reg[35][4]  ( .D(n9630), .CK(CLK), .Q(n30062), .QN(n38995)
         );
  DFF_X1 \REGISTERS_reg[35][63]  ( .D(n9571), .CK(CLK), .Q(n30003), .QN(n38926) );
  DFF_X1 \REGISTERS_reg[35][62]  ( .D(n9572), .CK(CLK), .Q(n30004), .QN(n38925) );
  DFF_X1 \REGISTERS_reg[35][61]  ( .D(n9573), .CK(CLK), .Q(n30005), .QN(n38924) );
  DFF_X1 \REGISTERS_reg[35][60]  ( .D(n9574), .CK(CLK), .Q(n30006), .QN(n38994) );
  DFF_X1 \REGISTERS_reg[35][59]  ( .D(n9575), .CK(CLK), .Q(n30007), .QN(n32384) );
  DFF_X1 \REGISTERS_reg[35][58]  ( .D(n9576), .CK(CLK), .Q(n30008), .QN(n38993) );
  DFF_X1 \REGISTERS_reg[35][57]  ( .D(n9577), .CK(CLK), .Q(n30009), .QN(n38992) );
  DFF_X1 \REGISTERS_reg[35][56]  ( .D(n9578), .CK(CLK), .Q(n30010), .QN(n38991) );
  DFF_X1 \REGISTERS_reg[35][55]  ( .D(n9579), .CK(CLK), .Q(n30011), .QN(n38990) );
  DFF_X1 \REGISTERS_reg[35][54]  ( .D(n9580), .CK(CLK), .Q(n30012), .QN(n38989) );
  DFF_X1 \REGISTERS_reg[35][53]  ( .D(n9581), .CK(CLK), .Q(n30013), .QN(n38988) );
  DFF_X1 \REGISTERS_reg[35][52]  ( .D(n9582), .CK(CLK), .Q(n30014), .QN(n38987) );
  DFF_X1 \REGISTERS_reg[36][51]  ( .D(n9647), .CK(CLK), .Q(n30079), .QN(n38919) );
  DFF_X1 \REGISTERS_reg[36][50]  ( .D(n9648), .CK(CLK), .Q(n30080), .QN(n38918) );
  DFF_X1 \REGISTERS_reg[36][49]  ( .D(n9649), .CK(CLK), .Q(n30081), .QN(n38917) );
  DFF_X1 \REGISTERS_reg[36][48]  ( .D(n9650), .CK(CLK), .Q(n30082), .QN(n38916) );
  DFF_X1 \REGISTERS_reg[36][47]  ( .D(n9651), .CK(CLK), .Q(n30083), .QN(n38915) );
  DFF_X1 \REGISTERS_reg[36][46]  ( .D(n9652), .CK(CLK), .Q(n30084), .QN(n38914) );
  DFF_X1 \REGISTERS_reg[36][45]  ( .D(n9653), .CK(CLK), .Q(n30085), .QN(n38913) );
  DFF_X1 \REGISTERS_reg[36][44]  ( .D(n9654), .CK(CLK), .Q(n30086), .QN(n38912) );
  DFF_X1 \REGISTERS_reg[36][43]  ( .D(n9655), .CK(CLK), .Q(n30087), .QN(n38911) );
  DFF_X1 \REGISTERS_reg[36][42]  ( .D(n9656), .CK(CLK), .Q(n30088), .QN(n38910) );
  DFF_X1 \REGISTERS_reg[36][41]  ( .D(n9657), .CK(CLK), .Q(n30089), .QN(n38909) );
  DFF_X1 \REGISTERS_reg[36][40]  ( .D(n9658), .CK(CLK), .Q(n30090), .QN(n38908) );
  DFF_X1 \REGISTERS_reg[36][39]  ( .D(n9659), .CK(CLK), .Q(n30091), .QN(n38907) );
  DFF_X1 \REGISTERS_reg[36][38]  ( .D(n9660), .CK(CLK), .Q(n30092), .QN(n38906) );
  DFF_X1 \REGISTERS_reg[36][37]  ( .D(n9661), .CK(CLK), .Q(n30093), .QN(n38905) );
  DFF_X1 \REGISTERS_reg[36][36]  ( .D(n9662), .CK(CLK), .Q(n30094), .QN(n38904) );
  DFF_X1 \REGISTERS_reg[36][35]  ( .D(n9663), .CK(CLK), .Q(n30095), .QN(n38903) );
  DFF_X1 \REGISTERS_reg[36][34]  ( .D(n9664), .CK(CLK), .Q(n30096), .QN(n38902) );
  DFF_X1 \REGISTERS_reg[36][33]  ( .D(n9665), .CK(CLK), .Q(n30097), .QN(n38901) );
  DFF_X1 \REGISTERS_reg[36][32]  ( .D(n9666), .CK(CLK), .Q(n30098), .QN(n38900) );
  DFF_X1 \REGISTERS_reg[36][31]  ( .D(n9667), .CK(CLK), .Q(n30099), .QN(n38899) );
  DFF_X1 \REGISTERS_reg[36][30]  ( .D(n9668), .CK(CLK), .Q(n30100), .QN(n38898) );
  DFF_X1 \REGISTERS_reg[36][29]  ( .D(n9669), .CK(CLK), .Q(n30101), .QN(n38897) );
  DFF_X1 \REGISTERS_reg[36][28]  ( .D(n9670), .CK(CLK), .Q(n30102), .QN(n38896) );
  DFF_X1 \REGISTERS_reg[36][27]  ( .D(n9671), .CK(CLK), .Q(n30103), .QN(n38895) );
  DFF_X1 \REGISTERS_reg[36][26]  ( .D(n9672), .CK(CLK), .Q(n30104), .QN(n38894) );
  DFF_X1 \REGISTERS_reg[36][25]  ( .D(n9673), .CK(CLK), .Q(n30105), .QN(n38893) );
  DFF_X1 \REGISTERS_reg[36][24]  ( .D(n9674), .CK(CLK), .Q(n30106), .QN(n38892) );
  DFF_X1 \REGISTERS_reg[36][23]  ( .D(n9675), .CK(CLK), .Q(n30107), .QN(n38891) );
  DFF_X1 \REGISTERS_reg[36][22]  ( .D(n9676), .CK(CLK), .Q(n30108), .QN(n38890) );
  DFF_X1 \REGISTERS_reg[36][21]  ( .D(n9677), .CK(CLK), .Q(n30109), .QN(n38889) );
  DFF_X1 \REGISTERS_reg[36][20]  ( .D(n9678), .CK(CLK), .Q(n30110), .QN(n38888) );
  DFF_X1 \REGISTERS_reg[36][19]  ( .D(n9679), .CK(CLK), .Q(n30111), .QN(n38887) );
  DFF_X1 \REGISTERS_reg[36][18]  ( .D(n9680), .CK(CLK), .Q(n30112), .QN(n38886) );
  DFF_X1 \REGISTERS_reg[36][17]  ( .D(n9681), .CK(CLK), .Q(n30113), .QN(n38885) );
  DFF_X1 \REGISTERS_reg[36][16]  ( .D(n9682), .CK(CLK), .Q(n30114), .QN(n38884) );
  DFF_X1 \REGISTERS_reg[36][15]  ( .D(n9683), .CK(CLK), .Q(n30115), .QN(n38883) );
  DFF_X1 \REGISTERS_reg[36][14]  ( .D(n9684), .CK(CLK), .Q(n30116), .QN(n38882) );
  DFF_X1 \REGISTERS_reg[36][13]  ( .D(n9685), .CK(CLK), .Q(n30117), .QN(n38881) );
  DFF_X1 \REGISTERS_reg[36][12]  ( .D(n9686), .CK(CLK), .Q(n30118), .QN(n38880) );
  DFF_X1 \REGISTERS_reg[36][11]  ( .D(n9687), .CK(CLK), .Q(n30119), .QN(n38879) );
  DFF_X1 \REGISTERS_reg[36][10]  ( .D(n9688), .CK(CLK), .Q(n30120), .QN(n38878) );
  DFF_X1 \REGISTERS_reg[36][9]  ( .D(n9689), .CK(CLK), .Q(n30121), .QN(n38877)
         );
  DFF_X1 \REGISTERS_reg[36][8]  ( .D(n9690), .CK(CLK), .Q(n30122), .QN(n38876)
         );
  DFF_X1 \REGISTERS_reg[36][7]  ( .D(n9691), .CK(CLK), .Q(n30123), .QN(n38875)
         );
  DFF_X1 \REGISTERS_reg[36][6]  ( .D(n9692), .CK(CLK), .Q(n30124), .QN(n38874)
         );
  DFF_X1 \REGISTERS_reg[36][5]  ( .D(n9693), .CK(CLK), .Q(n30125), .QN(n38873)
         );
  DFF_X1 \REGISTERS_reg[36][4]  ( .D(n9694), .CK(CLK), .Q(n30126), .QN(n38872)
         );
  DFF_X1 \REGISTERS_reg[36][63]  ( .D(n9635), .CK(CLK), .Q(n30067), .QN(n38793) );
  DFF_X1 \REGISTERS_reg[36][62]  ( .D(n9636), .CK(CLK), .Q(n30068), .QN(n38792) );
  DFF_X1 \REGISTERS_reg[36][61]  ( .D(n9637), .CK(CLK), .Q(n30069), .QN(n38791) );
  DFF_X1 \REGISTERS_reg[36][60]  ( .D(n9638), .CK(CLK), .Q(n30070), .QN(n38871) );
  DFF_X1 \REGISTERS_reg[36][59]  ( .D(n9639), .CK(CLK), .Q(n30071), .QN(n32444) );
  DFF_X1 \REGISTERS_reg[36][58]  ( .D(n9640), .CK(CLK), .Q(n30072), .QN(n38870) );
  DFF_X1 \REGISTERS_reg[36][57]  ( .D(n9641), .CK(CLK), .Q(n30073), .QN(n38869) );
  DFF_X1 \REGISTERS_reg[36][56]  ( .D(n9642), .CK(CLK), .Q(n30074), .QN(n38868) );
  DFF_X1 \REGISTERS_reg[36][55]  ( .D(n9643), .CK(CLK), .Q(n30075), .QN(n38867) );
  DFF_X1 \REGISTERS_reg[36][54]  ( .D(n9644), .CK(CLK), .Q(n30076), .QN(n38866) );
  DFF_X1 \REGISTERS_reg[36][53]  ( .D(n9645), .CK(CLK), .Q(n30077), .QN(n38865) );
  DFF_X1 \REGISTERS_reg[36][52]  ( .D(n9646), .CK(CLK), .Q(n30078), .QN(n38864) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n8415), .CK(CLK), .Q(n28847), .QN(n38863)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n8416), .CK(CLK), .Q(n28848), .QN(n38862)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n8417), .CK(CLK), .Q(n28849), .QN(n38861)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n8418), .CK(CLK), .Q(n28850), .QN(n38860)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n9055), .CK(CLK), .Q(n29487), .QN(n32460)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n9056), .CK(CLK), .Q(n29488), .QN(n32461)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n9057), .CK(CLK), .Q(n29489), .QN(n32462)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n9058), .CK(CLK), .Q(n29490), .QN(n32463)
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n8991), .CK(CLK), .Q(n29423), .QN(n32464)
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n8992), .CK(CLK), .Q(n29424), .QN(n32465)
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n8993), .CK(CLK), .Q(n29425), .QN(n32466)
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n8994), .CK(CLK), .Q(n29426), .QN(n32467)
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n8735), .CK(CLK), .Q(n29167), .QN(n32476)
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n8736), .CK(CLK), .Q(n29168), .QN(n32477)
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n8737), .CK(CLK), .Q(n29169), .QN(n32478)
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n8738), .CK(CLK), .Q(n29170), .QN(n32479)
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n8671), .CK(CLK), .Q(n29103), .QN(n32480)
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n8672), .CK(CLK), .Q(n29104), .QN(n32481)
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n8673), .CK(CLK), .Q(n29105), .QN(n32482)
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n8674), .CK(CLK), .Q(n29106), .QN(n32483)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n9311), .CK(CLK), .Q(n29743), .QN(n38986)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n9312), .CK(CLK), .Q(n29744), .QN(n38985)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n9313), .CK(CLK), .Q(n29745), .QN(n38984)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n9314), .CK(CLK), .Q(n29746), .QN(n38983)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n9375), .CK(CLK), .Q(n29807), .QN(n38859)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n9376), .CK(CLK), .Q(n29808), .QN(n38858)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n9377), .CK(CLK), .Q(n29809), .QN(n38857)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n9378), .CK(CLK), .Q(n29810), .QN(n38856)
         );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n8409), .CK(CLK), .Q(n28841), .QN(n38855)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n8410), .CK(CLK), .Q(n28842), .QN(n38854)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n8411), .CK(CLK), .Q(n28843), .QN(n38853)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n8413), .CK(CLK), .Q(n28845), .QN(n38852)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n8414), .CK(CLK), .Q(n28846), .QN(n38851)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n8412), .CK(CLK), .Q(n28844), .QN(n38850)
         );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7407), .CK(CLK), .Q(n27956), .QN(n32547)
         );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7408), .CK(CLK), .Q(n27957), .QN(n32548)
         );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7409), .CK(CLK), .Q(n27958), .QN(n32549)
         );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7410), .CK(CLK), .Q(n27959), .QN(n32550)
         );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7411), .CK(CLK), .Q(n27960), .QN(n32551)
         );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7412), .CK(CLK), .Q(n27961), .QN(n32552)
         );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7413), .CK(CLK), .Q(n27962), .QN(n32553)
         );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7414), .CK(CLK), .Q(n27963), .QN(n32554)
         );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7415), .CK(CLK), .Q(n27964), .QN(n32555)
         );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7416), .CK(CLK), .Q(n27965), .QN(n32556)
         );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7417), .CK(CLK), .Q(n27966), .QN(n32557)
         );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7418), .CK(CLK), .Q(n27967), .QN(n32558)
         );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7419), .CK(CLK), .Q(n27968), .QN(n32559)
         );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7420), .CK(CLK), .Q(n27969), .QN(n32560)
         );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7421), .CK(CLK), .Q(n27970), .QN(n32561)
         );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7422), .CK(CLK), .Q(n27971), .QN(n32562)
         );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7423), .CK(CLK), .Q(n27972), .QN(n32563)
         );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7424), .CK(CLK), .Q(n27973), .QN(n32564)
         );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7425), .CK(CLK), .Q(n27974), .QN(n32565)
         );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7426), .CK(CLK), .Q(n27975), .QN(n32566)
         );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7427), .CK(CLK), .Q(n27976), .QN(n32567)
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7428), .CK(CLK), .Q(n27977), .QN(n32568)
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7429), .CK(CLK), .Q(n27978), .QN(n32569)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7430), .CK(CLK), .Q(n27979), .QN(n32570)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7431), .CK(CLK), .Q(n27980), .QN(n32571)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7432), .CK(CLK), .Q(n27981), .QN(n32572)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7433), .CK(CLK), .Q(n27982), .QN(n32573)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7434), .CK(CLK), .Q(n27983), .QN(n32574)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7435), .CK(CLK), .Q(n27984), .QN(n32575)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7436), .CK(CLK), .Q(n27985), .QN(n32576)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7437), .CK(CLK), .Q(n27986), .QN(n32577)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7438), .CK(CLK), .Q(n27987), .QN(n32578)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n7439), .CK(CLK), .Q(n27988), .QN(n32579)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n7440), .CK(CLK), .Q(n27989), .QN(n32580)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n7441), .CK(CLK), .Q(n27990), .QN(n32581)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n7442), .CK(CLK), .Q(n27991), .QN(n32582)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n7443), .CK(CLK), .Q(n27992), .QN(n32583)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n7444), .CK(CLK), .Q(n27993), .QN(n32584)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n7445), .CK(CLK), .Q(n27994), .QN(n32585)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n7446), .CK(CLK), .Q(n27995), .QN(n32586)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n7447), .CK(CLK), .Q(n27996), .QN(n32587)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n7448), .CK(CLK), .Q(n27997), .QN(n32588)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n7449), .CK(CLK), .Q(n27998), .QN(n32589)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n7450), .CK(CLK), .Q(n27999), .QN(n32590)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n7451), .CK(CLK), .Q(n28000), .QN(n32591)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n7452), .CK(CLK), .Q(n28001), .QN(n32592)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n7453), .CK(CLK), .Q(n28002), .QN(n32593)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n7454), .CK(CLK), .Q(n28003), .QN(n32594)
         );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n9007), .CK(CLK), .Q(n29439), .QN(n32595) );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n9008), .CK(CLK), .Q(n29440), .QN(n32596) );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n9009), .CK(CLK), .Q(n29441), .QN(n32597) );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n9010), .CK(CLK), .Q(n29442), .QN(n32598) );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n9011), .CK(CLK), .Q(n29443), .QN(n32599) );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n9012), .CK(CLK), .Q(n29444), .QN(n32600) );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n9013), .CK(CLK), .Q(n29445), .QN(n32601) );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n9014), .CK(CLK), .Q(n29446), .QN(n32602) );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n9015), .CK(CLK), .Q(n29447), .QN(n32603) );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n9016), .CK(CLK), .Q(n29448), .QN(n32604) );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n9017), .CK(CLK), .Q(n29449), .QN(n32605) );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n9018), .CK(CLK), .Q(n29450), .QN(n32606) );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n9019), .CK(CLK), .Q(n29451), .QN(n32607) );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n9020), .CK(CLK), .Q(n29452), .QN(n32608) );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n9021), .CK(CLK), .Q(n29453), .QN(n32609) );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n9022), .CK(CLK), .Q(n29454), .QN(n32610) );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n9023), .CK(CLK), .Q(n29455), .QN(n32611) );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n9024), .CK(CLK), .Q(n29456), .QN(n32612) );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n9025), .CK(CLK), .Q(n29457), .QN(n32613) );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n9026), .CK(CLK), .Q(n29458), .QN(n32614) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n9027), .CK(CLK), .Q(n29459), .QN(n32615) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n9028), .CK(CLK), .Q(n29460), .QN(n32616) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n9029), .CK(CLK), .Q(n29461), .QN(n32617) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n9030), .CK(CLK), .Q(n29462), .QN(n32618) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n9031), .CK(CLK), .Q(n29463), .QN(n32619) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n9032), .CK(CLK), .Q(n29464), .QN(n32620) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n9033), .CK(CLK), .Q(n29465), .QN(n32621) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n9034), .CK(CLK), .Q(n29466), .QN(n32622) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n9035), .CK(CLK), .Q(n29467), .QN(n32623) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n9036), .CK(CLK), .Q(n29468), .QN(n32624) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n9037), .CK(CLK), .Q(n29469), .QN(n32625) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n9038), .CK(CLK), .Q(n29470), .QN(n32626) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n9039), .CK(CLK), .Q(n29471), .QN(n32627) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n9040), .CK(CLK), .Q(n29472), .QN(n32628) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n9041), .CK(CLK), .Q(n29473), .QN(n32629) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n9042), .CK(CLK), .Q(n29474), .QN(n32630) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n9043), .CK(CLK), .Q(n29475), .QN(n32631) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n9044), .CK(CLK), .Q(n29476), .QN(n32632) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n9045), .CK(CLK), .Q(n29477), .QN(n32633) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n9046), .CK(CLK), .Q(n29478), .QN(n32634) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n9047), .CK(CLK), .Q(n29479), .QN(n32635) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n9048), .CK(CLK), .Q(n29480), .QN(n32636) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n9049), .CK(CLK), .Q(n29481), .QN(n32637)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n9050), .CK(CLK), .Q(n29482), .QN(n32638)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n9051), .CK(CLK), .Q(n29483), .QN(n32639)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n9052), .CK(CLK), .Q(n29484), .QN(n32640)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n9053), .CK(CLK), .Q(n29485), .QN(n32641)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n9054), .CK(CLK), .Q(n29486), .QN(n32642)
         );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n8943), .CK(CLK), .Q(n29375), .QN(n32643) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n8944), .CK(CLK), .Q(n29376), .QN(n32644) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n8945), .CK(CLK), .Q(n29377), .QN(n32645) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n8946), .CK(CLK), .Q(n29378), .QN(n32646) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n8947), .CK(CLK), .Q(n29379), .QN(n32647) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n8948), .CK(CLK), .Q(n29380), .QN(n32648) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n8949), .CK(CLK), .Q(n29381), .QN(n32649) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n8950), .CK(CLK), .Q(n29382), .QN(n32650) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n8951), .CK(CLK), .Q(n29383), .QN(n32651) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n8952), .CK(CLK), .Q(n29384), .QN(n32652) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n8953), .CK(CLK), .Q(n29385), .QN(n32653) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n8954), .CK(CLK), .Q(n29386), .QN(n32654) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n8955), .CK(CLK), .Q(n29387), .QN(n32655) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n8956), .CK(CLK), .Q(n29388), .QN(n32656) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n8957), .CK(CLK), .Q(n29389), .QN(n32657) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n8958), .CK(CLK), .Q(n29390), .QN(n32658) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n8959), .CK(CLK), .Q(n29391), .QN(n32659) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n8960), .CK(CLK), .Q(n29392), .QN(n32660) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n8961), .CK(CLK), .Q(n29393), .QN(n32661) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n8962), .CK(CLK), .Q(n29394), .QN(n32662) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n8963), .CK(CLK), .Q(n29395), .QN(n32663) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n8964), .CK(CLK), .Q(n29396), .QN(n32664) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n8965), .CK(CLK), .Q(n29397), .QN(n32665) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n8966), .CK(CLK), .Q(n29398), .QN(n32666) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n8967), .CK(CLK), .Q(n29399), .QN(n32667) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n8968), .CK(CLK), .Q(n29400), .QN(n32668) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n8969), .CK(CLK), .Q(n29401), .QN(n32669) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n8970), .CK(CLK), .Q(n29402), .QN(n32670) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n8971), .CK(CLK), .Q(n29403), .QN(n32671) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n8972), .CK(CLK), .Q(n29404), .QN(n32672) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n8973), .CK(CLK), .Q(n29405), .QN(n32673) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n8974), .CK(CLK), .Q(n29406), .QN(n32674) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n8975), .CK(CLK), .Q(n29407), .QN(n32675) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n8976), .CK(CLK), .Q(n29408), .QN(n32676) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n8977), .CK(CLK), .Q(n29409), .QN(n32677) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n8978), .CK(CLK), .Q(n29410), .QN(n32678) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n8979), .CK(CLK), .Q(n29411), .QN(n32679) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n8980), .CK(CLK), .Q(n29412), .QN(n32680) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n8981), .CK(CLK), .Q(n29413), .QN(n32681) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n8982), .CK(CLK), .Q(n29414), .QN(n32682) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n8983), .CK(CLK), .Q(n29415), .QN(n32683) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n8984), .CK(CLK), .Q(n29416), .QN(n32684) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n8985), .CK(CLK), .Q(n29417), .QN(n32685)
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n8986), .CK(CLK), .Q(n29418), .QN(n32686)
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n8987), .CK(CLK), .Q(n29419), .QN(n32687)
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n8988), .CK(CLK), .Q(n29420), .QN(n32688)
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n8989), .CK(CLK), .Q(n29421), .QN(n32689)
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n8990), .CK(CLK), .Q(n29422), .QN(n32690)
         );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n7395), .CK(CLK), .Q(n27944), .QN(n32691)
         );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n7396), .CK(CLK), .Q(n27945), .QN(n32692)
         );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7397), .CK(CLK), .Q(n27946), .QN(n32693)
         );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7398), .CK(CLK), .Q(n27947), .QN(n32694)
         );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7399), .CK(CLK), .Q(n27948), .QN(n32695)
         );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7400), .CK(CLK), .Q(n27949), .QN(n32696)
         );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7401), .CK(CLK), .Q(n27950), .QN(n32697)
         );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7402), .CK(CLK), .Q(n27951), .QN(n32698)
         );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7403), .CK(CLK), .Q(n27952), .QN(n32699)
         );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7404), .CK(CLK), .Q(n27953), .QN(n32700)
         );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7405), .CK(CLK), .Q(n27954), .QN(n32701)
         );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7406), .CK(CLK), .Q(n27955), .QN(n32702)
         );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n8995), .CK(CLK), .Q(n29427), .QN(n32703) );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n8996), .CK(CLK), .Q(n29428), .QN(n32704) );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n8997), .CK(CLK), .Q(n29429), .QN(n32705) );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n8998), .CK(CLK), .Q(n29430), .QN(n32706) );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n8999), .CK(CLK), .Q(n29431), .QN(n32707) );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n9000), .CK(CLK), .Q(n29432), .QN(n32708) );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n9001), .CK(CLK), .Q(n29433), .QN(n32709) );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n9002), .CK(CLK), .Q(n29434), .QN(n32710) );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n9003), .CK(CLK), .Q(n29435), .QN(n32711) );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n9004), .CK(CLK), .Q(n29436), .QN(n32712) );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n9005), .CK(CLK), .Q(n29437), .QN(n32713) );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n9006), .CK(CLK), .Q(n29438), .QN(n32714) );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n8931), .CK(CLK), .Q(n29363), .QN(n32715) );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n8932), .CK(CLK), .Q(n29364), .QN(n32716) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n8933), .CK(CLK), .Q(n29365), .QN(n32717) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n8934), .CK(CLK), .Q(n29366), .QN(n32718) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n8935), .CK(CLK), .Q(n29367), .QN(n32719) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n8936), .CK(CLK), .Q(n29368), .QN(n32720) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n8937), .CK(CLK), .Q(n29369), .QN(n32721) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n8938), .CK(CLK), .Q(n29370), .QN(n32722) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n8939), .CK(CLK), .Q(n29371), .QN(n32723) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n8940), .CK(CLK), .Q(n29372), .QN(n32724) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n8941), .CK(CLK), .Q(n29373), .QN(n32725) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n8942), .CK(CLK), .Q(n29374), .QN(n32726) );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n8687), .CK(CLK), .Q(n29119), .QN(n32847) );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n8688), .CK(CLK), .Q(n29120), .QN(n32848) );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n8689), .CK(CLK), .Q(n29121), .QN(n32849) );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n8690), .CK(CLK), .Q(n29122), .QN(n32850) );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n8691), .CK(CLK), .Q(n29123), .QN(n32851) );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n8692), .CK(CLK), .Q(n29124), .QN(n32852) );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n8693), .CK(CLK), .Q(n29125), .QN(n32853) );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n8694), .CK(CLK), .Q(n29126), .QN(n32854) );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n8695), .CK(CLK), .Q(n29127), .QN(n32855) );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n8696), .CK(CLK), .Q(n29128), .QN(n32856) );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n8697), .CK(CLK), .Q(n29129), .QN(n32857) );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n8698), .CK(CLK), .Q(n29130), .QN(n32858) );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n8699), .CK(CLK), .Q(n29131), .QN(n32859) );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n8700), .CK(CLK), .Q(n29132), .QN(n32860) );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n8701), .CK(CLK), .Q(n29133), .QN(n32861) );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n8702), .CK(CLK), .Q(n29134), .QN(n32862) );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n8703), .CK(CLK), .Q(n29135), .QN(n32863) );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n8704), .CK(CLK), .Q(n29136), .QN(n32864) );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n8705), .CK(CLK), .Q(n29137), .QN(n32865) );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n8706), .CK(CLK), .Q(n29138), .QN(n32866) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n8707), .CK(CLK), .Q(n29139), .QN(n32867) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n8708), .CK(CLK), .Q(n29140), .QN(n32868) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n8709), .CK(CLK), .Q(n29141), .QN(n32869) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n8710), .CK(CLK), .Q(n29142), .QN(n32870) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n8711), .CK(CLK), .Q(n29143), .QN(n32871) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n8712), .CK(CLK), .Q(n29144), .QN(n32872) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n8713), .CK(CLK), .Q(n29145), .QN(n32873) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n8714), .CK(CLK), .Q(n29146), .QN(n32874) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n8715), .CK(CLK), .Q(n29147), .QN(n32875) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n8716), .CK(CLK), .Q(n29148), .QN(n32876) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n8717), .CK(CLK), .Q(n29149), .QN(n32877) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n8718), .CK(CLK), .Q(n29150), .QN(n32878) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n8719), .CK(CLK), .Q(n29151), .QN(n32879) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n8720), .CK(CLK), .Q(n29152), .QN(n32880) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n8721), .CK(CLK), .Q(n29153), .QN(n32881) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n8722), .CK(CLK), .Q(n29154), .QN(n32882) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n8723), .CK(CLK), .Q(n29155), .QN(n32883) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n8724), .CK(CLK), .Q(n29156), .QN(n32884) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n8725), .CK(CLK), .Q(n29157), .QN(n32885) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n8726), .CK(CLK), .Q(n29158), .QN(n32886) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n8727), .CK(CLK), .Q(n29159), .QN(n32887) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n8728), .CK(CLK), .Q(n29160), .QN(n32888) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n8729), .CK(CLK), .Q(n29161), .QN(n32889)
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n8730), .CK(CLK), .Q(n29162), .QN(n32890)
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n8731), .CK(CLK), .Q(n29163), .QN(n32891)
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n8732), .CK(CLK), .Q(n29164), .QN(n32892)
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n8733), .CK(CLK), .Q(n29165), .QN(n32893)
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n8734), .CK(CLK), .Q(n29166), .QN(n32894)
         );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n8623), .CK(CLK), .Q(n29055), .QN(n32895) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n8624), .CK(CLK), .Q(n29056), .QN(n32896) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n8625), .CK(CLK), .Q(n29057), .QN(n32897) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n8626), .CK(CLK), .Q(n29058), .QN(n32898) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n8627), .CK(CLK), .Q(n29059), .QN(n32899) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n8628), .CK(CLK), .Q(n29060), .QN(n32900) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n8629), .CK(CLK), .Q(n29061), .QN(n32901) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n8630), .CK(CLK), .Q(n29062), .QN(n32902) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n8631), .CK(CLK), .Q(n29063), .QN(n32903) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n8632), .CK(CLK), .Q(n29064), .QN(n32904) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n8633), .CK(CLK), .Q(n29065), .QN(n32905) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n8634), .CK(CLK), .Q(n29066), .QN(n32906) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n8635), .CK(CLK), .Q(n29067), .QN(n32907) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n8636), .CK(CLK), .Q(n29068), .QN(n32908) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n8637), .CK(CLK), .Q(n29069), .QN(n32909) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n8638), .CK(CLK), .Q(n29070), .QN(n32910) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n8639), .CK(CLK), .Q(n29071), .QN(n32911) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n8640), .CK(CLK), .Q(n29072), .QN(n32912) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n8641), .CK(CLK), .Q(n29073), .QN(n32913) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n8642), .CK(CLK), .Q(n29074), .QN(n32914) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n8643), .CK(CLK), .Q(n29075), .QN(n32915) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n8644), .CK(CLK), .Q(n29076), .QN(n32916) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n8645), .CK(CLK), .Q(n29077), .QN(n32917) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n8646), .CK(CLK), .Q(n29078), .QN(n32918) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n8647), .CK(CLK), .Q(n29079), .QN(n32919) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n8648), .CK(CLK), .Q(n29080), .QN(n32920) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n8649), .CK(CLK), .Q(n29081), .QN(n32921) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n8650), .CK(CLK), .Q(n29082), .QN(n32922) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n8651), .CK(CLK), .Q(n29083), .QN(n32923) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n8652), .CK(CLK), .Q(n29084), .QN(n32924) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n8653), .CK(CLK), .Q(n29085), .QN(n32925) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n8654), .CK(CLK), .Q(n29086), .QN(n32926) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n8655), .CK(CLK), .Q(n29087), .QN(n32927) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n8656), .CK(CLK), .Q(n29088), .QN(n32928) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n8657), .CK(CLK), .Q(n29089), .QN(n32929) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n8658), .CK(CLK), .Q(n29090), .QN(n32930) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n8659), .CK(CLK), .Q(n29091), .QN(n32931) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n8660), .CK(CLK), .Q(n29092), .QN(n32932) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n8661), .CK(CLK), .Q(n29093), .QN(n32933) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n8662), .CK(CLK), .Q(n29094), .QN(n32934) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n8663), .CK(CLK), .Q(n29095), .QN(n32935) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n8664), .CK(CLK), .Q(n29096), .QN(n32936) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n8665), .CK(CLK), .Q(n29097), .QN(n32937)
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n8666), .CK(CLK), .Q(n29098), .QN(n32938)
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n8667), .CK(CLK), .Q(n29099), .QN(n32939)
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n8668), .CK(CLK), .Q(n29100), .QN(n32940)
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n8669), .CK(CLK), .Q(n29101), .QN(n32941)
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n8670), .CK(CLK), .Q(n29102), .QN(n32942)
         );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n9263), .CK(CLK), .Q(n29695), .QN(n38982) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n9264), .CK(CLK), .Q(n29696), .QN(n38981) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n9265), .CK(CLK), .Q(n29697), .QN(n38980) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n9266), .CK(CLK), .Q(n29698), .QN(n38979) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n9267), .CK(CLK), .Q(n29699), .QN(n38978) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n9268), .CK(CLK), .Q(n29700), .QN(n38977) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n9269), .CK(CLK), .Q(n29701), .QN(n38976) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n9270), .CK(CLK), .Q(n29702), .QN(n38975) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n9271), .CK(CLK), .Q(n29703), .QN(n38974) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n9272), .CK(CLK), .Q(n29704), .QN(n38973) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n9273), .CK(CLK), .Q(n29705), .QN(n38972) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n9274), .CK(CLK), .Q(n29706), .QN(n38971) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n9275), .CK(CLK), .Q(n29707), .QN(n38970) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n9276), .CK(CLK), .Q(n29708), .QN(n38969) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n9277), .CK(CLK), .Q(n29709), .QN(n38968) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n9278), .CK(CLK), .Q(n29710), .QN(n38967) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n9279), .CK(CLK), .Q(n29711), .QN(n38966) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n9280), .CK(CLK), .Q(n29712), .QN(n38965) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n9281), .CK(CLK), .Q(n29713), .QN(n38964) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n9282), .CK(CLK), .Q(n29714), .QN(n38963) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n9283), .CK(CLK), .Q(n29715), .QN(n38962) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n9284), .CK(CLK), .Q(n29716), .QN(n38961) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n9285), .CK(CLK), .Q(n29717), .QN(n38960) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n9286), .CK(CLK), .Q(n29718), .QN(n38959) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n9287), .CK(CLK), .Q(n29719), .QN(n38958) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n9288), .CK(CLK), .Q(n29720), .QN(n38957) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n9289), .CK(CLK), .Q(n29721), .QN(n38956) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n9290), .CK(CLK), .Q(n29722), .QN(n38955) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n9291), .CK(CLK), .Q(n29723), .QN(n38954) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n9292), .CK(CLK), .Q(n29724), .QN(n38953) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n9293), .CK(CLK), .Q(n29725), .QN(n38952) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n9294), .CK(CLK), .Q(n29726), .QN(n38951) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n9295), .CK(CLK), .Q(n29727), .QN(n38950) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n9296), .CK(CLK), .Q(n29728), .QN(n38949) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n9297), .CK(CLK), .Q(n29729), .QN(n38948) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n9298), .CK(CLK), .Q(n29730), .QN(n38947) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n9299), .CK(CLK), .Q(n29731), .QN(n38946) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n9300), .CK(CLK), .Q(n29732), .QN(n38945) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n9301), .CK(CLK), .Q(n29733), .QN(n38944) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n9302), .CK(CLK), .Q(n29734), .QN(n38943) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n9303), .CK(CLK), .Q(n29735), .QN(n38942) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n9304), .CK(CLK), .Q(n29736), .QN(n38941) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n9305), .CK(CLK), .Q(n29737), .QN(n38940)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n9306), .CK(CLK), .Q(n29738), .QN(n38939)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n9307), .CK(CLK), .Q(n29739), .QN(n38938)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n9308), .CK(CLK), .Q(n29740), .QN(n38937)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n9309), .CK(CLK), .Q(n29741), .QN(n38936)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n9310), .CK(CLK), .Q(n29742), .QN(n38935)
         );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n8675), .CK(CLK), .Q(n29107), .QN(n33087) );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n8676), .CK(CLK), .Q(n29108), .QN(n33088) );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n8677), .CK(CLK), .Q(n29109), .QN(n33089) );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n8678), .CK(CLK), .Q(n29110), .QN(n33090) );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n8679), .CK(CLK), .Q(n29111), .QN(n33091) );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n8680), .CK(CLK), .Q(n29112), .QN(n33092) );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n8681), .CK(CLK), .Q(n29113), .QN(n33093) );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n8682), .CK(CLK), .Q(n29114), .QN(n33094) );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n8683), .CK(CLK), .Q(n29115), .QN(n33095) );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n8684), .CK(CLK), .Q(n29116), .QN(n33096) );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n8685), .CK(CLK), .Q(n29117), .QN(n33097) );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n8686), .CK(CLK), .Q(n29118), .QN(n33098) );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n8611), .CK(CLK), .Q(n29043), .QN(n33099) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n8612), .CK(CLK), .Q(n29044), .QN(n33100) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n8613), .CK(CLK), .Q(n29045), .QN(n33101) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n8614), .CK(CLK), .Q(n29046), .QN(n33102) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n8615), .CK(CLK), .Q(n29047), .QN(n33103) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n8616), .CK(CLK), .Q(n29048), .QN(n33104) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n8617), .CK(CLK), .Q(n29049), .QN(n33105) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n8618), .CK(CLK), .Q(n29050), .QN(n33106) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n8619), .CK(CLK), .Q(n29051), .QN(n33107) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n8620), .CK(CLK), .Q(n29052), .QN(n33108) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n8621), .CK(CLK), .Q(n29053), .QN(n33109) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n8622), .CK(CLK), .Q(n29054), .QN(n33110) );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n9251), .CK(CLK), .Q(n29683), .QN(n33135) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n9252), .CK(CLK), .Q(n29684), .QN(n33136) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n9253), .CK(CLK), .Q(n29685), .QN(n33137) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n9254), .CK(CLK), .Q(n29686), .QN(n38934) );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n9255), .CK(CLK), .Q(n29687), .QN(n33139) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n9256), .CK(CLK), .Q(n29688), .QN(n38933) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n9257), .CK(CLK), .Q(n29689), .QN(n38932) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n9258), .CK(CLK), .Q(n29690), .QN(n38931) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n9259), .CK(CLK), .Q(n29691), .QN(n38930) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n9260), .CK(CLK), .Q(n29692), .QN(n38929) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n9261), .CK(CLK), .Q(n29693), .QN(n38928) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n9262), .CK(CLK), .Q(n29694), .QN(n38927) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n9327), .CK(CLK), .Q(n29759), .QN(n38849) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n9328), .CK(CLK), .Q(n29760), .QN(n38848) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n9329), .CK(CLK), .Q(n29761), .QN(n38847) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n9330), .CK(CLK), .Q(n29762), .QN(n38846) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n9331), .CK(CLK), .Q(n29763), .QN(n38845) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n9332), .CK(CLK), .Q(n29764), .QN(n38844) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n9333), .CK(CLK), .Q(n29765), .QN(n38843) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n9334), .CK(CLK), .Q(n29766), .QN(n38842) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n9335), .CK(CLK), .Q(n29767), .QN(n38841) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n9336), .CK(CLK), .Q(n29768), .QN(n38840) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n9337), .CK(CLK), .Q(n29769), .QN(n38839) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n9338), .CK(CLK), .Q(n29770), .QN(n38838) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n9339), .CK(CLK), .Q(n29771), .QN(n38837) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n9340), .CK(CLK), .Q(n29772), .QN(n38836) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n9341), .CK(CLK), .Q(n29773), .QN(n38835) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n9342), .CK(CLK), .Q(n29774), .QN(n38834) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n9343), .CK(CLK), .Q(n29775), .QN(n38833) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n9344), .CK(CLK), .Q(n29776), .QN(n38832) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n9345), .CK(CLK), .Q(n29777), .QN(n38831) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n9346), .CK(CLK), .Q(n29778), .QN(n38830) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n9347), .CK(CLK), .Q(n29779), .QN(n38829) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n9348), .CK(CLK), .Q(n29780), .QN(n38828) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n9349), .CK(CLK), .Q(n29781), .QN(n38827) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n9350), .CK(CLK), .Q(n29782), .QN(n38826) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n9351), .CK(CLK), .Q(n29783), .QN(n38825) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n9352), .CK(CLK), .Q(n29784), .QN(n38824) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n9353), .CK(CLK), .Q(n29785), .QN(n38823) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n9354), .CK(CLK), .Q(n29786), .QN(n38822) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n9355), .CK(CLK), .Q(n29787), .QN(n38821) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n9356), .CK(CLK), .Q(n29788), .QN(n38820) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n9357), .CK(CLK), .Q(n29789), .QN(n38819) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n9358), .CK(CLK), .Q(n29790), .QN(n38818) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n9359), .CK(CLK), .Q(n29791), .QN(n38817) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n9360), .CK(CLK), .Q(n29792), .QN(n38816) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n9361), .CK(CLK), .Q(n29793), .QN(n38815) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n9362), .CK(CLK), .Q(n29794), .QN(n38814) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n9363), .CK(CLK), .Q(n29795), .QN(n38813) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n9364), .CK(CLK), .Q(n29796), .QN(n38812) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n9365), .CK(CLK), .Q(n29797), .QN(n38811) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n9366), .CK(CLK), .Q(n29798), .QN(n38810) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n9367), .CK(CLK), .Q(n29799), .QN(n38809) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n9368), .CK(CLK), .Q(n29800), .QN(n38808) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n9369), .CK(CLK), .Q(n29801), .QN(n38807)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n9370), .CK(CLK), .Q(n29802), .QN(n38806)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n9371), .CK(CLK), .Q(n29803), .QN(n38805)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n9372), .CK(CLK), .Q(n29804), .QN(n38804)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n9373), .CK(CLK), .Q(n29805), .QN(n38803)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n9374), .CK(CLK), .Q(n29806), .QN(n38802)
         );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n9315), .CK(CLK), .Q(n29747), .QN(n33195) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n9316), .CK(CLK), .Q(n29748), .QN(n33196) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n9317), .CK(CLK), .Q(n29749), .QN(n33197) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n9318), .CK(CLK), .Q(n29750), .QN(n38801) );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n9319), .CK(CLK), .Q(n29751), .QN(n33199) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n9320), .CK(CLK), .Q(n29752), .QN(n38800) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n9321), .CK(CLK), .Q(n29753), .QN(n38799) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n9322), .CK(CLK), .Q(n29754), .QN(n38798) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n9323), .CK(CLK), .Q(n29755), .QN(n38797) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n9324), .CK(CLK), .Q(n29756), .QN(n38796) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n9325), .CK(CLK), .Q(n29757), .QN(n38795) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n9326), .CK(CLK), .Q(n29758), .QN(n38794) );
  NAND3_X1 U26382 ( .A1(n33212), .A2(n41370), .A3(n2695), .ZN(n33214) );
  XOR2_X1 U26383 ( .A(n32323), .B(n2683), .Z(n33241) );
  NAND3_X1 U26384 ( .A1(n33249), .A2(n32255), .A3(n2709), .ZN(n33248) );
  NAND3_X1 U26385 ( .A1(n32153), .A2(n40581), .A3(n33257), .ZN(n33252) );
  NAND3_X1 U26386 ( .A1(n33257), .A2(n40561), .A3(n32154), .ZN(n33261) );
  NAND3_X1 U26387 ( .A1(n33257), .A2(n40541), .A3(n32155), .ZN(n33266) );
  NAND3_X1 U26388 ( .A1(n33257), .A2(n40521), .A3(n32156), .ZN(n33271) );
  NAND3_X1 U26389 ( .A1(n33257), .A2(n40501), .A3(n33279), .ZN(n33276) );
  NAND3_X1 U26390 ( .A1(n33257), .A2(n40481), .A3(n33284), .ZN(n33281) );
  NAND3_X1 U26391 ( .A1(n33257), .A2(n40461), .A3(n33289), .ZN(n33286) );
  NAND3_X1 U26392 ( .A1(WR), .A2(n32150), .A3(n33294), .ZN(n33256) );
  NAND3_X1 U26393 ( .A1(n33257), .A2(n40441), .A3(n33295), .ZN(n33291) );
  NAND3_X1 U26394 ( .A1(n33297), .A2(ENABLE), .A3(n33298), .ZN(n33259) );
  NAND3_X1 U26395 ( .A1(n33294), .A2(n32150), .A3(n33299), .ZN(n33258) );
  NAND3_X1 U26396 ( .A1(n32153), .A2(n40421), .A3(n33306), .ZN(n33302) );
  NAND3_X1 U26397 ( .A1(n32154), .A2(n40401), .A3(n33306), .ZN(n33309) );
  NAND3_X1 U26398 ( .A1(n32155), .A2(n40381), .A3(n33306), .ZN(n33312) );
  NAND3_X1 U26399 ( .A1(n32156), .A2(n40361), .A3(n33306), .ZN(n33315) );
  NAND3_X1 U26400 ( .A1(n33279), .A2(n40341), .A3(n33306), .ZN(n33318) );
  NAND3_X1 U26401 ( .A1(n33284), .A2(n40321), .A3(n33306), .ZN(n33321) );
  NAND3_X1 U26402 ( .A1(n33289), .A2(n40301), .A3(n33306), .ZN(n33324) );
  NAND3_X1 U26403 ( .A1(N932), .A2(N931), .A3(n33330), .ZN(n33305) );
  NAND3_X1 U26404 ( .A1(n33295), .A2(n40281), .A3(n33306), .ZN(n33327) );
  NAND3_X1 U26405 ( .A1(n32239), .A2(n33332), .A3(N813), .ZN(n33308) );
  NAND3_X1 U26406 ( .A1(N931), .A2(n33333), .A3(N932), .ZN(n33307) );
  NAND3_X1 U26407 ( .A1(n32153), .A2(n40261), .A3(n33338), .ZN(n33334) );
  NAND3_X1 U26408 ( .A1(n32154), .A2(n40241), .A3(n33338), .ZN(n33341) );
  NAND3_X1 U26409 ( .A1(n32155), .A2(n40221), .A3(n33338), .ZN(n33344) );
  NAND3_X1 U26410 ( .A1(n32156), .A2(n40201), .A3(n33338), .ZN(n33347) );
  NAND3_X1 U26411 ( .A1(n33279), .A2(n40181), .A3(n33338), .ZN(n33350) );
  NAND3_X1 U26412 ( .A1(n33284), .A2(n40161), .A3(n33338), .ZN(n33353) );
  NAND3_X1 U26413 ( .A1(n33289), .A2(n40141), .A3(n33338), .ZN(n33356) );
  NAND3_X1 U26414 ( .A1(N932), .A2(n32152), .A3(n33330), .ZN(n33337) );
  NAND3_X1 U26415 ( .A1(n33295), .A2(n40121), .A3(n33338), .ZN(n33359) );
  NAND3_X1 U26416 ( .A1(n32239), .A2(n32247), .A3(n33332), .ZN(n33340) );
  NAND3_X1 U26417 ( .A1(n33333), .A2(n32152), .A3(N932), .ZN(n33339) );
  NAND3_X1 U26418 ( .A1(n32153), .A2(n40101), .A3(n33367), .ZN(n33363) );
  NAND3_X1 U26419 ( .A1(n32154), .A2(n40082), .A3(n33367), .ZN(n33370) );
  NAND3_X1 U26420 ( .A1(n32155), .A2(n40062), .A3(n33367), .ZN(n33373) );
  NAND3_X1 U26421 ( .A1(n32156), .A2(n40042), .A3(n33367), .ZN(n33376) );
  NAND3_X1 U26422 ( .A1(n33279), .A2(n40021), .A3(n33367), .ZN(n33379) );
  NAND3_X1 U26423 ( .A1(n33284), .A2(n40002), .A3(n33367), .ZN(n33382) );
  NAND3_X1 U26424 ( .A1(n33289), .A2(n39984), .A3(n33367), .ZN(n33385) );
  NAND3_X1 U26425 ( .A1(N931), .A2(n32151), .A3(n33330), .ZN(n33366) );
  NAND3_X1 U26426 ( .A1(n33295), .A2(n39964), .A3(n33367), .ZN(n33388) );
  NAND3_X1 U26427 ( .A1(n33332), .A2(n33362), .A3(N813), .ZN(n33369) );
  NAND3_X1 U26428 ( .A1(n33333), .A2(n32151), .A3(N931), .ZN(n33368) );
  NAND3_X1 U26429 ( .A1(n32153), .A2(n39944), .A3(n33395), .ZN(n33391) );
  NAND3_X1 U26430 ( .A1(N811), .A2(n33398), .A3(N812), .ZN(n33260) );
  NAND3_X1 U26432 ( .A1(n32154), .A2(n39923), .A3(n33395), .ZN(n33399) );
  NAND3_X1 U26433 ( .A1(N812), .A2(N811), .A3(n32254), .ZN(n33265) );
  NAND3_X1 U26434 ( .A1(N930), .A2(N929), .A3(n33402), .ZN(n33264) );
  NAND3_X1 U26435 ( .A1(n32155), .A2(n39904), .A3(n33395), .ZN(n33403) );
  NAND3_X1 U26436 ( .A1(n33398), .A2(n32251), .A3(N812), .ZN(n33270) );
  NAND3_X1 U26437 ( .A1(n32163), .A2(n32161), .A3(N930), .ZN(n33269) );
  NAND3_X1 U26438 ( .A1(n32156), .A2(n39886), .A3(n33395), .ZN(n33406) );
  NAND3_X1 U26439 ( .A1(N812), .A2(n32251), .A3(n32254), .ZN(n33275) );
  NAND3_X1 U26440 ( .A1(N930), .A2(n32161), .A3(n33402), .ZN(n33274) );
  NAND3_X1 U26441 ( .A1(n33279), .A2(n39866), .A3(n33395), .ZN(n33409) );
  NAND3_X1 U26442 ( .A1(n33398), .A2(n32249), .A3(N811), .ZN(n33280) );
  NAND3_X1 U26443 ( .A1(n33284), .A2(n39846), .A3(n33395), .ZN(n33412) );
  NAND3_X1 U26444 ( .A1(N811), .A2(n32249), .A3(n32254), .ZN(n33285) );
  NAND3_X1 U26445 ( .A1(n33289), .A2(n39826), .A3(n33395), .ZN(n33415) );
  NAND3_X1 U26446 ( .A1(n32251), .A2(n32249), .A3(n33398), .ZN(n33290) );
  NAND3_X1 U26447 ( .A1(n33295), .A2(n39804), .A3(n33395), .ZN(n33418) );
  NAND3_X1 U26448 ( .A1(n33362), .A2(n32247), .A3(n33332), .ZN(n33396) );
  XOR2_X1 U26449 ( .A(\add_146/carry[4] ), .B(n2695), .Z(n33362) );
  NAND3_X1 U26450 ( .A1(n32251), .A2(n32249), .A3(n32254), .ZN(n33296) );
  XOR2_X1 U26451 ( .A(n33422), .B(\r498/carry[5] ), .Z(n33301) );
  XOR2_X1 U26452 ( .A(n33423), .B(ADD_WR[0]), .Z(n33402) );
  XOR2_X1 U26453 ( .A(n34696), .B(ADD_RD1[0]), .Z(n34694) );
  XOR2_X1 U26454 ( .A(n35970), .B(ADD_RD2[0]), .Z(n35968) );
  XOR2_X1 U26455 ( .A(n27874), .B(n2697), .Z(n33243) );
  XOR2_X1 U26456 ( .A(n27871), .B(n2699), .Z(n33242) );
  XOR2_X1 U26457 ( .A(n27870), .B(n33215), .Z(n35978) );
  XOR2_X1 U26458 ( .A(n32258), .B(N661), .Z(n33245) );
  XOR2_X1 U26459 ( .A(n38790), .B(n2698), .Z(n33239) );
  XOR2_X1 U26460 ( .A(\add_136/carry[4] ), .B(n2695), .Z(n37240) );
  NAND3_X1 U26461 ( .A1(\i[1] ), .A2(n32255), .A3(n33249), .ZN(n33250) );
  DFF_X1 \CWP_reg[3]  ( .D(n9904), .CK(CLK), .Q(N661), .QN(n2696) );
  DFF_X1 \CWP_reg[2]  ( .D(n9905), .CK(CLK), .Q(N660), .QN(n2697) );
  DFF_X1 \CWP_reg[1]  ( .D(n9906), .CK(CLK), .Q(N659), .QN(n2698) );
  DFF_X1 \i_reg[3]  ( .D(n25394), .CK(CLK), .Q(\i[3] ), .QN(n2706) );
  DFF_X1 \i_reg[1]  ( .D(n9892), .CK(CLK), .Q(\i[1] ), .QN(n2709) );
  DFF_X1 \i_reg[2]  ( .D(n9891), .CK(CLK), .Q(\i[2] ), .QN(n2707) );
  DFF_X1 STORE_DATA_reg ( .D(n7202), .CK(CLK), .Q(SPILL), .QN(n2700) );
  DFF_X1 RETRIEVE_DATA_reg ( .D(n9893), .CK(CLK), .Q(FILL), .QN(n23853) );
  DFF_X1 \BUSout_reg[63]  ( .D(n7201), .CK(CLK), .Q(BUSout[63]), .QN(n16941)
         );
  DFF_X1 \BUSout_reg[62]  ( .D(n7200), .CK(CLK), .Q(BUSout[62]), .QN(n16940)
         );
  DFF_X1 \BUSout_reg[61]  ( .D(n7199), .CK(CLK), .Q(BUSout[61]), .QN(n16939)
         );
  DFF_X1 \BUSout_reg[60]  ( .D(n7198), .CK(CLK), .Q(BUSout[60]), .QN(n16938)
         );
  DFF_X1 \BUSout_reg[5]  ( .D(n7143), .CK(CLK), .Q(BUSout[5]), .QN(n16883) );
  DFF_X1 \BUSout_reg[4]  ( .D(n7142), .CK(CLK), .Q(BUSout[4]), .QN(n16882) );
  DFF_X1 \BUSout_reg[3]  ( .D(n7141), .CK(CLK), .Q(BUSout[3]), .QN(n16881) );
  DFF_X1 \BUSout_reg[2]  ( .D(n7140), .CK(CLK), .Q(BUSout[2]), .QN(n16880) );
  DFF_X1 \BUSout_reg[1]  ( .D(n7139), .CK(CLK), .Q(BUSout[1]), .QN(n16879) );
  DFF_X1 \BUSout_reg[53]  ( .D(n7191), .CK(CLK), .Q(BUSout[53]), .QN(n16931)
         );
  DFF_X1 \BUSout_reg[52]  ( .D(n7190), .CK(CLK), .Q(BUSout[52]), .QN(n16930)
         );
  DFF_X1 \BUSout_reg[51]  ( .D(n7189), .CK(CLK), .Q(BUSout[51]), .QN(n16929)
         );
  DFF_X1 \BUSout_reg[50]  ( .D(n7188), .CK(CLK), .Q(BUSout[50]), .QN(n16928)
         );
  DFF_X1 \BUSout_reg[49]  ( .D(n7187), .CK(CLK), .Q(BUSout[49]), .QN(n16927)
         );
  DFF_X1 \BUSout_reg[48]  ( .D(n7186), .CK(CLK), .Q(BUSout[48]), .QN(n16926)
         );
  DFF_X1 \BUSout_reg[47]  ( .D(n7185), .CK(CLK), .Q(BUSout[47]), .QN(n16925)
         );
  DFF_X1 \BUSout_reg[46]  ( .D(n7184), .CK(CLK), .Q(BUSout[46]), .QN(n16924)
         );
  DFF_X1 \BUSout_reg[45]  ( .D(n7183), .CK(CLK), .Q(BUSout[45]), .QN(n16923)
         );
  DFF_X1 \BUSout_reg[44]  ( .D(n7182), .CK(CLK), .Q(BUSout[44]), .QN(n16922)
         );
  DFF_X1 \BUSout_reg[43]  ( .D(n7181), .CK(CLK), .Q(BUSout[43]), .QN(n16921)
         );
  DFF_X1 \BUSout_reg[42]  ( .D(n7180), .CK(CLK), .Q(BUSout[42]), .QN(n16920)
         );
  DFF_X1 \BUSout_reg[41]  ( .D(n7179), .CK(CLK), .Q(BUSout[41]), .QN(n16919)
         );
  DFF_X1 \BUSout_reg[40]  ( .D(n7178), .CK(CLK), .Q(BUSout[40]), .QN(n16918)
         );
  DFF_X1 \BUSout_reg[39]  ( .D(n7177), .CK(CLK), .Q(BUSout[39]), .QN(n16917)
         );
  DFF_X1 \BUSout_reg[38]  ( .D(n7176), .CK(CLK), .Q(BUSout[38]), .QN(n16916)
         );
  DFF_X1 \BUSout_reg[37]  ( .D(n7175), .CK(CLK), .Q(BUSout[37]), .QN(n16915)
         );
  DFF_X1 \BUSout_reg[36]  ( .D(n7174), .CK(CLK), .Q(BUSout[36]), .QN(n16914)
         );
  DFF_X1 \BUSout_reg[35]  ( .D(n7173), .CK(CLK), .Q(BUSout[35]), .QN(n16913)
         );
  DFF_X1 \BUSout_reg[34]  ( .D(n7172), .CK(CLK), .Q(BUSout[34]), .QN(n16912)
         );
  DFF_X1 \BUSout_reg[33]  ( .D(n7171), .CK(CLK), .Q(BUSout[33]), .QN(n16911)
         );
  DFF_X1 \BUSout_reg[32]  ( .D(n7170), .CK(CLK), .Q(BUSout[32]), .QN(n16910)
         );
  DFF_X1 \BUSout_reg[31]  ( .D(n7169), .CK(CLK), .Q(BUSout[31]), .QN(n16909)
         );
  DFF_X1 \BUSout_reg[30]  ( .D(n7168), .CK(CLK), .Q(BUSout[30]), .QN(n16908)
         );
  DFF_X1 \BUSout_reg[29]  ( .D(n7167), .CK(CLK), .Q(BUSout[29]), .QN(n16907)
         );
  DFF_X1 \BUSout_reg[28]  ( .D(n7166), .CK(CLK), .Q(BUSout[28]), .QN(n16906)
         );
  DFF_X1 \BUSout_reg[27]  ( .D(n7165), .CK(CLK), .Q(BUSout[27]), .QN(n16905)
         );
  DFF_X1 \BUSout_reg[26]  ( .D(n7164), .CK(CLK), .Q(BUSout[26]), .QN(n16904)
         );
  DFF_X1 \BUSout_reg[25]  ( .D(n7163), .CK(CLK), .Q(BUSout[25]), .QN(n16903)
         );
  DFF_X1 \BUSout_reg[24]  ( .D(n7162), .CK(CLK), .Q(BUSout[24]), .QN(n16902)
         );
  DFF_X1 \BUSout_reg[23]  ( .D(n7161), .CK(CLK), .Q(BUSout[23]), .QN(n16901)
         );
  DFF_X1 \BUSout_reg[22]  ( .D(n7160), .CK(CLK), .Q(BUSout[22]), .QN(n16900)
         );
  DFF_X1 \BUSout_reg[21]  ( .D(n7159), .CK(CLK), .Q(BUSout[21]), .QN(n16899)
         );
  DFF_X1 \BUSout_reg[20]  ( .D(n7158), .CK(CLK), .Q(BUSout[20]), .QN(n16898)
         );
  DFF_X1 \BUSout_reg[19]  ( .D(n7157), .CK(CLK), .Q(BUSout[19]), .QN(n16897)
         );
  DFF_X1 \BUSout_reg[18]  ( .D(n7156), .CK(CLK), .Q(BUSout[18]), .QN(n16896)
         );
  DFF_X1 \BUSout_reg[17]  ( .D(n7155), .CK(CLK), .Q(BUSout[17]), .QN(n16895)
         );
  DFF_X1 \BUSout_reg[16]  ( .D(n7154), .CK(CLK), .Q(BUSout[16]), .QN(n16894)
         );
  DFF_X1 \BUSout_reg[15]  ( .D(n7153), .CK(CLK), .Q(BUSout[15]), .QN(n16893)
         );
  DFF_X1 \BUSout_reg[14]  ( .D(n7152), .CK(CLK), .Q(BUSout[14]), .QN(n16892)
         );
  DFF_X1 \BUSout_reg[13]  ( .D(n7151), .CK(CLK), .Q(BUSout[13]), .QN(n16891)
         );
  DFF_X1 \BUSout_reg[12]  ( .D(n7150), .CK(CLK), .Q(BUSout[12]), .QN(n16890)
         );
  DFF_X1 \BUSout_reg[11]  ( .D(n7149), .CK(CLK), .Q(BUSout[11]), .QN(n16889)
         );
  DFF_X1 \BUSout_reg[10]  ( .D(n7148), .CK(CLK), .Q(BUSout[10]), .QN(n16888)
         );
  DFF_X1 \BUSout_reg[9]  ( .D(n7147), .CK(CLK), .Q(BUSout[9]), .QN(n16887) );
  DFF_X1 \BUSout_reg[8]  ( .D(n7146), .CK(CLK), .Q(BUSout[8]), .QN(n16886) );
  DFF_X1 \BUSout_reg[7]  ( .D(n7145), .CK(CLK), .Q(BUSout[7]), .QN(n16885) );
  DFF_X1 \BUSout_reg[6]  ( .D(n7144), .CK(CLK), .Q(BUSout[6]), .QN(n16884) );
  DFF_X1 \SWP_reg[4]  ( .D(n9896), .CK(CLK), .Q(n27872), .QN(n32322) );
  DFF_X1 \SWP_reg[3]  ( .D(n9897), .CK(CLK), .Q(n38789), .QN(n32258) );
  DFF_X1 \SWP_reg[1]  ( .D(n9899), .CK(CLK), .Q(n38790), .QN(n32260) );
  DFF_X1 \SWP_reg[5]  ( .D(n9901), .CK(CLK), .Q(n27870), .QN(n32323) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n7583), .CK(CLK), .QN(n30605) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n7584), .CK(CLK), .QN(n30606) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n7585), .CK(CLK), .QN(n30607) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n7586), .CK(CLK), .QN(n30608) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n7519), .CK(CLK), .QN(n30541) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n7520), .CK(CLK), .QN(n30542) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n7521), .CK(CLK), .QN(n30543) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n7522), .CK(CLK), .QN(n30544) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n7455), .CK(CLK), .Q(n28004), .QN(n32456)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n7456), .CK(CLK), .Q(n28005), .QN(n32457)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n7457), .CK(CLK), .Q(n28006), .QN(n32458)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n7458), .CK(CLK), .Q(n28007), .QN(n32459)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n7647), .CK(CLK), .QN(n30669) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n7648), .CK(CLK), .QN(n30670) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n7649), .CK(CLK), .QN(n30671) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n7650), .CK(CLK), .QN(n30672) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n7839), .CK(CLK), .QN(n30733) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n7840), .CK(CLK), .QN(n30734) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n7841), .CK(CLK), .QN(n30735) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n7842), .CK(CLK), .QN(n30736) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n7967), .CK(CLK), .QN(n30861) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n7968), .CK(CLK), .QN(n30862) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n7969), .CK(CLK), .QN(n30863) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n7970), .CK(CLK), .QN(n30864) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n7903), .CK(CLK), .QN(n30797) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n7904), .CK(CLK), .QN(n30798) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n7905), .CK(CLK), .QN(n30799) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n7906), .CK(CLK), .QN(n30800) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n8607), .CK(CLK), .QN(n31363) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n8608), .CK(CLK), .QN(n31364) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n8609), .CK(CLK), .QN(n31365) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n8610), .CK(CLK), .QN(n31366) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n8543), .CK(CLK), .QN(n31299) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n8544), .CK(CLK), .QN(n31300) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n8545), .CK(CLK), .QN(n31301) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n8546), .CK(CLK), .QN(n31302) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n8479), .CK(CLK), .QN(n31235) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n8480), .CK(CLK), .QN(n31236) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n8481), .CK(CLK), .QN(n31237) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n8482), .CK(CLK), .QN(n31238) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n7526), .CK(CLK), .QN(n30548) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n7528), .CK(CLK), .QN(n30550) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n7529), .CK(CLK), .QN(n30551) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n7530), .CK(CLK), .QN(n30552) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n7531), .CK(CLK), .QN(n30553) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n7532), .CK(CLK), .QN(n30554) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n7533), .CK(CLK), .QN(n30555) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n7534), .CK(CLK), .QN(n30556) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n7535), .CK(CLK), .QN(n30557) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n7536), .CK(CLK), .QN(n30558) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n7537), .CK(CLK), .QN(n30559) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n7538), .CK(CLK), .QN(n30560) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n7539), .CK(CLK), .QN(n30561) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n7540), .CK(CLK), .QN(n30562) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n7541), .CK(CLK), .QN(n30563) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n7542), .CK(CLK), .QN(n30564) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n7543), .CK(CLK), .QN(n30565) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n7544), .CK(CLK), .QN(n30566) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n7545), .CK(CLK), .QN(n30567) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n7546), .CK(CLK), .QN(n30568) );
  DFF_X1 \CWP_reg[4]  ( .D(n9903), .CK(CLK), .Q(n32242), .QN(n2695) );
  DFF_X1 \CWP_reg[5]  ( .D(n9902), .CK(CLK), .Q(n32244), .QN(n2683) );
  DFF_X1 \i_reg[0]  ( .D(n9895), .CK(CLK), .Q(n32255), .QN(n2710) );
  DFF_X1 \CWP_reg[0]  ( .D(n9907), .CK(CLK), .Q(n32253), .QN(n2699) );
  DFF_X1 \SWP_reg[2]  ( .D(n9898), .CK(CLK), .Q(n32259), .QN(n27874) );
  DFF_X1 \SWP_reg[0]  ( .D(n9900), .CK(CLK), .Q(n32261), .QN(n27871) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n7775), .CK(CLK), .Q(n32484), .QN(n503) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n7776), .CK(CLK), .Q(n32485), .QN(n504) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n7777), .CK(CLK), .Q(n32486), .QN(n505) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n7778), .CK(CLK), .Q(n32487), .QN(n506) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n7711), .CK(CLK), .Q(n32488), .QN(n439) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n7712), .CK(CLK), .Q(n32489), .QN(n440) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n7713), .CK(CLK), .Q(n32490), .QN(n441) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n7714), .CK(CLK), .Q(n32491), .QN(n442) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n7391), .CK(CLK), .Q(n30477), .QN(n27940)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n7392), .CK(CLK), .Q(n30478), .QN(n27941)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n7393), .CK(CLK), .Q(n30479), .QN(n27942)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n7394), .CK(CLK), .Q(n30480), .QN(n27943)
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n8095), .CK(CLK), .Q(n32468), .QN(n823)
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n8096), .CK(CLK), .Q(n32469), .QN(n824)
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n8097), .CK(CLK), .Q(n32470), .QN(n825)
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n8098), .CK(CLK), .Q(n32471), .QN(n826)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n8031), .CK(CLK), .Q(n32472), .QN(n759)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n8032), .CK(CLK), .Q(n32473), .QN(n760)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n8033), .CK(CLK), .Q(n32474), .QN(n761)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n8034), .CK(CLK), .Q(n32475), .QN(n762)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n8351), .CK(CLK), .Q(n31117), .QN(n25401)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n8352), .CK(CLK), .Q(n31118), .QN(n25400)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n8353), .CK(CLK), .Q(n31119), .QN(n25399)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n8354), .CK(CLK), .Q(n31120), .QN(n25398)
         );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n7727), .CK(CLK), .Q(n32943), .QN(n455)
         );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n7728), .CK(CLK), .Q(n32944), .QN(n456)
         );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n7729), .CK(CLK), .Q(n32945), .QN(n457)
         );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n7730), .CK(CLK), .Q(n32946), .QN(n458)
         );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n7731), .CK(CLK), .Q(n32947), .QN(n459)
         );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n7732), .CK(CLK), .Q(n32948), .QN(n460)
         );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n7733), .CK(CLK), .Q(n32949), .QN(n461)
         );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n7734), .CK(CLK), .Q(n32950), .QN(n462)
         );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n7735), .CK(CLK), .Q(n32951), .QN(n463)
         );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n7736), .CK(CLK), .Q(n32952), .QN(n464)
         );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n7737), .CK(CLK), .Q(n32953), .QN(n465)
         );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n7738), .CK(CLK), .Q(n32954), .QN(n466)
         );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n7739), .CK(CLK), .Q(n32955), .QN(n467)
         );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n7740), .CK(CLK), .Q(n32956), .QN(n468)
         );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n7741), .CK(CLK), .Q(n32957), .QN(n469)
         );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n7742), .CK(CLK), .Q(n32958), .QN(n470)
         );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n7743), .CK(CLK), .Q(n32959), .QN(n471)
         );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n7744), .CK(CLK), .Q(n32960), .QN(n472)
         );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n7745), .CK(CLK), .Q(n32961), .QN(n473)
         );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n7746), .CK(CLK), .Q(n32962), .QN(n474)
         );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n7747), .CK(CLK), .Q(n32963), .QN(n475)
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n7748), .CK(CLK), .Q(n32964), .QN(n476)
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n7749), .CK(CLK), .Q(n32965), .QN(n477)
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n7750), .CK(CLK), .Q(n32966), .QN(n478)
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n7751), .CK(CLK), .Q(n32967), .QN(n479)
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n7752), .CK(CLK), .Q(n32968), .QN(n480)
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n7753), .CK(CLK), .Q(n32969), .QN(n481)
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n7754), .CK(CLK), .Q(n32970), .QN(n482)
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n7755), .CK(CLK), .Q(n32971), .QN(n483)
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n7756), .CK(CLK), .Q(n32972), .QN(n484)
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n7757), .CK(CLK), .Q(n32973), .QN(n485)
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n7758), .CK(CLK), .Q(n32974), .QN(n486)
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n7759), .CK(CLK), .Q(n32975), .QN(n487)
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n7760), .CK(CLK), .Q(n32976), .QN(n488)
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n7761), .CK(CLK), .Q(n32977), .QN(n489)
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n7762), .CK(CLK), .Q(n32978), .QN(n490)
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n7763), .CK(CLK), .Q(n32979), .QN(n491)
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n7764), .CK(CLK), .Q(n32980), .QN(n492)
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n7765), .CK(CLK), .Q(n32981), .QN(n493)
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n7766), .CK(CLK), .Q(n32982), .QN(n494)
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n7767), .CK(CLK), .Q(n32983), .QN(n495)
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n7768), .CK(CLK), .Q(n32984), .QN(n496)
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n7769), .CK(CLK), .Q(n32985), .QN(n497) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n7770), .CK(CLK), .Q(n32986), .QN(n498) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n7771), .CK(CLK), .Q(n32987), .QN(n499) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n7772), .CK(CLK), .Q(n32988), .QN(n500) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n7773), .CK(CLK), .Q(n32989), .QN(n501) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n7774), .CK(CLK), .Q(n32990), .QN(n502) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n7715), .CK(CLK), .Q(n33111), .QN(n443)
         );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n7716), .CK(CLK), .Q(n33112), .QN(n444)
         );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n7717), .CK(CLK), .Q(n33113), .QN(n445)
         );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n7718), .CK(CLK), .Q(n33114), .QN(n446)
         );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n7719), .CK(CLK), .Q(n33115), .QN(n447)
         );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n7720), .CK(CLK), .Q(n33116), .QN(n448)
         );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n7721), .CK(CLK), .Q(n33117), .QN(n449)
         );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n7722), .CK(CLK), .Q(n33118), .QN(n450)
         );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n7723), .CK(CLK), .Q(n33119), .QN(n451)
         );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n7724), .CK(CLK), .Q(n33120), .QN(n452)
         );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n7725), .CK(CLK), .Q(n33121), .QN(n453)
         );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n7726), .CK(CLK), .Q(n33122), .QN(n454)
         );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n7663), .CK(CLK), .Q(n32991), .QN(n391)
         );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n7664), .CK(CLK), .Q(n32992), .QN(n392)
         );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n7665), .CK(CLK), .Q(n32993), .QN(n393)
         );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n7666), .CK(CLK), .Q(n32994), .QN(n394)
         );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n7667), .CK(CLK), .Q(n32995), .QN(n395)
         );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n7668), .CK(CLK), .Q(n32996), .QN(n396)
         );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n7669), .CK(CLK), .Q(n32997), .QN(n397)
         );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n7670), .CK(CLK), .Q(n32998), .QN(n398)
         );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n7671), .CK(CLK), .Q(n32999), .QN(n399)
         );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n7672), .CK(CLK), .Q(n33000), .QN(n400)
         );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n7673), .CK(CLK), .Q(n33001), .QN(n401)
         );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n7674), .CK(CLK), .Q(n33002), .QN(n402)
         );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n7675), .CK(CLK), .Q(n33003), .QN(n403)
         );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n7676), .CK(CLK), .Q(n33004), .QN(n404)
         );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n7677), .CK(CLK), .Q(n33005), .QN(n405)
         );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n7678), .CK(CLK), .Q(n33006), .QN(n406)
         );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n7679), .CK(CLK), .Q(n33007), .QN(n407)
         );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n7680), .CK(CLK), .Q(n33008), .QN(n408)
         );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n7681), .CK(CLK), .Q(n33009), .QN(n409)
         );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n7682), .CK(CLK), .Q(n33010), .QN(n410)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n7683), .CK(CLK), .Q(n33011), .QN(n411)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n7684), .CK(CLK), .Q(n33012), .QN(n412)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n7685), .CK(CLK), .Q(n33013), .QN(n413)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n7686), .CK(CLK), .Q(n33014), .QN(n414)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n7687), .CK(CLK), .Q(n33015), .QN(n415)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n7688), .CK(CLK), .Q(n33016), .QN(n416)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n7689), .CK(CLK), .Q(n33017), .QN(n417)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n7690), .CK(CLK), .Q(n33018), .QN(n418)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n7691), .CK(CLK), .Q(n33019), .QN(n419)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n7692), .CK(CLK), .Q(n33020), .QN(n420)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n7693), .CK(CLK), .Q(n33021), .QN(n421)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n7694), .CK(CLK), .Q(n33022), .QN(n422)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n7695), .CK(CLK), .Q(n33023), .QN(n423)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n7696), .CK(CLK), .Q(n33024), .QN(n424)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n7697), .CK(CLK), .Q(n33025), .QN(n425)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n7698), .CK(CLK), .Q(n33026), .QN(n426)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n7699), .CK(CLK), .Q(n33027), .QN(n427)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n7700), .CK(CLK), .Q(n33028), .QN(n428)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n7701), .CK(CLK), .Q(n33029), .QN(n429)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n7702), .CK(CLK), .Q(n33030), .QN(n430)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n7703), .CK(CLK), .Q(n33031), .QN(n431)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n7704), .CK(CLK), .Q(n33032), .QN(n432)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n7705), .CK(CLK), .Q(n33033), .QN(n433) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n7706), .CK(CLK), .Q(n33034), .QN(n434) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n7707), .CK(CLK), .Q(n33035), .QN(n435) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n7708), .CK(CLK), .Q(n33036), .QN(n436) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n7709), .CK(CLK), .Q(n33037), .QN(n437) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n7710), .CK(CLK), .Q(n33038), .QN(n438) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n7651), .CK(CLK), .Q(n33123), .QN(n379)
         );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n7652), .CK(CLK), .Q(n33124), .QN(n380)
         );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n7653), .CK(CLK), .Q(n33125), .QN(n381)
         );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n7654), .CK(CLK), .Q(n33126), .QN(n382)
         );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n7655), .CK(CLK), .Q(n33127), .QN(n383)
         );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n7656), .CK(CLK), .Q(n33128), .QN(n384)
         );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n7657), .CK(CLK), .Q(n33129), .QN(n385)
         );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n7658), .CK(CLK), .Q(n33130), .QN(n386)
         );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n7659), .CK(CLK), .Q(n33131), .QN(n387)
         );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n7660), .CK(CLK), .Q(n33132), .QN(n388)
         );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n7661), .CK(CLK), .Q(n33133), .QN(n389)
         );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n7662), .CK(CLK), .Q(n33134), .QN(n390)
         );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n8357), .CK(CLK), .Q(n31123), .QN(n25509) );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n8355), .CK(CLK), .Q(n31121), .QN(n25511) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n8356), .CK(CLK), .Q(n31122), .QN(n25510) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n8358), .CK(CLK), .Q(n31124), .QN(n25508) );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n8359), .CK(CLK), .Q(n31125), .QN(n25507) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n8360), .CK(CLK), .Q(n31126), .QN(n25506) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n8361), .CK(CLK), .Q(n31127), .QN(n25505) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n8362), .CK(CLK), .Q(n31128), .QN(n25504) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n8363), .CK(CLK), .Q(n31129), .QN(n25503) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n8364), .CK(CLK), .Q(n31130), .QN(n25502) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n8365), .CK(CLK), .Q(n31131), .QN(n25501) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n8366), .CK(CLK), .Q(n31132), .QN(n25500) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n8367), .CK(CLK), .Q(n31133), .QN(n25499) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n8368), .CK(CLK), .Q(n31134), .QN(n25498) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n8369), .CK(CLK), .Q(n31135), .QN(n25497) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n8370), .CK(CLK), .Q(n31136), .QN(n25496) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n8371), .CK(CLK), .Q(n31137), .QN(n25495) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n8372), .CK(CLK), .Q(n31138), .QN(n25494) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n8373), .CK(CLK), .Q(n31139), .QN(n25493) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n8374), .CK(CLK), .Q(n31140), .QN(n25492) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n8375), .CK(CLK), .Q(n31141), .QN(n25491) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n8376), .CK(CLK), .Q(n31142), .QN(n25490) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n8377), .CK(CLK), .Q(n31143), .QN(n25489) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n8378), .CK(CLK), .Q(n31144), .QN(n25488) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n8379), .CK(CLK), .Q(n31145), .QN(n25487) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n8380), .CK(CLK), .Q(n31146), .QN(n25486) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n8381), .CK(CLK), .Q(n31147), .QN(n25485) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n8382), .CK(CLK), .Q(n31148), .QN(n25484) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n8383), .CK(CLK), .Q(n31149), .QN(n25483) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n8384), .CK(CLK), .Q(n31150), .QN(n25482) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n8385), .CK(CLK), .Q(n31151), .QN(n25481) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n8386), .CK(CLK), .Q(n31152), .QN(n25480) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n8387), .CK(CLK), .Q(n31153), .QN(n25479) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n8388), .CK(CLK), .Q(n31154), .QN(n25478) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n8389), .CK(CLK), .Q(n31155), .QN(n25477) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n8390), .CK(CLK), .Q(n31156), .QN(n25476) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n8391), .CK(CLK), .Q(n31157), .QN(n25475) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n8392), .CK(CLK), .Q(n31158), .QN(n25474) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n8393), .CK(CLK), .Q(n31159), .QN(n25473) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n8394), .CK(CLK), .Q(n31160), .QN(n25472) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n8395), .CK(CLK), .Q(n31161), .QN(n25471) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n8396), .CK(CLK), .Q(n31162), .QN(n25470) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n8397), .CK(CLK), .Q(n31163), .QN(n25469) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n8398), .CK(CLK), .Q(n31164), .QN(n25468) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n8399), .CK(CLK), .Q(n31165), .QN(n25467) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n8400), .CK(CLK), .Q(n31166), .QN(n25466) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n8401), .CK(CLK), .Q(n31167), .QN(n25465) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n8402), .CK(CLK), .Q(n31168), .QN(n25464) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n8403), .CK(CLK), .Q(n31169), .QN(n25463) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n8404), .CK(CLK), .Q(n31170), .QN(n25462) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n8405), .CK(CLK), .Q(n31171), .QN(n25461) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n8406), .CK(CLK), .Q(n31172), .QN(n25460) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n8407), .CK(CLK), .Q(n31173), .QN(n25459) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n8408), .CK(CLK), .Q(n31174), .QN(n25458) );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7343), .CK(CLK), .Q(n32518), .QN(n71) );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7344), .CK(CLK), .Q(n32519), .QN(n72) );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7345), .CK(CLK), .Q(n32520), .QN(n73) );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7346), .CK(CLK), .Q(n32521), .QN(n74) );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7347), .CK(CLK), .Q(n32522), .QN(n75) );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7348), .CK(CLK), .Q(n32523), .QN(n76) );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7349), .CK(CLK), .Q(n32524), .QN(n77) );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7350), .CK(CLK), .Q(n32525), .QN(n78) );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7351), .CK(CLK), .Q(n32526), .QN(n79) );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7352), .CK(CLK), .Q(n32527), .QN(n80) );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7353), .CK(CLK), .Q(n32528), .QN(n81) );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7354), .CK(CLK), .Q(n32529), .QN(n82) );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7355), .CK(CLK), .Q(n32530), .QN(n83) );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7356), .CK(CLK), .Q(n32531), .QN(n84) );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7357), .CK(CLK), .Q(n32532), .QN(n85) );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7358), .CK(CLK), .Q(n32533), .QN(n86) );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7359), .CK(CLK), .Q(n32534), .QN(n87) );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7360), .CK(CLK), .Q(n32535), .QN(n88) );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7361), .CK(CLK), .Q(n32536), .QN(n89) );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7362), .CK(CLK), .Q(n32537), .QN(n90) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7363), .CK(CLK), .Q(n32538), .QN(n91) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7364), .CK(CLK), .Q(n32539), .QN(n92) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7365), .CK(CLK), .Q(n32540), .QN(n93) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7366), .CK(CLK), .Q(n32541), .QN(n94) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7367), .CK(CLK), .Q(n32542), .QN(n95) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7368), .CK(CLK), .Q(n32543), .QN(n96) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7369), .CK(CLK), .Q(n32544), .QN(n97) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7370), .CK(CLK), .Q(n32545), .QN(n98) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7371), .CK(CLK), .Q(n32546), .QN(n99) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7372), .CK(CLK), .Q(n30458), .QN(n27921)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7373), .CK(CLK), .Q(n30459), .QN(n27922)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7374), .CK(CLK), .Q(n30460), .QN(n27923)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7375), .CK(CLK), .Q(n30461), .QN(n27924)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7376), .CK(CLK), .Q(n30462), .QN(n27925)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7377), .CK(CLK), .Q(n30463), .QN(n27926)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7378), .CK(CLK), .Q(n30464), .QN(n27927)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7379), .CK(CLK), .Q(n30465), .QN(n27928)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7380), .CK(CLK), .Q(n30466), .QN(n27929)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7381), .CK(CLK), .Q(n30467), .QN(n27930)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7382), .CK(CLK), .Q(n30468), .QN(n27931)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n7383), .CK(CLK), .Q(n30469), .QN(n27932)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n7384), .CK(CLK), .Q(n30470), .QN(n27933)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n7385), .CK(CLK), .Q(n30471), .QN(n27934)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n7386), .CK(CLK), .Q(n30472), .QN(n27935)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n7387), .CK(CLK), .Q(n30473), .QN(n27936)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n7388), .CK(CLK), .Q(n30474), .QN(n27937)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n7389), .CK(CLK), .Q(n30475), .QN(n27938)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n7390), .CK(CLK), .Q(n30476), .QN(n27939)
         );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7331), .CK(CLK), .Q(n32508), .QN(n59) );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7332), .CK(CLK), .Q(n32509), .QN(n60) );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7333), .CK(CLK), .Q(n32506), .QN(n61) );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7334), .CK(CLK), .Q(n32507), .QN(n62) );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7335), .CK(CLK), .Q(n32510), .QN(n63) );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7336), .CK(CLK), .Q(n32511), .QN(n64) );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7337), .CK(CLK), .Q(n32512), .QN(n65) );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7338), .CK(CLK), .Q(n32513), .QN(n66) );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7339), .CK(CLK), .Q(n32514), .QN(n67) );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7340), .CK(CLK), .Q(n32515), .QN(n68) );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7341), .CK(CLK), .Q(n32516), .QN(n69) );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7342), .CK(CLK), .Q(n32517), .QN(n70) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n8047), .CK(CLK), .Q(n32727), .QN(n775)
         );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n8048), .CK(CLK), .Q(n32728), .QN(n776)
         );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n8049), .CK(CLK), .Q(n32729), .QN(n777)
         );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n8050), .CK(CLK), .Q(n32730), .QN(n778)
         );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n8051), .CK(CLK), .Q(n32731), .QN(n779)
         );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n8052), .CK(CLK), .Q(n32732), .QN(n780)
         );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n8053), .CK(CLK), .Q(n32733), .QN(n781)
         );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n8054), .CK(CLK), .Q(n32734), .QN(n782)
         );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n8055), .CK(CLK), .Q(n32735), .QN(n783)
         );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n8056), .CK(CLK), .Q(n32736), .QN(n784)
         );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n8057), .CK(CLK), .Q(n32737), .QN(n785)
         );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n8058), .CK(CLK), .Q(n32738), .QN(n786)
         );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n8059), .CK(CLK), .Q(n32739), .QN(n787)
         );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n8060), .CK(CLK), .Q(n32740), .QN(n788)
         );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n8061), .CK(CLK), .Q(n32741), .QN(n789)
         );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n8062), .CK(CLK), .Q(n32742), .QN(n790)
         );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n8063), .CK(CLK), .Q(n32743), .QN(n791)
         );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n8064), .CK(CLK), .Q(n32744), .QN(n792)
         );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n8065), .CK(CLK), .Q(n32745), .QN(n793)
         );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n8066), .CK(CLK), .Q(n32746), .QN(n794)
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n8067), .CK(CLK), .Q(n32747), .QN(n795)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n8068), .CK(CLK), .Q(n32748), .QN(n796)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n8069), .CK(CLK), .Q(n32749), .QN(n797)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n8070), .CK(CLK), .Q(n32750), .QN(n798)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n8071), .CK(CLK), .Q(n32751), .QN(n799)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n8072), .CK(CLK), .Q(n32752), .QN(n800)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n8073), .CK(CLK), .Q(n32753), .QN(n801)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n8074), .CK(CLK), .Q(n32754), .QN(n802)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n8075), .CK(CLK), .Q(n32755), .QN(n803)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n8076), .CK(CLK), .Q(n32756), .QN(n804)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n8077), .CK(CLK), .Q(n32757), .QN(n805)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n8078), .CK(CLK), .Q(n32758), .QN(n806)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n8079), .CK(CLK), .Q(n32759), .QN(n807)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n8080), .CK(CLK), .Q(n32760), .QN(n808)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n8081), .CK(CLK), .Q(n32761), .QN(n809)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n8082), .CK(CLK), .Q(n32762), .QN(n810)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n8083), .CK(CLK), .Q(n32763), .QN(n811)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n8084), .CK(CLK), .Q(n32764), .QN(n812)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n8085), .CK(CLK), .Q(n32765), .QN(n813)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n8086), .CK(CLK), .Q(n32766), .QN(n814)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n8087), .CK(CLK), .Q(n32767), .QN(n815)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n8088), .CK(CLK), .Q(n32768), .QN(n816)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n8089), .CK(CLK), .Q(n32769), .QN(n817)
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n8090), .CK(CLK), .Q(n32770), .QN(n818)
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n8091), .CK(CLK), .Q(n32771), .QN(n819)
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n8092), .CK(CLK), .Q(n32772), .QN(n820)
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n8093), .CK(CLK), .Q(n32773), .QN(n821)
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n8094), .CK(CLK), .Q(n32774), .QN(n822)
         );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n7983), .CK(CLK), .Q(n32775), .QN(n711)
         );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n7984), .CK(CLK), .Q(n32776), .QN(n712)
         );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n7985), .CK(CLK), .Q(n32777), .QN(n713)
         );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n7986), .CK(CLK), .Q(n32778), .QN(n714)
         );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n7987), .CK(CLK), .Q(n32779), .QN(n715)
         );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n7988), .CK(CLK), .Q(n32780), .QN(n716)
         );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n7989), .CK(CLK), .Q(n32781), .QN(n717)
         );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n7990), .CK(CLK), .Q(n32782), .QN(n718)
         );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n7991), .CK(CLK), .Q(n32783), .QN(n719)
         );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n7992), .CK(CLK), .Q(n32784), .QN(n720)
         );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n7993), .CK(CLK), .Q(n32785), .QN(n721)
         );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n7994), .CK(CLK), .Q(n32786), .QN(n722)
         );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n7995), .CK(CLK), .Q(n32787), .QN(n723)
         );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n7996), .CK(CLK), .Q(n32788), .QN(n724)
         );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n7997), .CK(CLK), .Q(n32789), .QN(n725)
         );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n7998), .CK(CLK), .Q(n32790), .QN(n726)
         );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n7999), .CK(CLK), .Q(n32791), .QN(n727)
         );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n8000), .CK(CLK), .Q(n32792), .QN(n728)
         );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n8001), .CK(CLK), .Q(n32793), .QN(n729)
         );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n8002), .CK(CLK), .Q(n32794), .QN(n730)
         );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n8003), .CK(CLK), .Q(n32795), .QN(n731)
         );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n8004), .CK(CLK), .Q(n32796), .QN(n732)
         );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n8005), .CK(CLK), .Q(n32797), .QN(n733)
         );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n8006), .CK(CLK), .Q(n32798), .QN(n734)
         );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n8007), .CK(CLK), .Q(n32799), .QN(n735)
         );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n8008), .CK(CLK), .Q(n32800), .QN(n736)
         );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n8009), .CK(CLK), .Q(n32801), .QN(n737)
         );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n8010), .CK(CLK), .Q(n32802), .QN(n738)
         );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n8011), .CK(CLK), .Q(n32803), .QN(n739)
         );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n8012), .CK(CLK), .Q(n32804), .QN(n740)
         );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n8013), .CK(CLK), .Q(n32805), .QN(n741)
         );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n8014), .CK(CLK), .Q(n32806), .QN(n742)
         );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n8015), .CK(CLK), .Q(n32807), .QN(n743)
         );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n8016), .CK(CLK), .Q(n32808), .QN(n744)
         );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n8017), .CK(CLK), .Q(n32809), .QN(n745)
         );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n8018), .CK(CLK), .Q(n32810), .QN(n746)
         );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n8019), .CK(CLK), .Q(n32811), .QN(n747)
         );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n8020), .CK(CLK), .Q(n32812), .QN(n748)
         );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n8021), .CK(CLK), .Q(n32813), .QN(n749)
         );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n8022), .CK(CLK), .Q(n32814), .QN(n750)
         );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n8023), .CK(CLK), .Q(n32815), .QN(n751)
         );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n8024), .CK(CLK), .Q(n32816), .QN(n752)
         );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n8025), .CK(CLK), .Q(n32817), .QN(n753)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n8026), .CK(CLK), .Q(n32818), .QN(n754)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n8027), .CK(CLK), .Q(n32819), .QN(n755)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n8028), .CK(CLK), .Q(n32820), .QN(n756)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n8029), .CK(CLK), .Q(n32821), .QN(n757)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n8030), .CK(CLK), .Q(n32822), .QN(n758)
         );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n8035), .CK(CLK), .Q(n32823), .QN(n763)
         );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n8036), .CK(CLK), .Q(n32824), .QN(n764)
         );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n8037), .CK(CLK), .Q(n32825), .QN(n765)
         );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n8038), .CK(CLK), .Q(n32826), .QN(n766)
         );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n8039), .CK(CLK), .Q(n32827), .QN(n767)
         );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n8040), .CK(CLK), .Q(n32828), .QN(n768)
         );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n8041), .CK(CLK), .Q(n32829), .QN(n769)
         );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n8042), .CK(CLK), .Q(n32830), .QN(n770)
         );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n8043), .CK(CLK), .Q(n32831), .QN(n771)
         );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n8044), .CK(CLK), .Q(n32832), .QN(n772)
         );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n8045), .CK(CLK), .Q(n32833), .QN(n773)
         );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n8046), .CK(CLK), .Q(n32834), .QN(n774)
         );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n7971), .CK(CLK), .Q(n32835), .QN(n699)
         );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n7972), .CK(CLK), .Q(n32836), .QN(n700)
         );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n7973), .CK(CLK), .Q(n32837), .QN(n701)
         );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n7974), .CK(CLK), .Q(n32838), .QN(n702)
         );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n7975), .CK(CLK), .Q(n32839), .QN(n703)
         );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n7976), .CK(CLK), .Q(n32840), .QN(n704)
         );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n7977), .CK(CLK), .Q(n32841), .QN(n705)
         );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n7978), .CK(CLK), .Q(n32842), .QN(n706)
         );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n7979), .CK(CLK), .Q(n32843), .QN(n707)
         );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n7980), .CK(CLK), .Q(n32844), .QN(n708)
         );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n7981), .CK(CLK), .Q(n32845), .QN(n709)
         );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n7982), .CK(CLK), .Q(n32846), .QN(n710)
         );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n8303), .CK(CLK), .Q(n31069), .QN(n25449) );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n8304), .CK(CLK), .Q(n31070), .QN(n25448) );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n8305), .CK(CLK), .Q(n31071), .QN(n25447) );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n8306), .CK(CLK), .Q(n31072), .QN(n25446) );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n8307), .CK(CLK), .Q(n31073), .QN(n25445) );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n8308), .CK(CLK), .Q(n31074), .QN(n25444) );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n8309), .CK(CLK), .Q(n31075), .QN(n25443) );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n8310), .CK(CLK), .Q(n31076), .QN(n25442) );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n8311), .CK(CLK), .Q(n31077), .QN(n25441) );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n8312), .CK(CLK), .Q(n31078), .QN(n25440) );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n8313), .CK(CLK), .Q(n31079), .QN(n25439) );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n8314), .CK(CLK), .Q(n31080), .QN(n25438) );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n8315), .CK(CLK), .Q(n31081), .QN(n25437) );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n8316), .CK(CLK), .Q(n31082), .QN(n25436) );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n8317), .CK(CLK), .Q(n31083), .QN(n25435) );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n8318), .CK(CLK), .Q(n31084), .QN(n25434) );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n8319), .CK(CLK), .Q(n31085), .QN(n25433) );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n8320), .CK(CLK), .Q(n31086), .QN(n25432) );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n8321), .CK(CLK), .Q(n31087), .QN(n25431) );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n8322), .CK(CLK), .Q(n31088), .QN(n25430) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n8323), .CK(CLK), .Q(n31089), .QN(n25429) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n8324), .CK(CLK), .Q(n31090), .QN(n25428) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n8325), .CK(CLK), .Q(n31091), .QN(n25427) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n8326), .CK(CLK), .Q(n31092), .QN(n25426) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n8327), .CK(CLK), .Q(n31093), .QN(n25425) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n8328), .CK(CLK), .Q(n31094), .QN(n25424) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n8329), .CK(CLK), .Q(n31095), .QN(n25423) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n8330), .CK(CLK), .Q(n31096), .QN(n25422) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n8331), .CK(CLK), .Q(n31097), .QN(n25421) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n8332), .CK(CLK), .Q(n31098), .QN(n25420) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n8333), .CK(CLK), .Q(n31099), .QN(n25419) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n8334), .CK(CLK), .Q(n31100), .QN(n25418) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n8335), .CK(CLK), .Q(n31101), .QN(n25417) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n8336), .CK(CLK), .Q(n31102), .QN(n25416) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n8337), .CK(CLK), .Q(n31103), .QN(n25415) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n8338), .CK(CLK), .Q(n31104), .QN(n25414) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n8339), .CK(CLK), .Q(n31105), .QN(n25413) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n8340), .CK(CLK), .Q(n31106), .QN(n25412) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n8341), .CK(CLK), .Q(n31107), .QN(n25411) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n8342), .CK(CLK), .Q(n31108), .QN(n25410) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n8343), .CK(CLK), .Q(n31109), .QN(n25409) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n8344), .CK(CLK), .Q(n31110), .QN(n25408) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n8345), .CK(CLK), .Q(n31111), .QN(n25407)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n8346), .CK(CLK), .Q(n31112), .QN(n25406)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n8347), .CK(CLK), .Q(n31113), .QN(n25405)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n8348), .CK(CLK), .Q(n31114), .QN(n25404)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n8349), .CK(CLK), .Q(n31115), .QN(n25403)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n8350), .CK(CLK), .Q(n31116), .QN(n25402)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n8291), .CK(CLK), .Q(n31057), .QN(n25397) );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n8292), .CK(CLK), .Q(n31058), .QN(n25396) );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n8293), .CK(CLK), .Q(n31059), .QN(n25395) );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n8294), .CK(CLK), .Q(n31060), .QN(n25457) );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n8295), .CK(CLK), .Q(n31061), .QN(n28840) );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n8296), .CK(CLK), .Q(n31062), .QN(n25456) );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n8297), .CK(CLK), .Q(n31063), .QN(n25455) );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n8298), .CK(CLK), .Q(n31064), .QN(n25454) );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n8299), .CK(CLK), .Q(n31065), .QN(n25453) );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n8300), .CK(CLK), .Q(n31066), .QN(n25452) );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n8301), .CK(CLK), .Q(n31067), .QN(n25451) );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n8302), .CK(CLK), .Q(n31068), .QN(n25450) );
  NOR3_X1 U26462 ( .A1(n32243), .A2(N690), .A3(n37226), .ZN(n37249) );
  NOR3_X1 U26463 ( .A1(N6272), .A2(N6273), .A3(n34672), .ZN(n34693) );
  NOR3_X1 U26464 ( .A1(N6397), .A2(N6398), .A3(n35946), .ZN(n35967) );
  XNOR2_X1 U26465 ( .A(n37251), .B(n32244), .ZN(n37226) );
  XNOR2_X1 U26466 ( .A(n34697), .B(\r504/carry[5] ), .ZN(n34672) );
  XNOR2_X1 U26467 ( .A(n35971), .B(\r510/carry[5] ), .ZN(n35946) );
  XNOR2_X1 U26468 ( .A(n32255), .B(n2699), .ZN(n33398) );
  BUF_X1 U26469 ( .A(n36016), .Z(n39163) );
  BUF_X1 U26470 ( .A(n36016), .Z(n39164) );
  BUF_X1 U26471 ( .A(n36016), .Z(n39165) );
  BUF_X1 U26472 ( .A(n36016), .Z(n39162) );
  BUF_X1 U26473 ( .A(n36016), .Z(n39166) );
  BUF_X1 U26474 ( .A(n39913), .Z(n39914) );
  BUF_X1 U26475 ( .A(n39932), .Z(n39933) );
  BUF_X1 U26476 ( .A(n39913), .Z(n39918) );
  BUF_X1 U26477 ( .A(n39913), .Z(n39917) );
  BUF_X1 U26478 ( .A(n39913), .Z(n39916) );
  BUF_X1 U26479 ( .A(n39913), .Z(n39915) );
  BUF_X1 U26480 ( .A(n39932), .Z(n39937) );
  BUF_X1 U26481 ( .A(n39932), .Z(n39936) );
  BUF_X1 U26482 ( .A(n39932), .Z(n39935) );
  BUF_X1 U26483 ( .A(n39932), .Z(n39934) );
  BUF_X1 U26484 ( .A(n39952), .Z(n39957) );
  BUF_X1 U26485 ( .A(n39952), .Z(n39956) );
  BUF_X1 U26486 ( .A(n39952), .Z(n39955) );
  BUF_X1 U26487 ( .A(n39952), .Z(n39954) );
  BUF_X1 U26488 ( .A(n39952), .Z(n39953) );
  BUF_X1 U26489 ( .A(n39894), .Z(n39899) );
  BUF_X1 U26490 ( .A(n39894), .Z(n39898) );
  BUF_X1 U26491 ( .A(n39894), .Z(n39897) );
  BUF_X1 U26492 ( .A(n39894), .Z(n39896) );
  BUF_X1 U26493 ( .A(n39894), .Z(n39895) );
  BUF_X1 U26494 ( .A(n36028), .Z(n39103) );
  BUF_X1 U26495 ( .A(n36034), .Z(n39073) );
  BUF_X1 U26496 ( .A(n36028), .Z(n39104) );
  BUF_X1 U26497 ( .A(n36034), .Z(n39074) );
  BUF_X1 U26498 ( .A(n36028), .Z(n39105) );
  BUF_X1 U26499 ( .A(n36034), .Z(n39075) );
  BUF_X1 U26500 ( .A(n36028), .Z(n39102) );
  BUF_X1 U26501 ( .A(n36034), .Z(n39072) );
  BUF_X1 U26502 ( .A(n36028), .Z(n39106) );
  BUF_X1 U26503 ( .A(n36034), .Z(n39076) );
  BUF_X1 U26504 ( .A(n33473), .Z(n39608) );
  BUF_X1 U26505 ( .A(n33479), .Z(n39578) );
  BUF_X1 U26506 ( .A(n34747), .Z(n39356) );
  BUF_X1 U26507 ( .A(n34753), .Z(n39326) );
  BUF_X1 U26508 ( .A(n33473), .Z(n39607) );
  BUF_X1 U26509 ( .A(n33479), .Z(n39577) );
  BUF_X1 U26510 ( .A(n34747), .Z(n39355) );
  BUF_X1 U26511 ( .A(n34753), .Z(n39325) );
  BUF_X1 U26512 ( .A(n33473), .Z(n39606) );
  BUF_X1 U26513 ( .A(n33479), .Z(n39576) );
  BUF_X1 U26514 ( .A(n34747), .Z(n39354) );
  BUF_X1 U26515 ( .A(n34753), .Z(n39324) );
  BUF_X1 U26516 ( .A(n33473), .Z(n39605) );
  BUF_X1 U26517 ( .A(n33479), .Z(n39575) );
  BUF_X1 U26518 ( .A(n34747), .Z(n39353) );
  BUF_X1 U26519 ( .A(n34753), .Z(n39323) );
  BUF_X1 U26520 ( .A(n33473), .Z(n39604) );
  BUF_X1 U26521 ( .A(n33479), .Z(n39574) );
  BUF_X1 U26522 ( .A(n34747), .Z(n39352) );
  BUF_X1 U26523 ( .A(n34753), .Z(n39322) );
  BUF_X1 U26524 ( .A(n36022), .Z(n39133) );
  BUF_X1 U26525 ( .A(n36006), .Z(n39193) );
  BUF_X1 U26526 ( .A(n36000), .Z(n39223) );
  BUF_X1 U26527 ( .A(n35988), .Z(n39283) );
  BUF_X1 U26528 ( .A(n35994), .Z(n39253) );
  BUF_X1 U26529 ( .A(n36022), .Z(n39134) );
  BUF_X1 U26530 ( .A(n36006), .Z(n39194) );
  BUF_X1 U26531 ( .A(n36000), .Z(n39224) );
  BUF_X1 U26532 ( .A(n35988), .Z(n39284) );
  BUF_X1 U26533 ( .A(n35994), .Z(n39254) );
  BUF_X1 U26534 ( .A(n36022), .Z(n39135) );
  BUF_X1 U26535 ( .A(n36006), .Z(n39195) );
  BUF_X1 U26536 ( .A(n36000), .Z(n39225) );
  BUF_X1 U26537 ( .A(n35988), .Z(n39285) );
  BUF_X1 U26538 ( .A(n35994), .Z(n39255) );
  BUF_X1 U26539 ( .A(n36022), .Z(n39132) );
  BUF_X1 U26540 ( .A(n36006), .Z(n39192) );
  BUF_X1 U26541 ( .A(n36000), .Z(n39222) );
  BUF_X1 U26542 ( .A(n35988), .Z(n39282) );
  BUF_X1 U26543 ( .A(n35994), .Z(n39252) );
  BUF_X1 U26544 ( .A(n36022), .Z(n39136) );
  BUF_X1 U26545 ( .A(n36006), .Z(n39196) );
  BUF_X1 U26546 ( .A(n36000), .Z(n39226) );
  BUF_X1 U26547 ( .A(n35988), .Z(n39286) );
  BUF_X1 U26548 ( .A(n35994), .Z(n39256) );
  BUF_X1 U26549 ( .A(n33467), .Z(n39638) );
  BUF_X1 U26550 ( .A(n33461), .Z(n39668) );
  BUF_X1 U26551 ( .A(n33433), .Z(n39788) );
  BUF_X1 U26552 ( .A(n33439), .Z(n39758) );
  BUF_X1 U26553 ( .A(n33445), .Z(n39728) );
  BUF_X1 U26554 ( .A(n33451), .Z(n39698) );
  BUF_X1 U26555 ( .A(n34741), .Z(n39386) );
  BUF_X1 U26556 ( .A(n34735), .Z(n39416) );
  BUF_X1 U26557 ( .A(n34707), .Z(n39536) );
  BUF_X1 U26558 ( .A(n34713), .Z(n39506) );
  BUF_X1 U26559 ( .A(n34719), .Z(n39476) );
  BUF_X1 U26560 ( .A(n34725), .Z(n39446) );
  BUF_X1 U26561 ( .A(n33467), .Z(n39637) );
  BUF_X1 U26562 ( .A(n33461), .Z(n39667) );
  BUF_X1 U26563 ( .A(n33433), .Z(n39787) );
  BUF_X1 U26564 ( .A(n33439), .Z(n39757) );
  BUF_X1 U26565 ( .A(n33445), .Z(n39727) );
  BUF_X1 U26566 ( .A(n33451), .Z(n39697) );
  BUF_X1 U26567 ( .A(n34741), .Z(n39385) );
  BUF_X1 U26568 ( .A(n34735), .Z(n39415) );
  BUF_X1 U26569 ( .A(n34707), .Z(n39535) );
  BUF_X1 U26570 ( .A(n34713), .Z(n39505) );
  BUF_X1 U26571 ( .A(n34719), .Z(n39475) );
  BUF_X1 U26572 ( .A(n34725), .Z(n39445) );
  BUF_X1 U26573 ( .A(n33467), .Z(n39636) );
  BUF_X1 U26574 ( .A(n33461), .Z(n39666) );
  BUF_X1 U26575 ( .A(n33433), .Z(n39786) );
  BUF_X1 U26576 ( .A(n33439), .Z(n39756) );
  BUF_X1 U26577 ( .A(n33445), .Z(n39726) );
  BUF_X1 U26578 ( .A(n33451), .Z(n39696) );
  BUF_X1 U26579 ( .A(n34741), .Z(n39384) );
  BUF_X1 U26580 ( .A(n34735), .Z(n39414) );
  BUF_X1 U26581 ( .A(n34707), .Z(n39534) );
  BUF_X1 U26582 ( .A(n34713), .Z(n39504) );
  BUF_X1 U26583 ( .A(n34719), .Z(n39474) );
  BUF_X1 U26584 ( .A(n34725), .Z(n39444) );
  BUF_X1 U26585 ( .A(n33467), .Z(n39635) );
  BUF_X1 U26586 ( .A(n33461), .Z(n39665) );
  BUF_X1 U26587 ( .A(n33433), .Z(n39785) );
  BUF_X1 U26588 ( .A(n33439), .Z(n39755) );
  BUF_X1 U26589 ( .A(n33445), .Z(n39725) );
  BUF_X1 U26590 ( .A(n33451), .Z(n39695) );
  BUF_X1 U26591 ( .A(n34741), .Z(n39383) );
  BUF_X1 U26592 ( .A(n34735), .Z(n39413) );
  BUF_X1 U26593 ( .A(n34707), .Z(n39533) );
  BUF_X1 U26594 ( .A(n34713), .Z(n39503) );
  BUF_X1 U26595 ( .A(n34719), .Z(n39473) );
  BUF_X1 U26596 ( .A(n34725), .Z(n39443) );
  BUF_X1 U26597 ( .A(n33467), .Z(n39634) );
  BUF_X1 U26598 ( .A(n33461), .Z(n39664) );
  BUF_X1 U26599 ( .A(n33433), .Z(n39784) );
  BUF_X1 U26600 ( .A(n33439), .Z(n39754) );
  BUF_X1 U26601 ( .A(n33445), .Z(n39724) );
  BUF_X1 U26602 ( .A(n33451), .Z(n39694) );
  BUF_X1 U26603 ( .A(n34741), .Z(n39382) );
  BUF_X1 U26604 ( .A(n34735), .Z(n39412) );
  BUF_X1 U26605 ( .A(n34707), .Z(n39532) );
  BUF_X1 U26606 ( .A(n34713), .Z(n39502) );
  BUF_X1 U26607 ( .A(n34719), .Z(n39472) );
  BUF_X1 U26608 ( .A(n34725), .Z(n39442) );
  BUF_X1 U26609 ( .A(n36029), .Z(n39097) );
  BUF_X1 U26610 ( .A(n36035), .Z(n39067) );
  BUF_X1 U26611 ( .A(n36029), .Z(n39098) );
  BUF_X1 U26612 ( .A(n36035), .Z(n39068) );
  BUF_X1 U26613 ( .A(n36029), .Z(n39099) );
  BUF_X1 U26614 ( .A(n36035), .Z(n39069) );
  BUF_X1 U26615 ( .A(n36029), .Z(n39096) );
  BUF_X1 U26616 ( .A(n36035), .Z(n39066) );
  BUF_X1 U26617 ( .A(n36029), .Z(n39100) );
  BUF_X1 U26618 ( .A(n36035), .Z(n39070) );
  BUF_X1 U26619 ( .A(n33474), .Z(n39602) );
  BUF_X1 U26620 ( .A(n33480), .Z(n39572) );
  BUF_X1 U26621 ( .A(n34748), .Z(n39350) );
  BUF_X1 U26622 ( .A(n34754), .Z(n39320) );
  BUF_X1 U26623 ( .A(n33474), .Z(n39601) );
  BUF_X1 U26624 ( .A(n33480), .Z(n39571) );
  BUF_X1 U26625 ( .A(n34748), .Z(n39349) );
  BUF_X1 U26626 ( .A(n34754), .Z(n39319) );
  BUF_X1 U26627 ( .A(n33474), .Z(n39600) );
  BUF_X1 U26628 ( .A(n33480), .Z(n39570) );
  BUF_X1 U26629 ( .A(n34748), .Z(n39348) );
  BUF_X1 U26630 ( .A(n34754), .Z(n39318) );
  BUF_X1 U26631 ( .A(n33474), .Z(n39599) );
  BUF_X1 U26632 ( .A(n33480), .Z(n39569) );
  BUF_X1 U26633 ( .A(n34748), .Z(n39347) );
  BUF_X1 U26634 ( .A(n34754), .Z(n39317) );
  BUF_X1 U26635 ( .A(n33474), .Z(n39598) );
  BUF_X1 U26636 ( .A(n33480), .Z(n39568) );
  BUF_X1 U26637 ( .A(n34748), .Z(n39346) );
  BUF_X1 U26638 ( .A(n34754), .Z(n39316) );
  BUF_X1 U26639 ( .A(n36023), .Z(n39127) );
  BUF_X1 U26640 ( .A(n36017), .Z(n39157) );
  BUF_X1 U26641 ( .A(n36007), .Z(n39187) );
  BUF_X1 U26642 ( .A(n36001), .Z(n39217) );
  BUF_X1 U26643 ( .A(n35989), .Z(n39277) );
  BUF_X1 U26644 ( .A(n35995), .Z(n39247) );
  BUF_X1 U26645 ( .A(n36023), .Z(n39128) );
  BUF_X1 U26646 ( .A(n36017), .Z(n39158) );
  BUF_X1 U26647 ( .A(n36007), .Z(n39188) );
  BUF_X1 U26648 ( .A(n36001), .Z(n39218) );
  BUF_X1 U26649 ( .A(n35989), .Z(n39278) );
  BUF_X1 U26650 ( .A(n35995), .Z(n39248) );
  BUF_X1 U26651 ( .A(n36023), .Z(n39129) );
  BUF_X1 U26652 ( .A(n36017), .Z(n39159) );
  BUF_X1 U26653 ( .A(n36007), .Z(n39189) );
  BUF_X1 U26654 ( .A(n36001), .Z(n39219) );
  BUF_X1 U26655 ( .A(n35989), .Z(n39279) );
  BUF_X1 U26656 ( .A(n35995), .Z(n39249) );
  BUF_X1 U26657 ( .A(n36023), .Z(n39126) );
  BUF_X1 U26658 ( .A(n36017), .Z(n39156) );
  BUF_X1 U26659 ( .A(n36007), .Z(n39186) );
  BUF_X1 U26660 ( .A(n36001), .Z(n39216) );
  BUF_X1 U26661 ( .A(n35989), .Z(n39276) );
  BUF_X1 U26662 ( .A(n35995), .Z(n39246) );
  BUF_X1 U26663 ( .A(n36023), .Z(n39130) );
  BUF_X1 U26664 ( .A(n36017), .Z(n39160) );
  BUF_X1 U26665 ( .A(n36007), .Z(n39190) );
  BUF_X1 U26666 ( .A(n36001), .Z(n39220) );
  BUF_X1 U26667 ( .A(n35989), .Z(n39280) );
  BUF_X1 U26668 ( .A(n35995), .Z(n39250) );
  BUF_X1 U26669 ( .A(n33468), .Z(n39632) );
  BUF_X1 U26670 ( .A(n33462), .Z(n39662) );
  BUF_X1 U26671 ( .A(n33434), .Z(n39782) );
  BUF_X1 U26672 ( .A(n33440), .Z(n39752) );
  BUF_X1 U26673 ( .A(n33446), .Z(n39722) );
  BUF_X1 U26674 ( .A(n33452), .Z(n39692) );
  BUF_X1 U26675 ( .A(n34742), .Z(n39380) );
  BUF_X1 U26676 ( .A(n34736), .Z(n39410) );
  BUF_X1 U26677 ( .A(n34708), .Z(n39530) );
  BUF_X1 U26678 ( .A(n34714), .Z(n39500) );
  BUF_X1 U26679 ( .A(n34720), .Z(n39470) );
  BUF_X1 U26680 ( .A(n34726), .Z(n39440) );
  BUF_X1 U26681 ( .A(n33468), .Z(n39631) );
  BUF_X1 U26682 ( .A(n33462), .Z(n39661) );
  BUF_X1 U26683 ( .A(n33434), .Z(n39781) );
  BUF_X1 U26684 ( .A(n33440), .Z(n39751) );
  BUF_X1 U26685 ( .A(n33446), .Z(n39721) );
  BUF_X1 U26686 ( .A(n33452), .Z(n39691) );
  BUF_X1 U26687 ( .A(n34742), .Z(n39379) );
  BUF_X1 U26688 ( .A(n34736), .Z(n39409) );
  BUF_X1 U26689 ( .A(n34708), .Z(n39529) );
  BUF_X1 U26690 ( .A(n34714), .Z(n39499) );
  BUF_X1 U26691 ( .A(n34720), .Z(n39469) );
  BUF_X1 U26692 ( .A(n34726), .Z(n39439) );
  BUF_X1 U26693 ( .A(n33468), .Z(n39630) );
  BUF_X1 U26694 ( .A(n33462), .Z(n39660) );
  BUF_X1 U26695 ( .A(n33434), .Z(n39780) );
  BUF_X1 U26696 ( .A(n33440), .Z(n39750) );
  BUF_X1 U26697 ( .A(n33446), .Z(n39720) );
  BUF_X1 U26698 ( .A(n33452), .Z(n39690) );
  BUF_X1 U26699 ( .A(n34742), .Z(n39378) );
  BUF_X1 U26700 ( .A(n34736), .Z(n39408) );
  BUF_X1 U26701 ( .A(n34708), .Z(n39528) );
  BUF_X1 U26702 ( .A(n34714), .Z(n39498) );
  BUF_X1 U26703 ( .A(n34720), .Z(n39468) );
  BUF_X1 U26704 ( .A(n34726), .Z(n39438) );
  BUF_X1 U26705 ( .A(n33468), .Z(n39629) );
  BUF_X1 U26706 ( .A(n33462), .Z(n39659) );
  BUF_X1 U26707 ( .A(n33434), .Z(n39779) );
  BUF_X1 U26708 ( .A(n33440), .Z(n39749) );
  BUF_X1 U26709 ( .A(n33446), .Z(n39719) );
  BUF_X1 U26710 ( .A(n33452), .Z(n39689) );
  BUF_X1 U26711 ( .A(n34742), .Z(n39377) );
  BUF_X1 U26712 ( .A(n34736), .Z(n39407) );
  BUF_X1 U26713 ( .A(n34708), .Z(n39527) );
  BUF_X1 U26714 ( .A(n34714), .Z(n39497) );
  BUF_X1 U26715 ( .A(n34720), .Z(n39467) );
  BUF_X1 U26716 ( .A(n34726), .Z(n39437) );
  BUF_X1 U26717 ( .A(n33468), .Z(n39628) );
  BUF_X1 U26718 ( .A(n33462), .Z(n39658) );
  BUF_X1 U26719 ( .A(n33434), .Z(n39778) );
  BUF_X1 U26720 ( .A(n33440), .Z(n39748) );
  BUF_X1 U26721 ( .A(n33446), .Z(n39718) );
  BUF_X1 U26722 ( .A(n33452), .Z(n39688) );
  BUF_X1 U26723 ( .A(n34742), .Z(n39376) );
  BUF_X1 U26724 ( .A(n34736), .Z(n39406) );
  BUF_X1 U26725 ( .A(n34708), .Z(n39526) );
  BUF_X1 U26726 ( .A(n34714), .Z(n39496) );
  BUF_X1 U26727 ( .A(n34720), .Z(n39466) );
  BUF_X1 U26728 ( .A(n34726), .Z(n39436) );
  BUF_X1 U26729 ( .A(n33438), .Z(n39764) );
  BUF_X1 U26730 ( .A(n33444), .Z(n39734) );
  BUF_X1 U26731 ( .A(n34712), .Z(n39512) );
  BUF_X1 U26732 ( .A(n34718), .Z(n39482) );
  BUF_X1 U26733 ( .A(n33438), .Z(n39763) );
  BUF_X1 U26734 ( .A(n33444), .Z(n39733) );
  BUF_X1 U26735 ( .A(n34712), .Z(n39511) );
  BUF_X1 U26736 ( .A(n34718), .Z(n39481) );
  BUF_X1 U26737 ( .A(n33438), .Z(n39762) );
  BUF_X1 U26738 ( .A(n33444), .Z(n39732) );
  BUF_X1 U26739 ( .A(n34712), .Z(n39510) );
  BUF_X1 U26740 ( .A(n34718), .Z(n39480) );
  BUF_X1 U26741 ( .A(n33438), .Z(n39761) );
  BUF_X1 U26742 ( .A(n33444), .Z(n39731) );
  BUF_X1 U26743 ( .A(n34712), .Z(n39509) );
  BUF_X1 U26744 ( .A(n34718), .Z(n39479) );
  BUF_X1 U26745 ( .A(n33438), .Z(n39760) );
  BUF_X1 U26746 ( .A(n33444), .Z(n39730) );
  BUF_X1 U26747 ( .A(n34712), .Z(n39508) );
  BUF_X1 U26748 ( .A(n34718), .Z(n39478) );
  BUF_X1 U26749 ( .A(n35993), .Z(n39259) );
  BUF_X1 U26750 ( .A(n35999), .Z(n39229) );
  BUF_X1 U26751 ( .A(n35993), .Z(n39260) );
  BUF_X1 U26752 ( .A(n35999), .Z(n39230) );
  BUF_X1 U26753 ( .A(n35993), .Z(n39261) );
  BUF_X1 U26754 ( .A(n35999), .Z(n39231) );
  BUF_X1 U26755 ( .A(n35993), .Z(n39258) );
  BUF_X1 U26756 ( .A(n35999), .Z(n39228) );
  BUF_X1 U26757 ( .A(n35993), .Z(n39262) );
  BUF_X1 U26758 ( .A(n35999), .Z(n39232) );
  BUF_X1 U26759 ( .A(n33478), .Z(n39584) );
  BUF_X1 U26760 ( .A(n33450), .Z(n39704) );
  BUF_X1 U26761 ( .A(n34752), .Z(n39332) );
  BUF_X1 U26762 ( .A(n34724), .Z(n39452) );
  BUF_X1 U26763 ( .A(n33478), .Z(n39583) );
  BUF_X1 U26764 ( .A(n33450), .Z(n39703) );
  BUF_X1 U26765 ( .A(n34752), .Z(n39331) );
  BUF_X1 U26766 ( .A(n34724), .Z(n39451) );
  BUF_X1 U26767 ( .A(n33478), .Z(n39582) );
  BUF_X1 U26768 ( .A(n33450), .Z(n39702) );
  BUF_X1 U26769 ( .A(n34752), .Z(n39330) );
  BUF_X1 U26770 ( .A(n34724), .Z(n39450) );
  BUF_X1 U26771 ( .A(n33478), .Z(n39581) );
  BUF_X1 U26772 ( .A(n33450), .Z(n39701) );
  BUF_X1 U26773 ( .A(n34752), .Z(n39329) );
  BUF_X1 U26774 ( .A(n34724), .Z(n39449) );
  BUF_X1 U26775 ( .A(n33478), .Z(n39580) );
  BUF_X1 U26776 ( .A(n33450), .Z(n39700) );
  BUF_X1 U26777 ( .A(n34752), .Z(n39328) );
  BUF_X1 U26778 ( .A(n34724), .Z(n39448) );
  BUF_X1 U26779 ( .A(n33484), .Z(n39554) );
  BUF_X1 U26780 ( .A(n33484), .Z(n39553) );
  BUF_X1 U26781 ( .A(n36033), .Z(n39079) );
  BUF_X1 U26782 ( .A(n36039), .Z(n39049) );
  BUF_X1 U26783 ( .A(n36021), .Z(n39139) );
  BUF_X1 U26784 ( .A(n36011), .Z(n39169) );
  BUF_X1 U26785 ( .A(n36033), .Z(n39080) );
  BUF_X1 U26786 ( .A(n36039), .Z(n39050) );
  BUF_X1 U26787 ( .A(n36021), .Z(n39140) );
  BUF_X1 U26788 ( .A(n36011), .Z(n39170) );
  BUF_X1 U26789 ( .A(n36033), .Z(n39081) );
  BUF_X1 U26790 ( .A(n36039), .Z(n39051) );
  BUF_X1 U26791 ( .A(n36021), .Z(n39141) );
  BUF_X1 U26792 ( .A(n36011), .Z(n39171) );
  BUF_X1 U26793 ( .A(n36033), .Z(n39078) );
  BUF_X1 U26794 ( .A(n36039), .Z(n39048) );
  BUF_X1 U26795 ( .A(n36021), .Z(n39138) );
  BUF_X1 U26796 ( .A(n36011), .Z(n39168) );
  BUF_X1 U26797 ( .A(n36033), .Z(n39082) );
  BUF_X1 U26798 ( .A(n36039), .Z(n39052) );
  BUF_X1 U26799 ( .A(n36021), .Z(n39142) );
  BUF_X1 U26800 ( .A(n36011), .Z(n39172) );
  BUF_X1 U26801 ( .A(n33466), .Z(n39644) );
  BUF_X1 U26802 ( .A(n34758), .Z(n39302) );
  BUF_X1 U26803 ( .A(n34740), .Z(n39392) );
  BUF_X1 U26804 ( .A(n33466), .Z(n39643) );
  BUF_X1 U26805 ( .A(n34758), .Z(n39301) );
  BUF_X1 U26806 ( .A(n34740), .Z(n39391) );
  BUF_X1 U26807 ( .A(n33484), .Z(n39552) );
  BUF_X1 U26808 ( .A(n33466), .Z(n39642) );
  BUF_X1 U26809 ( .A(n34758), .Z(n39300) );
  BUF_X1 U26810 ( .A(n34740), .Z(n39390) );
  BUF_X1 U26811 ( .A(n33484), .Z(n39551) );
  BUF_X1 U26812 ( .A(n33466), .Z(n39641) );
  BUF_X1 U26813 ( .A(n34758), .Z(n39299) );
  BUF_X1 U26814 ( .A(n34740), .Z(n39389) );
  BUF_X1 U26815 ( .A(n33484), .Z(n39550) );
  BUF_X1 U26816 ( .A(n33466), .Z(n39640) );
  BUF_X1 U26817 ( .A(n34758), .Z(n39298) );
  BUF_X1 U26818 ( .A(n34740), .Z(n39388) );
  BUF_X1 U26819 ( .A(n36005), .Z(n39199) );
  BUF_X1 U26820 ( .A(n36005), .Z(n39200) );
  BUF_X1 U26821 ( .A(n36005), .Z(n39201) );
  BUF_X1 U26822 ( .A(n36005), .Z(n39198) );
  BUF_X1 U26823 ( .A(n36005), .Z(n39202) );
  BUF_X1 U26824 ( .A(n36027), .Z(n39109) );
  BUF_X1 U26825 ( .A(n36027), .Z(n39110) );
  BUF_X1 U26826 ( .A(n36027), .Z(n39111) );
  BUF_X1 U26827 ( .A(n36027), .Z(n39108) );
  BUF_X1 U26828 ( .A(n36027), .Z(n39112) );
  BUF_X1 U26829 ( .A(n33472), .Z(n39614) );
  BUF_X1 U26830 ( .A(n34746), .Z(n39362) );
  BUF_X1 U26831 ( .A(n33472), .Z(n39613) );
  BUF_X1 U26832 ( .A(n34746), .Z(n39361) );
  BUF_X1 U26833 ( .A(n33472), .Z(n39612) );
  BUF_X1 U26834 ( .A(n34746), .Z(n39360) );
  BUF_X1 U26835 ( .A(n33472), .Z(n39611) );
  BUF_X1 U26836 ( .A(n34746), .Z(n39359) );
  BUF_X1 U26837 ( .A(n33472), .Z(n39610) );
  BUF_X1 U26838 ( .A(n34746), .Z(n39358) );
  BUF_X1 U26839 ( .A(n33456), .Z(n39674) );
  BUF_X1 U26840 ( .A(n34730), .Z(n39422) );
  BUF_X1 U26841 ( .A(n33456), .Z(n39673) );
  BUF_X1 U26842 ( .A(n34730), .Z(n39421) );
  BUF_X1 U26843 ( .A(n33456), .Z(n39672) );
  BUF_X1 U26844 ( .A(n34730), .Z(n39420) );
  BUF_X1 U26845 ( .A(n33456), .Z(n39671) );
  BUF_X1 U26846 ( .A(n34730), .Z(n39419) );
  BUF_X1 U26847 ( .A(n33456), .Z(n39670) );
  BUF_X1 U26848 ( .A(n34730), .Z(n39418) );
  BUF_X1 U26849 ( .A(n33436), .Z(n39776) );
  BUF_X1 U26850 ( .A(n33442), .Z(n39746) );
  BUF_X1 U26851 ( .A(n34710), .Z(n39524) );
  BUF_X1 U26852 ( .A(n34716), .Z(n39494) );
  BUF_X1 U26853 ( .A(n33436), .Z(n39775) );
  BUF_X1 U26854 ( .A(n33442), .Z(n39745) );
  BUF_X1 U26855 ( .A(n34710), .Z(n39523) );
  BUF_X1 U26856 ( .A(n34716), .Z(n39493) );
  BUF_X1 U26857 ( .A(n33436), .Z(n39774) );
  BUF_X1 U26858 ( .A(n33442), .Z(n39744) );
  BUF_X1 U26859 ( .A(n34710), .Z(n39522) );
  BUF_X1 U26860 ( .A(n34716), .Z(n39492) );
  BUF_X1 U26861 ( .A(n33436), .Z(n39773) );
  BUF_X1 U26862 ( .A(n33442), .Z(n39743) );
  BUF_X1 U26863 ( .A(n34710), .Z(n39521) );
  BUF_X1 U26864 ( .A(n34716), .Z(n39491) );
  BUF_X1 U26865 ( .A(n33436), .Z(n39772) );
  BUF_X1 U26866 ( .A(n33442), .Z(n39742) );
  BUF_X1 U26867 ( .A(n34710), .Z(n39520) );
  BUF_X1 U26868 ( .A(n34716), .Z(n39490) );
  BUF_X1 U26869 ( .A(n35991), .Z(n39271) );
  BUF_X1 U26870 ( .A(n35997), .Z(n39241) );
  BUF_X1 U26871 ( .A(n35991), .Z(n39272) );
  BUF_X1 U26872 ( .A(n35997), .Z(n39242) );
  BUF_X1 U26873 ( .A(n35991), .Z(n39273) );
  BUF_X1 U26874 ( .A(n35997), .Z(n39243) );
  BUF_X1 U26875 ( .A(n35991), .Z(n39270) );
  BUF_X1 U26876 ( .A(n35997), .Z(n39240) );
  BUF_X1 U26877 ( .A(n35991), .Z(n39274) );
  BUF_X1 U26878 ( .A(n35997), .Z(n39244) );
  BUF_X1 U26879 ( .A(n33482), .Z(n39566) );
  BUF_X1 U26880 ( .A(n34756), .Z(n39314) );
  BUF_X1 U26881 ( .A(n33482), .Z(n39565) );
  BUF_X1 U26882 ( .A(n34756), .Z(n39313) );
  BUF_X1 U26883 ( .A(n33482), .Z(n39564) );
  BUF_X1 U26884 ( .A(n34756), .Z(n39312) );
  BUF_X1 U26885 ( .A(n33482), .Z(n39563) );
  BUF_X1 U26886 ( .A(n34756), .Z(n39311) );
  BUF_X1 U26887 ( .A(n33482), .Z(n39562) );
  BUF_X1 U26888 ( .A(n34756), .Z(n39310) );
  BUF_X1 U26889 ( .A(n36037), .Z(n39061) );
  BUF_X1 U26890 ( .A(n36019), .Z(n39151) );
  BUF_X1 U26891 ( .A(n36009), .Z(n39181) );
  BUF_X1 U26892 ( .A(n36037), .Z(n39062) );
  BUF_X1 U26893 ( .A(n36019), .Z(n39152) );
  BUF_X1 U26894 ( .A(n36009), .Z(n39182) );
  BUF_X1 U26895 ( .A(n36037), .Z(n39063) );
  BUF_X1 U26896 ( .A(n36019), .Z(n39153) );
  BUF_X1 U26897 ( .A(n36009), .Z(n39183) );
  BUF_X1 U26898 ( .A(n36037), .Z(n39060) );
  BUF_X1 U26899 ( .A(n36019), .Z(n39150) );
  BUF_X1 U26900 ( .A(n36009), .Z(n39180) );
  BUF_X1 U26901 ( .A(n36037), .Z(n39064) );
  BUF_X1 U26902 ( .A(n36019), .Z(n39154) );
  BUF_X1 U26903 ( .A(n36009), .Z(n39184) );
  BUF_X1 U26904 ( .A(n36003), .Z(n39211) );
  BUF_X1 U26905 ( .A(n36003), .Z(n39212) );
  BUF_X1 U26906 ( .A(n36003), .Z(n39213) );
  BUF_X1 U26907 ( .A(n36003), .Z(n39210) );
  BUF_X1 U26908 ( .A(n36003), .Z(n39214) );
  BUF_X1 U26909 ( .A(n33470), .Z(n39626) );
  BUF_X1 U26910 ( .A(n33454), .Z(n39686) );
  BUF_X1 U26911 ( .A(n34744), .Z(n39374) );
  BUF_X1 U26912 ( .A(n34728), .Z(n39434) );
  BUF_X1 U26913 ( .A(n33470), .Z(n39625) );
  BUF_X1 U26914 ( .A(n33454), .Z(n39685) );
  BUF_X1 U26915 ( .A(n34744), .Z(n39373) );
  BUF_X1 U26916 ( .A(n34728), .Z(n39433) );
  BUF_X1 U26917 ( .A(n33470), .Z(n39624) );
  BUF_X1 U26918 ( .A(n33454), .Z(n39684) );
  BUF_X1 U26919 ( .A(n34744), .Z(n39372) );
  BUF_X1 U26920 ( .A(n34728), .Z(n39432) );
  BUF_X1 U26921 ( .A(n33470), .Z(n39623) );
  BUF_X1 U26922 ( .A(n33454), .Z(n39683) );
  BUF_X1 U26923 ( .A(n34744), .Z(n39371) );
  BUF_X1 U26924 ( .A(n34728), .Z(n39431) );
  BUF_X1 U26925 ( .A(n33470), .Z(n39622) );
  BUF_X1 U26926 ( .A(n33454), .Z(n39682) );
  BUF_X1 U26927 ( .A(n34744), .Z(n39370) );
  BUF_X1 U26928 ( .A(n34728), .Z(n39430) );
  BUF_X1 U26929 ( .A(n36031), .Z(n39091) );
  BUF_X1 U26930 ( .A(n36031), .Z(n39092) );
  BUF_X1 U26931 ( .A(n36031), .Z(n39093) );
  BUF_X1 U26932 ( .A(n36031), .Z(n39090) );
  BUF_X1 U26933 ( .A(n36031), .Z(n39094) );
  BUF_X1 U26934 ( .A(n33476), .Z(n39596) );
  BUF_X1 U26935 ( .A(n33448), .Z(n39716) );
  BUF_X1 U26936 ( .A(n34750), .Z(n39344) );
  BUF_X1 U26937 ( .A(n34722), .Z(n39464) );
  BUF_X1 U26938 ( .A(n33476), .Z(n39595) );
  BUF_X1 U26939 ( .A(n33448), .Z(n39715) );
  BUF_X1 U26940 ( .A(n34750), .Z(n39343) );
  BUF_X1 U26941 ( .A(n34722), .Z(n39463) );
  BUF_X1 U26942 ( .A(n33476), .Z(n39594) );
  BUF_X1 U26943 ( .A(n33448), .Z(n39714) );
  BUF_X1 U26944 ( .A(n34750), .Z(n39342) );
  BUF_X1 U26945 ( .A(n34722), .Z(n39462) );
  BUF_X1 U26946 ( .A(n33476), .Z(n39593) );
  BUF_X1 U26947 ( .A(n33448), .Z(n39713) );
  BUF_X1 U26948 ( .A(n34750), .Z(n39341) );
  BUF_X1 U26949 ( .A(n34722), .Z(n39461) );
  BUF_X1 U26950 ( .A(n33476), .Z(n39592) );
  BUF_X1 U26951 ( .A(n33448), .Z(n39712) );
  BUF_X1 U26952 ( .A(n34750), .Z(n39340) );
  BUF_X1 U26953 ( .A(n34722), .Z(n39460) );
  BUF_X1 U26954 ( .A(n33437), .Z(n39770) );
  BUF_X1 U26955 ( .A(n33443), .Z(n39740) );
  BUF_X1 U26956 ( .A(n34711), .Z(n39518) );
  BUF_X1 U26957 ( .A(n34717), .Z(n39488) );
  BUF_X1 U26958 ( .A(n33437), .Z(n39769) );
  BUF_X1 U26959 ( .A(n33443), .Z(n39739) );
  BUF_X1 U26960 ( .A(n34711), .Z(n39517) );
  BUF_X1 U26961 ( .A(n34717), .Z(n39487) );
  BUF_X1 U26962 ( .A(n33437), .Z(n39768) );
  BUF_X1 U26963 ( .A(n33443), .Z(n39738) );
  BUF_X1 U26964 ( .A(n34711), .Z(n39516) );
  BUF_X1 U26965 ( .A(n34717), .Z(n39486) );
  BUF_X1 U26966 ( .A(n33437), .Z(n39767) );
  BUF_X1 U26967 ( .A(n33443), .Z(n39737) );
  BUF_X1 U26968 ( .A(n34711), .Z(n39515) );
  BUF_X1 U26969 ( .A(n34717), .Z(n39485) );
  BUF_X1 U26970 ( .A(n33437), .Z(n39766) );
  BUF_X1 U26971 ( .A(n33443), .Z(n39736) );
  BUF_X1 U26972 ( .A(n34711), .Z(n39514) );
  BUF_X1 U26973 ( .A(n34717), .Z(n39484) );
  BUF_X1 U26974 ( .A(n36025), .Z(n39121) );
  BUF_X1 U26975 ( .A(n36025), .Z(n39122) );
  BUF_X1 U26976 ( .A(n36025), .Z(n39123) );
  BUF_X1 U26977 ( .A(n36025), .Z(n39120) );
  BUF_X1 U26978 ( .A(n36025), .Z(n39124) );
  BUF_X1 U26979 ( .A(n33464), .Z(n39656) );
  BUF_X1 U26980 ( .A(n34738), .Z(n39404) );
  BUF_X1 U26981 ( .A(n33464), .Z(n39655) );
  BUF_X1 U26982 ( .A(n34738), .Z(n39403) );
  BUF_X1 U26983 ( .A(n33464), .Z(n39654) );
  BUF_X1 U26984 ( .A(n34738), .Z(n39402) );
  BUF_X1 U26985 ( .A(n33464), .Z(n39653) );
  BUF_X1 U26986 ( .A(n34738), .Z(n39401) );
  BUF_X1 U26987 ( .A(n33464), .Z(n39652) );
  BUF_X1 U26988 ( .A(n34738), .Z(n39400) );
  BUF_X1 U26989 ( .A(n33477), .Z(n39590) );
  BUF_X1 U26990 ( .A(n34751), .Z(n39338) );
  BUF_X1 U26991 ( .A(n33477), .Z(n39589) );
  BUF_X1 U26992 ( .A(n34751), .Z(n39337) );
  BUF_X1 U26993 ( .A(n33477), .Z(n39588) );
  BUF_X1 U26994 ( .A(n34751), .Z(n39336) );
  BUF_X1 U26995 ( .A(n33477), .Z(n39587) );
  BUF_X1 U26996 ( .A(n34751), .Z(n39335) );
  BUF_X1 U26997 ( .A(n33477), .Z(n39586) );
  BUF_X1 U26998 ( .A(n34751), .Z(n39334) );
  BUF_X1 U26999 ( .A(n35992), .Z(n39265) );
  BUF_X1 U27000 ( .A(n35998), .Z(n39235) );
  BUF_X1 U27001 ( .A(n35992), .Z(n39266) );
  BUF_X1 U27002 ( .A(n35998), .Z(n39236) );
  BUF_X1 U27003 ( .A(n35992), .Z(n39267) );
  BUF_X1 U27004 ( .A(n35998), .Z(n39237) );
  BUF_X1 U27005 ( .A(n35992), .Z(n39264) );
  BUF_X1 U27006 ( .A(n35998), .Z(n39234) );
  BUF_X1 U27007 ( .A(n35992), .Z(n39268) );
  BUF_X1 U27008 ( .A(n35998), .Z(n39238) );
  BUF_X1 U27009 ( .A(n33465), .Z(n39650) );
  BUF_X1 U27010 ( .A(n33449), .Z(n39710) );
  BUF_X1 U27011 ( .A(n34739), .Z(n39398) );
  BUF_X1 U27012 ( .A(n34723), .Z(n39458) );
  BUF_X1 U27013 ( .A(n33465), .Z(n39649) );
  BUF_X1 U27014 ( .A(n33449), .Z(n39709) );
  BUF_X1 U27015 ( .A(n34739), .Z(n39397) );
  BUF_X1 U27016 ( .A(n34723), .Z(n39457) );
  BUF_X1 U27017 ( .A(n33465), .Z(n39648) );
  BUF_X1 U27018 ( .A(n33449), .Z(n39708) );
  BUF_X1 U27019 ( .A(n34739), .Z(n39396) );
  BUF_X1 U27020 ( .A(n34723), .Z(n39456) );
  BUF_X1 U27021 ( .A(n33465), .Z(n39647) );
  BUF_X1 U27022 ( .A(n33449), .Z(n39707) );
  BUF_X1 U27023 ( .A(n34739), .Z(n39395) );
  BUF_X1 U27024 ( .A(n34723), .Z(n39455) );
  BUF_X1 U27025 ( .A(n33465), .Z(n39646) );
  BUF_X1 U27026 ( .A(n33449), .Z(n39706) );
  BUF_X1 U27027 ( .A(n34739), .Z(n39394) );
  BUF_X1 U27028 ( .A(n34723), .Z(n39454) );
  BUF_X1 U27029 ( .A(n33483), .Z(n39560) );
  BUF_X1 U27030 ( .A(n34757), .Z(n39308) );
  BUF_X1 U27031 ( .A(n33483), .Z(n39559) );
  BUF_X1 U27032 ( .A(n34757), .Z(n39307) );
  BUF_X1 U27033 ( .A(n33483), .Z(n39558) );
  BUF_X1 U27034 ( .A(n34757), .Z(n39306) );
  BUF_X1 U27035 ( .A(n33483), .Z(n39557) );
  BUF_X1 U27036 ( .A(n34757), .Z(n39305) );
  BUF_X1 U27037 ( .A(n33483), .Z(n39556) );
  BUF_X1 U27038 ( .A(n34757), .Z(n39304) );
  BUF_X1 U27039 ( .A(n36038), .Z(n39055) );
  BUF_X1 U27040 ( .A(n36010), .Z(n39175) );
  BUF_X1 U27041 ( .A(n36038), .Z(n39056) );
  BUF_X1 U27042 ( .A(n36010), .Z(n39176) );
  BUF_X1 U27043 ( .A(n36038), .Z(n39057) );
  BUF_X1 U27044 ( .A(n36010), .Z(n39177) );
  BUF_X1 U27045 ( .A(n36038), .Z(n39054) );
  BUF_X1 U27046 ( .A(n36010), .Z(n39174) );
  BUF_X1 U27047 ( .A(n36038), .Z(n39058) );
  BUF_X1 U27048 ( .A(n36010), .Z(n39178) );
  BUF_X1 U27049 ( .A(n36020), .Z(n39145) );
  BUF_X1 U27050 ( .A(n36020), .Z(n39146) );
  BUF_X1 U27051 ( .A(n36020), .Z(n39147) );
  BUF_X1 U27052 ( .A(n36020), .Z(n39144) );
  BUF_X1 U27053 ( .A(n36020), .Z(n39148) );
  BUF_X1 U27054 ( .A(n36004), .Z(n39205) );
  BUF_X1 U27055 ( .A(n36004), .Z(n39206) );
  BUF_X1 U27056 ( .A(n36004), .Z(n39207) );
  BUF_X1 U27057 ( .A(n36004), .Z(n39204) );
  BUF_X1 U27058 ( .A(n36004), .Z(n39208) );
  BUF_X1 U27059 ( .A(n36032), .Z(n39085) );
  BUF_X1 U27060 ( .A(n36026), .Z(n39115) );
  BUF_X1 U27061 ( .A(n36032), .Z(n39086) );
  BUF_X1 U27062 ( .A(n36026), .Z(n39116) );
  BUF_X1 U27063 ( .A(n36032), .Z(n39087) );
  BUF_X1 U27064 ( .A(n36026), .Z(n39117) );
  BUF_X1 U27065 ( .A(n36032), .Z(n39084) );
  BUF_X1 U27066 ( .A(n36026), .Z(n39114) );
  BUF_X1 U27067 ( .A(n36032), .Z(n39088) );
  BUF_X1 U27068 ( .A(n36026), .Z(n39118) );
  BUF_X1 U27069 ( .A(n33471), .Z(n39620) );
  BUF_X1 U27070 ( .A(n33455), .Z(n39680) );
  BUF_X1 U27071 ( .A(n34745), .Z(n39368) );
  BUF_X1 U27072 ( .A(n34729), .Z(n39428) );
  BUF_X1 U27073 ( .A(n33471), .Z(n39619) );
  BUF_X1 U27074 ( .A(n33455), .Z(n39679) );
  BUF_X1 U27075 ( .A(n34745), .Z(n39367) );
  BUF_X1 U27076 ( .A(n34729), .Z(n39427) );
  BUF_X1 U27077 ( .A(n33471), .Z(n39618) );
  BUF_X1 U27078 ( .A(n33455), .Z(n39678) );
  BUF_X1 U27079 ( .A(n34745), .Z(n39366) );
  BUF_X1 U27080 ( .A(n34729), .Z(n39426) );
  BUF_X1 U27081 ( .A(n33471), .Z(n39617) );
  BUF_X1 U27082 ( .A(n33455), .Z(n39677) );
  BUF_X1 U27083 ( .A(n34745), .Z(n39365) );
  BUF_X1 U27084 ( .A(n34729), .Z(n39425) );
  BUF_X1 U27085 ( .A(n33471), .Z(n39616) );
  BUF_X1 U27086 ( .A(n33455), .Z(n39676) );
  BUF_X1 U27087 ( .A(n34745), .Z(n39364) );
  BUF_X1 U27088 ( .A(n34729), .Z(n39424) );
  BUF_X1 U27089 ( .A(n33405), .Z(n39901) );
  BUF_X1 U27090 ( .A(n33401), .Z(n39920) );
  BUF_X1 U27091 ( .A(n33384), .Z(n39999) );
  BUF_X1 U27092 ( .A(n33381), .Z(n40018) );
  BUF_X1 U27093 ( .A(n33365), .Z(n40097) );
  BUF_X1 U27094 ( .A(n33420), .Z(n39802) );
  BUF_X1 U27095 ( .A(n33405), .Z(n39904) );
  BUF_X1 U27096 ( .A(n33405), .Z(n39903) );
  BUF_X1 U27097 ( .A(n33405), .Z(n39902) );
  BUF_X1 U27098 ( .A(n33401), .Z(n39923) );
  BUF_X1 U27099 ( .A(n33401), .Z(n39922) );
  BUF_X1 U27100 ( .A(n33401), .Z(n39921) );
  BUF_X1 U27101 ( .A(n33384), .Z(n40002) );
  BUF_X1 U27102 ( .A(n33384), .Z(n40001) );
  BUF_X1 U27103 ( .A(n33384), .Z(n40000) );
  BUF_X1 U27104 ( .A(n33381), .Z(n40021) );
  BUF_X1 U27105 ( .A(n33381), .Z(n40020) );
  BUF_X1 U27106 ( .A(n33381), .Z(n40019) );
  BUF_X1 U27107 ( .A(n33405), .Z(n39905) );
  BUF_X1 U27108 ( .A(n33401), .Z(n39924) );
  BUF_X1 U27109 ( .A(n33384), .Z(n40003) );
  BUF_X1 U27110 ( .A(n33381), .Z(n40022) );
  BUF_X1 U27111 ( .A(n33361), .Z(n40117) );
  BUF_X1 U27112 ( .A(n33361), .Z(n40118) );
  BUF_X1 U27113 ( .A(n33361), .Z(n40119) );
  BUF_X1 U27114 ( .A(n33361), .Z(n40120) );
  BUF_X1 U27115 ( .A(n33365), .Z(n40101) );
  BUF_X1 U27116 ( .A(n33365), .Z(n40100) );
  BUF_X1 U27117 ( .A(n33365), .Z(n40099) );
  BUF_X1 U27118 ( .A(n33365), .Z(n40098) );
  BUF_X1 U27119 ( .A(n33420), .Z(n39804) );
  BUF_X1 U27120 ( .A(n33420), .Z(n39803) );
  BUF_X1 U27121 ( .A(n33420), .Z(n39806) );
  BUF_X1 U27122 ( .A(n33420), .Z(n39805) );
  BUF_X1 U27123 ( .A(n33311), .Z(n40397) );
  BUF_X1 U27124 ( .A(n33311), .Z(n40398) );
  BUF_X1 U27125 ( .A(n33311), .Z(n40399) );
  BUF_X1 U27126 ( .A(n33311), .Z(n40400) );
  BUF_X1 U27127 ( .A(n33349), .Z(n40197) );
  BUF_X1 U27128 ( .A(n33349), .Z(n40198) );
  BUF_X1 U27129 ( .A(n33349), .Z(n40199) );
  BUF_X1 U27130 ( .A(n33349), .Z(n40200) );
  BUF_X1 U27131 ( .A(n33311), .Z(n40396) );
  BUF_X1 U27132 ( .A(n33349), .Z(n40196) );
  BUF_X1 U27133 ( .A(n33317), .Z(n40356) );
  BUF_X1 U27134 ( .A(n33317), .Z(n40357) );
  BUF_X1 U27135 ( .A(n33317), .Z(n40358) );
  BUF_X1 U27136 ( .A(n33317), .Z(n40359) );
  BUF_X1 U27137 ( .A(n33317), .Z(n40360) );
  BUF_X1 U27138 ( .A(n33343), .Z(n40236) );
  BUF_X1 U27139 ( .A(n33343), .Z(n40237) );
  BUF_X1 U27140 ( .A(n33343), .Z(n40238) );
  BUF_X1 U27141 ( .A(n33343), .Z(n40239) );
  BUF_X1 U27142 ( .A(n33343), .Z(n40240) );
  BUF_X1 U27143 ( .A(n33372), .Z(n40077) );
  BUF_X1 U27144 ( .A(n33372), .Z(n40078) );
  BUF_X1 U27145 ( .A(n33372), .Z(n40079) );
  BUF_X1 U27146 ( .A(n33372), .Z(n40080) );
  BUF_X1 U27147 ( .A(n33372), .Z(n40081) );
  BUF_X1 U27148 ( .A(n33378), .Z(n40037) );
  BUF_X1 U27149 ( .A(n33378), .Z(n40038) );
  BUF_X1 U27150 ( .A(n33378), .Z(n40039) );
  BUF_X1 U27151 ( .A(n33378), .Z(n40040) );
  BUF_X1 U27152 ( .A(n33378), .Z(n40041) );
  BUF_X1 U27153 ( .A(n33346), .Z(n40217) );
  BUF_X1 U27154 ( .A(n33346), .Z(n40218) );
  BUF_X1 U27155 ( .A(n33346), .Z(n40219) );
  BUF_X1 U27156 ( .A(n33346), .Z(n40220) );
  BUF_X1 U27157 ( .A(n33346), .Z(n40216) );
  BUF_X1 U27158 ( .A(n33314), .Z(n40376) );
  BUF_X1 U27159 ( .A(n33314), .Z(n40377) );
  BUF_X1 U27160 ( .A(n33314), .Z(n40378) );
  BUF_X1 U27161 ( .A(n33314), .Z(n40379) );
  BUF_X1 U27162 ( .A(n33314), .Z(n40380) );
  BUF_X1 U27163 ( .A(n33375), .Z(n40057) );
  BUF_X1 U27164 ( .A(n33375), .Z(n40058) );
  BUF_X1 U27165 ( .A(n33375), .Z(n40059) );
  BUF_X1 U27166 ( .A(n33375), .Z(n40060) );
  BUF_X1 U27167 ( .A(n33375), .Z(n40061) );
  BUF_X1 U27168 ( .A(n33304), .Z(n40417) );
  BUF_X1 U27169 ( .A(n33304), .Z(n40418) );
  BUF_X1 U27170 ( .A(n33304), .Z(n40419) );
  BUF_X1 U27171 ( .A(n33304), .Z(n40420) );
  BUF_X1 U27172 ( .A(n33326), .Z(n40297) );
  BUF_X1 U27173 ( .A(n33326), .Z(n40298) );
  BUF_X1 U27174 ( .A(n33326), .Z(n40299) );
  BUF_X1 U27175 ( .A(n33326), .Z(n40300) );
  BUF_X1 U27176 ( .A(n33323), .Z(n40317) );
  BUF_X1 U27177 ( .A(n33323), .Z(n40318) );
  BUF_X1 U27178 ( .A(n33323), .Z(n40319) );
  BUF_X1 U27179 ( .A(n33323), .Z(n40320) );
  BUF_X1 U27180 ( .A(n33417), .Z(n39822) );
  BUF_X1 U27181 ( .A(n33417), .Z(n39823) );
  BUF_X1 U27182 ( .A(n33417), .Z(n39824) );
  BUF_X1 U27183 ( .A(n33417), .Z(n39825) );
  BUF_X1 U27184 ( .A(n33304), .Z(n40416) );
  BUF_X1 U27185 ( .A(n33326), .Z(n40296) );
  BUF_X1 U27186 ( .A(n33323), .Z(n40316) );
  BUF_X1 U27187 ( .A(n33417), .Z(n39821) );
  BUF_X1 U27188 ( .A(n33320), .Z(n40336) );
  BUF_X1 U27189 ( .A(n33320), .Z(n40337) );
  BUF_X1 U27190 ( .A(n33320), .Z(n40338) );
  BUF_X1 U27191 ( .A(n33320), .Z(n40339) );
  BUF_X1 U27192 ( .A(n33320), .Z(n40340) );
  BUF_X1 U27193 ( .A(n33329), .Z(n40276) );
  BUF_X1 U27194 ( .A(n33329), .Z(n40277) );
  BUF_X1 U27195 ( .A(n33329), .Z(n40278) );
  BUF_X1 U27196 ( .A(n33329), .Z(n40279) );
  BUF_X1 U27197 ( .A(n33329), .Z(n40280) );
  BUF_X1 U27198 ( .A(n33336), .Z(n40256) );
  BUF_X1 U27199 ( .A(n33336), .Z(n40257) );
  BUF_X1 U27200 ( .A(n33336), .Z(n40258) );
  BUF_X1 U27201 ( .A(n33336), .Z(n40259) );
  BUF_X1 U27202 ( .A(n33336), .Z(n40260) );
  BUF_X1 U27203 ( .A(n33352), .Z(n40176) );
  BUF_X1 U27204 ( .A(n33352), .Z(n40177) );
  BUF_X1 U27205 ( .A(n33352), .Z(n40178) );
  BUF_X1 U27206 ( .A(n33352), .Z(n40179) );
  BUF_X1 U27207 ( .A(n33352), .Z(n40180) );
  BUF_X1 U27208 ( .A(n33355), .Z(n40156) );
  BUF_X1 U27209 ( .A(n33355), .Z(n40157) );
  BUF_X1 U27210 ( .A(n33355), .Z(n40158) );
  BUF_X1 U27211 ( .A(n33355), .Z(n40159) );
  BUF_X1 U27212 ( .A(n33355), .Z(n40160) );
  BUF_X1 U27213 ( .A(n33358), .Z(n40136) );
  BUF_X1 U27214 ( .A(n33358), .Z(n40137) );
  BUF_X1 U27215 ( .A(n33358), .Z(n40138) );
  BUF_X1 U27216 ( .A(n33358), .Z(n40139) );
  BUF_X1 U27217 ( .A(n33358), .Z(n40140) );
  BUF_X1 U27218 ( .A(n33387), .Z(n39979) );
  BUF_X1 U27219 ( .A(n33387), .Z(n39980) );
  BUF_X1 U27220 ( .A(n33387), .Z(n39981) );
  BUF_X1 U27221 ( .A(n33387), .Z(n39982) );
  BUF_X1 U27222 ( .A(n33387), .Z(n39983) );
  BUF_X1 U27223 ( .A(n33390), .Z(n39959) );
  BUF_X1 U27224 ( .A(n33390), .Z(n39960) );
  BUF_X1 U27225 ( .A(n33390), .Z(n39961) );
  BUF_X1 U27226 ( .A(n33390), .Z(n39962) );
  BUF_X1 U27227 ( .A(n33390), .Z(n39963) );
  BUF_X1 U27228 ( .A(n33393), .Z(n39939) );
  BUF_X1 U27229 ( .A(n33393), .Z(n39940) );
  BUF_X1 U27230 ( .A(n33393), .Z(n39941) );
  BUF_X1 U27231 ( .A(n33393), .Z(n39942) );
  BUF_X1 U27232 ( .A(n33393), .Z(n39943) );
  BUF_X1 U27233 ( .A(n33408), .Z(n39881) );
  BUF_X1 U27234 ( .A(n33408), .Z(n39882) );
  BUF_X1 U27235 ( .A(n33408), .Z(n39883) );
  BUF_X1 U27236 ( .A(n33408), .Z(n39884) );
  BUF_X1 U27237 ( .A(n33408), .Z(n39885) );
  BUF_X1 U27238 ( .A(n33411), .Z(n39861) );
  BUF_X1 U27239 ( .A(n33411), .Z(n39862) );
  BUF_X1 U27240 ( .A(n33411), .Z(n39863) );
  BUF_X1 U27241 ( .A(n33411), .Z(n39864) );
  BUF_X1 U27242 ( .A(n33411), .Z(n39865) );
  BUF_X1 U27243 ( .A(n33414), .Z(n39841) );
  BUF_X1 U27244 ( .A(n33414), .Z(n39842) );
  BUF_X1 U27245 ( .A(n33414), .Z(n39843) );
  BUF_X1 U27246 ( .A(n33414), .Z(n39844) );
  BUF_X1 U27247 ( .A(n33414), .Z(n39845) );
  BUF_X1 U27248 ( .A(n33361), .Z(n40116) );
  BUF_X1 U27249 ( .A(n40589), .Z(n40592) );
  BUF_X1 U27250 ( .A(n40589), .Z(n40591) );
  BUF_X1 U27251 ( .A(n40589), .Z(n40594) );
  BUF_X1 U27252 ( .A(n40589), .Z(n40593) );
  BUF_X1 U27253 ( .A(n40589), .Z(n40590) );
  BUF_X1 U27254 ( .A(n40429), .Z(n40430) );
  BUF_X1 U27255 ( .A(n40429), .Z(n40434) );
  BUF_X1 U27256 ( .A(n40429), .Z(n40433) );
  BUF_X1 U27257 ( .A(n40429), .Z(n40432) );
  BUF_X1 U27258 ( .A(n40429), .Z(n40431) );
  BUF_X1 U27259 ( .A(n40409), .Z(n40410) );
  BUF_X1 U27260 ( .A(n40209), .Z(n40210) );
  BUF_X1 U27261 ( .A(n40229), .Z(n40230) );
  BUF_X1 U27262 ( .A(n40409), .Z(n40414) );
  BUF_X1 U27263 ( .A(n40409), .Z(n40413) );
  BUF_X1 U27264 ( .A(n40409), .Z(n40412) );
  BUF_X1 U27265 ( .A(n40409), .Z(n40411) );
  BUF_X1 U27266 ( .A(n40209), .Z(n40214) );
  BUF_X1 U27267 ( .A(n40209), .Z(n40213) );
  BUF_X1 U27268 ( .A(n40209), .Z(n40212) );
  BUF_X1 U27269 ( .A(n40209), .Z(n40211) );
  BUF_X1 U27270 ( .A(n40229), .Z(n40234) );
  BUF_X1 U27271 ( .A(n40229), .Z(n40233) );
  BUF_X1 U27272 ( .A(n40229), .Z(n40232) );
  BUF_X1 U27273 ( .A(n40229), .Z(n40231) );
  BUF_X1 U27274 ( .A(n40011), .Z(n40012) );
  BUF_X1 U27275 ( .A(n40030), .Z(n40031) );
  BUF_X1 U27276 ( .A(n40011), .Z(n40016) );
  BUF_X1 U27277 ( .A(n40011), .Z(n40015) );
  BUF_X1 U27278 ( .A(n40011), .Z(n40014) );
  BUF_X1 U27279 ( .A(n40011), .Z(n40013) );
  BUF_X1 U27280 ( .A(n40030), .Z(n40035) );
  BUF_X1 U27281 ( .A(n40030), .Z(n40034) );
  BUF_X1 U27282 ( .A(n40030), .Z(n40033) );
  BUF_X1 U27283 ( .A(n40030), .Z(n40032) );
  BUF_X1 U27284 ( .A(n40309), .Z(n40310) );
  BUF_X1 U27285 ( .A(n40329), .Z(n40330) );
  BUF_X1 U27286 ( .A(n39834), .Z(n39835) );
  BUF_X1 U27287 ( .A(n40309), .Z(n40314) );
  BUF_X1 U27288 ( .A(n40309), .Z(n40313) );
  BUF_X1 U27289 ( .A(n40309), .Z(n40312) );
  BUF_X1 U27290 ( .A(n40309), .Z(n40311) );
  BUF_X1 U27291 ( .A(n40329), .Z(n40334) );
  BUF_X1 U27292 ( .A(n40329), .Z(n40333) );
  BUF_X1 U27293 ( .A(n40329), .Z(n40332) );
  BUF_X1 U27294 ( .A(n40329), .Z(n40331) );
  BUF_X1 U27295 ( .A(n39834), .Z(n39839) );
  BUF_X1 U27296 ( .A(n39834), .Z(n39838) );
  BUF_X1 U27297 ( .A(n39834), .Z(n39837) );
  BUF_X1 U27298 ( .A(n39834), .Z(n39836) );
  BUF_X1 U27299 ( .A(n39814), .Z(n39817) );
  BUF_X1 U27300 ( .A(n39814), .Z(n39816) );
  BUF_X1 U27301 ( .A(n39814), .Z(n39815) );
  BUF_X1 U27302 ( .A(n40529), .Z(n40530) );
  BUF_X1 U27303 ( .A(n40529), .Z(n40534) );
  BUF_X1 U27304 ( .A(n40529), .Z(n40533) );
  BUF_X1 U27305 ( .A(n40529), .Z(n40532) );
  BUF_X1 U27306 ( .A(n40529), .Z(n40531) );
  BUF_X1 U27307 ( .A(n40509), .Z(n40510) );
  BUF_X1 U27308 ( .A(n40509), .Z(n40514) );
  BUF_X1 U27309 ( .A(n40509), .Z(n40513) );
  BUF_X1 U27310 ( .A(n40509), .Z(n40512) );
  BUF_X1 U27311 ( .A(n40509), .Z(n40511) );
  BUF_X1 U27312 ( .A(n40569), .Z(n40574) );
  BUF_X1 U27313 ( .A(n40569), .Z(n40573) );
  BUF_X1 U27314 ( .A(n40569), .Z(n40572) );
  BUF_X1 U27315 ( .A(n40569), .Z(n40571) );
  BUF_X1 U27316 ( .A(n40569), .Z(n40570) );
  BUF_X1 U27317 ( .A(n40549), .Z(n40554) );
  BUF_X1 U27318 ( .A(n40549), .Z(n40553) );
  BUF_X1 U27319 ( .A(n40549), .Z(n40552) );
  BUF_X1 U27320 ( .A(n40549), .Z(n40551) );
  BUF_X1 U27321 ( .A(n40549), .Z(n40550) );
  BUF_X1 U27322 ( .A(n40489), .Z(n40494) );
  BUF_X1 U27323 ( .A(n40489), .Z(n40493) );
  BUF_X1 U27324 ( .A(n40489), .Z(n40492) );
  BUF_X1 U27325 ( .A(n40489), .Z(n40491) );
  BUF_X1 U27326 ( .A(n40489), .Z(n40490) );
  BUF_X1 U27327 ( .A(n40469), .Z(n40474) );
  BUF_X1 U27328 ( .A(n40469), .Z(n40473) );
  BUF_X1 U27329 ( .A(n40469), .Z(n40472) );
  BUF_X1 U27330 ( .A(n40469), .Z(n40471) );
  BUF_X1 U27331 ( .A(n40469), .Z(n40470) );
  BUF_X1 U27332 ( .A(n40449), .Z(n40454) );
  BUF_X1 U27333 ( .A(n40449), .Z(n40453) );
  BUF_X1 U27334 ( .A(n40449), .Z(n40452) );
  BUF_X1 U27335 ( .A(n40449), .Z(n40451) );
  BUF_X1 U27336 ( .A(n40449), .Z(n40450) );
  BUF_X1 U27337 ( .A(n40389), .Z(n40394) );
  BUF_X1 U27338 ( .A(n40389), .Z(n40393) );
  BUF_X1 U27339 ( .A(n40389), .Z(n40392) );
  BUF_X1 U27340 ( .A(n40389), .Z(n40391) );
  BUF_X1 U27341 ( .A(n40389), .Z(n40390) );
  BUF_X1 U27342 ( .A(n40369), .Z(n40374) );
  BUF_X1 U27343 ( .A(n40369), .Z(n40373) );
  BUF_X1 U27344 ( .A(n40369), .Z(n40372) );
  BUF_X1 U27345 ( .A(n40369), .Z(n40371) );
  BUF_X1 U27346 ( .A(n40369), .Z(n40370) );
  BUF_X1 U27347 ( .A(n40349), .Z(n40354) );
  BUF_X1 U27348 ( .A(n40349), .Z(n40353) );
  BUF_X1 U27349 ( .A(n40349), .Z(n40352) );
  BUF_X1 U27350 ( .A(n40349), .Z(n40351) );
  BUF_X1 U27351 ( .A(n40349), .Z(n40350) );
  BUF_X1 U27352 ( .A(n40289), .Z(n40294) );
  BUF_X1 U27353 ( .A(n40289), .Z(n40293) );
  BUF_X1 U27354 ( .A(n40289), .Z(n40292) );
  BUF_X1 U27355 ( .A(n40289), .Z(n40291) );
  BUF_X1 U27356 ( .A(n40289), .Z(n40290) );
  BUF_X1 U27357 ( .A(n40269), .Z(n40274) );
  BUF_X1 U27358 ( .A(n40269), .Z(n40273) );
  BUF_X1 U27359 ( .A(n40269), .Z(n40272) );
  BUF_X1 U27360 ( .A(n40269), .Z(n40271) );
  BUF_X1 U27361 ( .A(n40269), .Z(n40270) );
  BUF_X1 U27362 ( .A(n40249), .Z(n40254) );
  BUF_X1 U27363 ( .A(n40249), .Z(n40253) );
  BUF_X1 U27364 ( .A(n40249), .Z(n40252) );
  BUF_X1 U27365 ( .A(n40249), .Z(n40251) );
  BUF_X1 U27366 ( .A(n40249), .Z(n40250) );
  BUF_X1 U27367 ( .A(n40189), .Z(n40194) );
  BUF_X1 U27368 ( .A(n40189), .Z(n40193) );
  BUF_X1 U27369 ( .A(n40189), .Z(n40192) );
  BUF_X1 U27370 ( .A(n40189), .Z(n40191) );
  BUF_X1 U27371 ( .A(n40189), .Z(n40190) );
  BUF_X1 U27372 ( .A(n40169), .Z(n40174) );
  BUF_X1 U27373 ( .A(n40169), .Z(n40173) );
  BUF_X1 U27374 ( .A(n40169), .Z(n40172) );
  BUF_X1 U27375 ( .A(n40169), .Z(n40171) );
  BUF_X1 U27376 ( .A(n40169), .Z(n40170) );
  BUF_X1 U27377 ( .A(n40149), .Z(n40154) );
  BUF_X1 U27378 ( .A(n40149), .Z(n40153) );
  BUF_X1 U27379 ( .A(n40149), .Z(n40152) );
  BUF_X1 U27380 ( .A(n40149), .Z(n40151) );
  BUF_X1 U27381 ( .A(n40149), .Z(n40150) );
  BUF_X1 U27382 ( .A(n40129), .Z(n40134) );
  BUF_X1 U27383 ( .A(n40129), .Z(n40133) );
  BUF_X1 U27384 ( .A(n40129), .Z(n40132) );
  BUF_X1 U27385 ( .A(n40129), .Z(n40131) );
  BUF_X1 U27386 ( .A(n40129), .Z(n40130) );
  BUF_X1 U27387 ( .A(n40109), .Z(n40114) );
  BUF_X1 U27388 ( .A(n40109), .Z(n40113) );
  BUF_X1 U27389 ( .A(n40109), .Z(n40112) );
  BUF_X1 U27390 ( .A(n40109), .Z(n40111) );
  BUF_X1 U27391 ( .A(n40109), .Z(n40110) );
  BUF_X1 U27392 ( .A(n40090), .Z(n40095) );
  BUF_X1 U27393 ( .A(n40090), .Z(n40094) );
  BUF_X1 U27394 ( .A(n40090), .Z(n40093) );
  BUF_X1 U27395 ( .A(n40090), .Z(n40092) );
  BUF_X1 U27396 ( .A(n40090), .Z(n40091) );
  BUF_X1 U27397 ( .A(n40070), .Z(n40075) );
  BUF_X1 U27398 ( .A(n40070), .Z(n40074) );
  BUF_X1 U27399 ( .A(n40070), .Z(n40073) );
  BUF_X1 U27400 ( .A(n40070), .Z(n40072) );
  BUF_X1 U27401 ( .A(n40070), .Z(n40071) );
  BUF_X1 U27402 ( .A(n40050), .Z(n40055) );
  BUF_X1 U27403 ( .A(n40050), .Z(n40054) );
  BUF_X1 U27404 ( .A(n40050), .Z(n40053) );
  BUF_X1 U27405 ( .A(n40050), .Z(n40052) );
  BUF_X1 U27406 ( .A(n40050), .Z(n40051) );
  BUF_X1 U27407 ( .A(n39992), .Z(n39997) );
  BUF_X1 U27408 ( .A(n39992), .Z(n39996) );
  BUF_X1 U27409 ( .A(n39992), .Z(n39995) );
  BUF_X1 U27410 ( .A(n39992), .Z(n39994) );
  BUF_X1 U27411 ( .A(n39992), .Z(n39993) );
  BUF_X1 U27412 ( .A(n39972), .Z(n39977) );
  BUF_X1 U27413 ( .A(n39972), .Z(n39976) );
  BUF_X1 U27414 ( .A(n39972), .Z(n39975) );
  BUF_X1 U27415 ( .A(n39972), .Z(n39974) );
  BUF_X1 U27416 ( .A(n39972), .Z(n39973) );
  BUF_X1 U27417 ( .A(n39874), .Z(n39879) );
  BUF_X1 U27418 ( .A(n39874), .Z(n39878) );
  BUF_X1 U27419 ( .A(n39874), .Z(n39877) );
  BUF_X1 U27420 ( .A(n39874), .Z(n39876) );
  BUF_X1 U27421 ( .A(n39874), .Z(n39875) );
  BUF_X1 U27422 ( .A(n39854), .Z(n39859) );
  BUF_X1 U27423 ( .A(n39854), .Z(n39858) );
  BUF_X1 U27424 ( .A(n39854), .Z(n39857) );
  BUF_X1 U27425 ( .A(n39854), .Z(n39856) );
  BUF_X1 U27426 ( .A(n39854), .Z(n39855) );
  BUF_X1 U27427 ( .A(n39814), .Z(n39819) );
  BUF_X1 U27428 ( .A(n39814), .Z(n39818) );
  BUF_X1 U27429 ( .A(n40402), .Z(n40403) );
  BUF_X1 U27430 ( .A(n39906), .Z(n39907) );
  BUF_X1 U27431 ( .A(n39925), .Z(n39926) );
  BUF_X1 U27432 ( .A(n40202), .Z(n40203) );
  BUF_X1 U27433 ( .A(n40222), .Z(n40223) );
  BUF_X1 U27434 ( .A(n40402), .Z(n40407) );
  BUF_X1 U27435 ( .A(n40402), .Z(n40406) );
  BUF_X1 U27436 ( .A(n40402), .Z(n40405) );
  BUF_X1 U27437 ( .A(n40402), .Z(n40404) );
  BUF_X1 U27438 ( .A(n39906), .Z(n39911) );
  BUF_X1 U27439 ( .A(n39906), .Z(n39910) );
  BUF_X1 U27440 ( .A(n39906), .Z(n39909) );
  BUF_X1 U27441 ( .A(n39906), .Z(n39908) );
  BUF_X1 U27442 ( .A(n39925), .Z(n39930) );
  BUF_X1 U27443 ( .A(n39925), .Z(n39929) );
  BUF_X1 U27444 ( .A(n39925), .Z(n39928) );
  BUF_X1 U27445 ( .A(n39925), .Z(n39927) );
  BUF_X1 U27446 ( .A(n40202), .Z(n40207) );
  BUF_X1 U27447 ( .A(n40202), .Z(n40206) );
  BUF_X1 U27448 ( .A(n40202), .Z(n40205) );
  BUF_X1 U27449 ( .A(n40202), .Z(n40204) );
  BUF_X1 U27450 ( .A(n40222), .Z(n40227) );
  BUF_X1 U27451 ( .A(n40222), .Z(n40226) );
  BUF_X1 U27452 ( .A(n40222), .Z(n40225) );
  BUF_X1 U27453 ( .A(n40222), .Z(n40224) );
  BUF_X1 U27454 ( .A(n40043), .Z(n40046) );
  BUF_X1 U27455 ( .A(n40043), .Z(n40045) );
  BUF_X1 U27456 ( .A(n40043), .Z(n40044) );
  BUF_X1 U27457 ( .A(n39887), .Z(n39892) );
  BUF_X1 U27458 ( .A(n39887), .Z(n39891) );
  BUF_X1 U27459 ( .A(n39887), .Z(n39890) );
  BUF_X1 U27460 ( .A(n39887), .Z(n39889) );
  BUF_X1 U27461 ( .A(n39887), .Z(n39888) );
  BUF_X1 U27462 ( .A(n40422), .Z(n40423) );
  BUF_X1 U27463 ( .A(n40422), .Z(n40427) );
  BUF_X1 U27464 ( .A(n40422), .Z(n40426) );
  BUF_X1 U27465 ( .A(n40422), .Z(n40425) );
  BUF_X1 U27466 ( .A(n40422), .Z(n40424) );
  BUF_X1 U27467 ( .A(n40004), .Z(n40005) );
  BUF_X1 U27468 ( .A(n40023), .Z(n40024) );
  BUF_X1 U27469 ( .A(n40004), .Z(n40009) );
  BUF_X1 U27470 ( .A(n40004), .Z(n40008) );
  BUF_X1 U27471 ( .A(n40004), .Z(n40007) );
  BUF_X1 U27472 ( .A(n40004), .Z(n40006) );
  BUF_X1 U27473 ( .A(n40023), .Z(n40028) );
  BUF_X1 U27474 ( .A(n40023), .Z(n40027) );
  BUF_X1 U27475 ( .A(n40023), .Z(n40026) );
  BUF_X1 U27476 ( .A(n40023), .Z(n40025) );
  BUF_X1 U27477 ( .A(n40302), .Z(n40303) );
  BUF_X1 U27478 ( .A(n40322), .Z(n40323) );
  BUF_X1 U27479 ( .A(n40382), .Z(n40387) );
  BUF_X1 U27480 ( .A(n40382), .Z(n40386) );
  BUF_X1 U27481 ( .A(n40382), .Z(n40385) );
  BUF_X1 U27482 ( .A(n40382), .Z(n40384) );
  BUF_X1 U27483 ( .A(n40382), .Z(n40383) );
  BUF_X1 U27484 ( .A(n40362), .Z(n40367) );
  BUF_X1 U27485 ( .A(n40362), .Z(n40366) );
  BUF_X1 U27486 ( .A(n40362), .Z(n40365) );
  BUF_X1 U27487 ( .A(n40362), .Z(n40364) );
  BUF_X1 U27488 ( .A(n40362), .Z(n40363) );
  BUF_X1 U27489 ( .A(n40242), .Z(n40247) );
  BUF_X1 U27490 ( .A(n40242), .Z(n40246) );
  BUF_X1 U27491 ( .A(n40242), .Z(n40245) );
  BUF_X1 U27492 ( .A(n40242), .Z(n40244) );
  BUF_X1 U27493 ( .A(n40242), .Z(n40243) );
  BUF_X1 U27494 ( .A(n40083), .Z(n40088) );
  BUF_X1 U27495 ( .A(n40083), .Z(n40087) );
  BUF_X1 U27496 ( .A(n40083), .Z(n40086) );
  BUF_X1 U27497 ( .A(n40083), .Z(n40085) );
  BUF_X1 U27498 ( .A(n40083), .Z(n40084) );
  BUF_X1 U27499 ( .A(n40063), .Z(n40068) );
  BUF_X1 U27500 ( .A(n40063), .Z(n40067) );
  BUF_X1 U27501 ( .A(n40063), .Z(n40066) );
  BUF_X1 U27502 ( .A(n40063), .Z(n40065) );
  BUF_X1 U27503 ( .A(n40063), .Z(n40064) );
  BUF_X1 U27504 ( .A(n40043), .Z(n40048) );
  BUF_X1 U27505 ( .A(n40043), .Z(n40047) );
  BUF_X1 U27506 ( .A(n39827), .Z(n39828) );
  BUF_X1 U27507 ( .A(n40302), .Z(n40307) );
  BUF_X1 U27508 ( .A(n40302), .Z(n40306) );
  BUF_X1 U27509 ( .A(n40302), .Z(n40305) );
  BUF_X1 U27510 ( .A(n40302), .Z(n40304) );
  BUF_X1 U27511 ( .A(n40322), .Z(n40327) );
  BUF_X1 U27512 ( .A(n40322), .Z(n40326) );
  BUF_X1 U27513 ( .A(n40322), .Z(n40325) );
  BUF_X1 U27514 ( .A(n40322), .Z(n40324) );
  BUF_X1 U27515 ( .A(n39827), .Z(n39832) );
  BUF_X1 U27516 ( .A(n39827), .Z(n39831) );
  BUF_X1 U27517 ( .A(n39827), .Z(n39830) );
  BUF_X1 U27518 ( .A(n39827), .Z(n39829) );
  BUF_X1 U27519 ( .A(n39807), .Z(n39810) );
  BUF_X1 U27520 ( .A(n39807), .Z(n39809) );
  BUF_X1 U27521 ( .A(n39807), .Z(n39808) );
  BUF_X1 U27522 ( .A(n40342), .Z(n40347) );
  BUF_X1 U27523 ( .A(n40342), .Z(n40346) );
  BUF_X1 U27524 ( .A(n40342), .Z(n40345) );
  BUF_X1 U27525 ( .A(n40342), .Z(n40344) );
  BUF_X1 U27526 ( .A(n40342), .Z(n40343) );
  BUF_X1 U27527 ( .A(n40282), .Z(n40287) );
  BUF_X1 U27528 ( .A(n40282), .Z(n40286) );
  BUF_X1 U27529 ( .A(n40282), .Z(n40285) );
  BUF_X1 U27530 ( .A(n40282), .Z(n40284) );
  BUF_X1 U27531 ( .A(n40282), .Z(n40283) );
  BUF_X1 U27532 ( .A(n40262), .Z(n40267) );
  BUF_X1 U27533 ( .A(n40262), .Z(n40266) );
  BUF_X1 U27534 ( .A(n40262), .Z(n40265) );
  BUF_X1 U27535 ( .A(n40262), .Z(n40264) );
  BUF_X1 U27536 ( .A(n40262), .Z(n40263) );
  BUF_X1 U27537 ( .A(n40182), .Z(n40187) );
  BUF_X1 U27538 ( .A(n40182), .Z(n40186) );
  BUF_X1 U27539 ( .A(n40182), .Z(n40185) );
  BUF_X1 U27540 ( .A(n40182), .Z(n40184) );
  BUF_X1 U27541 ( .A(n40182), .Z(n40183) );
  BUF_X1 U27542 ( .A(n40162), .Z(n40167) );
  BUF_X1 U27543 ( .A(n40162), .Z(n40166) );
  BUF_X1 U27544 ( .A(n40162), .Z(n40165) );
  BUF_X1 U27545 ( .A(n40162), .Z(n40164) );
  BUF_X1 U27546 ( .A(n40162), .Z(n40163) );
  BUF_X1 U27547 ( .A(n40142), .Z(n40147) );
  BUF_X1 U27548 ( .A(n40142), .Z(n40146) );
  BUF_X1 U27549 ( .A(n40142), .Z(n40145) );
  BUF_X1 U27550 ( .A(n40142), .Z(n40144) );
  BUF_X1 U27551 ( .A(n40142), .Z(n40143) );
  BUF_X1 U27552 ( .A(n40122), .Z(n40127) );
  BUF_X1 U27553 ( .A(n40122), .Z(n40126) );
  BUF_X1 U27554 ( .A(n40122), .Z(n40125) );
  BUF_X1 U27555 ( .A(n40122), .Z(n40124) );
  BUF_X1 U27556 ( .A(n40122), .Z(n40123) );
  BUF_X1 U27557 ( .A(n40102), .Z(n40107) );
  BUF_X1 U27558 ( .A(n40102), .Z(n40106) );
  BUF_X1 U27559 ( .A(n40102), .Z(n40105) );
  BUF_X1 U27560 ( .A(n40102), .Z(n40104) );
  BUF_X1 U27561 ( .A(n40102), .Z(n40103) );
  BUF_X1 U27562 ( .A(n39985), .Z(n39990) );
  BUF_X1 U27563 ( .A(n39985), .Z(n39989) );
  BUF_X1 U27564 ( .A(n39985), .Z(n39988) );
  BUF_X1 U27565 ( .A(n39985), .Z(n39987) );
  BUF_X1 U27566 ( .A(n39985), .Z(n39986) );
  BUF_X1 U27567 ( .A(n39965), .Z(n39970) );
  BUF_X1 U27568 ( .A(n39965), .Z(n39969) );
  BUF_X1 U27569 ( .A(n39965), .Z(n39968) );
  BUF_X1 U27570 ( .A(n39965), .Z(n39967) );
  BUF_X1 U27571 ( .A(n39965), .Z(n39966) );
  BUF_X1 U27572 ( .A(n39945), .Z(n39950) );
  BUF_X1 U27573 ( .A(n39945), .Z(n39949) );
  BUF_X1 U27574 ( .A(n39945), .Z(n39948) );
  BUF_X1 U27575 ( .A(n39945), .Z(n39947) );
  BUF_X1 U27576 ( .A(n39945), .Z(n39946) );
  BUF_X1 U27577 ( .A(n39867), .Z(n39872) );
  BUF_X1 U27578 ( .A(n39867), .Z(n39871) );
  BUF_X1 U27579 ( .A(n39867), .Z(n39870) );
  BUF_X1 U27580 ( .A(n39867), .Z(n39869) );
  BUF_X1 U27581 ( .A(n39867), .Z(n39868) );
  BUF_X1 U27582 ( .A(n39847), .Z(n39852) );
  BUF_X1 U27583 ( .A(n39847), .Z(n39851) );
  BUF_X1 U27584 ( .A(n39847), .Z(n39850) );
  BUF_X1 U27585 ( .A(n39847), .Z(n39849) );
  BUF_X1 U27586 ( .A(n39847), .Z(n39848) );
  BUF_X1 U27587 ( .A(n39807), .Z(n39812) );
  BUF_X1 U27588 ( .A(n39807), .Z(n39811) );
  BUF_X1 U27589 ( .A(n33391), .Z(n39952) );
  BUF_X1 U27590 ( .A(n33406), .Z(n39894) );
  BUF_X1 U27591 ( .A(n33403), .Z(n39913) );
  BUF_X1 U27592 ( .A(n33399), .Z(n39932) );
  AND2_X1 U27593 ( .A1(n37228), .A2(n37246), .ZN(n36016) );
  BUF_X1 U27594 ( .A(n35981), .Z(n39289) );
  BUF_X1 U27595 ( .A(n35981), .Z(n39290) );
  BUF_X1 U27596 ( .A(n35981), .Z(n39291) );
  BUF_X1 U27597 ( .A(n35981), .Z(n39288) );
  BUF_X1 U27598 ( .A(n35981), .Z(n39292) );
  BUF_X1 U27599 ( .A(n33426), .Z(n39794) );
  BUF_X1 U27600 ( .A(n34700), .Z(n39542) );
  BUF_X1 U27601 ( .A(n33426), .Z(n39793) );
  BUF_X1 U27602 ( .A(n34700), .Z(n39541) );
  BUF_X1 U27603 ( .A(n33426), .Z(n39792) );
  BUF_X1 U27604 ( .A(n34700), .Z(n39540) );
  BUF_X1 U27605 ( .A(n33426), .Z(n39791) );
  BUF_X1 U27606 ( .A(n34700), .Z(n39539) );
  BUF_X1 U27607 ( .A(n33426), .Z(n39790) );
  BUF_X1 U27608 ( .A(n34700), .Z(n39538) );
  OAI221_X1 U27609 ( .B1(n33264), .B2(n33307), .C1(n33265), .C2(n33308), .A(
        n41366), .ZN(n33311) );
  OAI221_X1 U27610 ( .B1(n33274), .B2(n33339), .C1(n33275), .C2(n33340), .A(
        n41366), .ZN(n33349) );
  OAI221_X1 U27611 ( .B1(n33274), .B2(n33307), .C1(n33275), .C2(n33308), .A(
        n41366), .ZN(n33317) );
  OAI221_X1 U27612 ( .B1(n33264), .B2(n33339), .C1(n33265), .C2(n33340), .A(
        n41366), .ZN(n33343) );
  OAI221_X1 U27613 ( .B1(n33264), .B2(n33368), .C1(n33265), .C2(n33369), .A(
        n41366), .ZN(n33372) );
  OAI221_X1 U27614 ( .B1(n33274), .B2(n33368), .C1(n33275), .C2(n33369), .A(
        n41365), .ZN(n33378) );
  OAI221_X1 U27615 ( .B1(n33269), .B2(n33339), .C1(n33270), .C2(n33340), .A(
        n41366), .ZN(n33346) );
  OAI221_X1 U27616 ( .B1(n33269), .B2(n33307), .C1(n33270), .C2(n33308), .A(
        n41366), .ZN(n33314) );
  OAI221_X1 U27617 ( .B1(n33269), .B2(n33368), .C1(n33270), .C2(n33369), .A(
        n41364), .ZN(n33375) );
  OAI221_X1 U27618 ( .B1(n33270), .B2(n33396), .C1(n33269), .C2(n33397), .A(
        n41365), .ZN(n33405) );
  OAI221_X1 U27619 ( .B1(n33265), .B2(n33396), .C1(n33264), .C2(n33397), .A(
        n41365), .ZN(n33401) );
  OAI221_X1 U27620 ( .B1(n33290), .B2(n33396), .C1(n32159), .C2(n33397), .A(
        n41364), .ZN(n33417) );
  OAI221_X1 U27621 ( .B1(n33260), .B2(n33396), .C1(n33255), .C2(n33397), .A(
        n41365), .ZN(n33393) );
  OAI221_X1 U27622 ( .B1(n33275), .B2(n33396), .C1(n33274), .C2(n33397), .A(
        n41364), .ZN(n33408) );
  OAI221_X1 U27623 ( .B1(n33280), .B2(n33396), .C1(n32157), .C2(n33397), .A(
        n41364), .ZN(n33411) );
  OAI221_X1 U27624 ( .B1(n33285), .B2(n33396), .C1(n32158), .C2(n33397), .A(
        n41364), .ZN(n33414) );
  OAI221_X1 U27625 ( .B1(n33255), .B2(n33307), .C1(n33260), .C2(n33308), .A(
        n41365), .ZN(n33304) );
  OAI221_X1 U27626 ( .B1(n32158), .B2(n33368), .C1(n33285), .C2(n33369), .A(
        n41365), .ZN(n33384) );
  OAI221_X1 U27627 ( .B1(n32157), .B2(n33368), .C1(n33280), .C2(n33369), .A(
        n41365), .ZN(n33381) );
  OAI221_X1 U27628 ( .B1(n32159), .B2(n33307), .C1(n33290), .C2(n33308), .A(
        n41367), .ZN(n33326) );
  OAI221_X1 U27629 ( .B1(n32158), .B2(n33307), .C1(n33285), .C2(n33308), .A(
        n41366), .ZN(n33323) );
  OAI221_X1 U27630 ( .B1(n32157), .B2(n33307), .C1(n33280), .C2(n33308), .A(
        n41367), .ZN(n33320) );
  OAI221_X1 U27631 ( .B1(n32160), .B2(n33307), .C1(n33296), .C2(n33308), .A(
        n41365), .ZN(n33329) );
  OAI221_X1 U27632 ( .B1(n33255), .B2(n33339), .C1(n33260), .C2(n33340), .A(
        n41367), .ZN(n33336) );
  OAI221_X1 U27633 ( .B1(n32157), .B2(n33339), .C1(n33280), .C2(n33340), .A(
        n41366), .ZN(n33352) );
  OAI221_X1 U27634 ( .B1(n32158), .B2(n33339), .C1(n33285), .C2(n33340), .A(
        n41366), .ZN(n33355) );
  OAI221_X1 U27635 ( .B1(n32159), .B2(n33339), .C1(n33290), .C2(n33340), .A(
        n41366), .ZN(n33358) );
  OAI221_X1 U27636 ( .B1(n32160), .B2(n33339), .C1(n33296), .C2(n33340), .A(
        n41366), .ZN(n33361) );
  OAI221_X1 U27637 ( .B1(n33255), .B2(n33368), .C1(n33260), .C2(n33369), .A(
        n41366), .ZN(n33365) );
  OAI221_X1 U27638 ( .B1(n32159), .B2(n33368), .C1(n33290), .C2(n33369), .A(
        n41365), .ZN(n33387) );
  OAI221_X1 U27639 ( .B1(n32160), .B2(n33368), .C1(n33296), .C2(n33369), .A(
        n41365), .ZN(n33390) );
  OAI221_X1 U27640 ( .B1(n32160), .B2(n33397), .C1(n33296), .C2(n33396), .A(
        n41364), .ZN(n33420) );
  NOR3_X1 U27641 ( .A1(n32251), .A2(n32254), .A3(n32248), .ZN(n37228) );
  NOR2_X1 U27642 ( .A1(n32246), .A2(n32243), .ZN(n37246) );
  NOR3_X1 U27643 ( .A1(n32168), .A2(n32166), .A3(n32165), .ZN(n34674) );
  NOR3_X1 U27644 ( .A1(n32173), .A2(n32171), .A3(n32170), .ZN(n35948) );
  INV_X1 U27645 ( .A(n33295), .ZN(n32160) );
  INV_X1 U27646 ( .A(n33289), .ZN(n32159) );
  INV_X1 U27647 ( .A(n33279), .ZN(n32157) );
  INV_X1 U27648 ( .A(n33284), .ZN(n32158) );
  NAND2_X1 U27649 ( .A1(n33333), .A2(n33294), .ZN(n33397) );
  INV_X1 U27650 ( .A(n33264), .ZN(n32154) );
  INV_X1 U27651 ( .A(n33274), .ZN(n32156) );
  INV_X1 U27652 ( .A(n33269), .ZN(n32155) );
  NAND2_X1 U27653 ( .A1(n37249), .A2(n37228), .ZN(n36033) );
  NAND2_X1 U27654 ( .A1(n37249), .A2(n37234), .ZN(n36039) );
  NAND2_X1 U27655 ( .A1(n37249), .A2(n37230), .ZN(n36038) );
  NAND2_X1 U27656 ( .A1(n37249), .A2(n37231), .ZN(n36037) );
  NAND2_X1 U27657 ( .A1(n34693), .A2(n34673), .ZN(n33478) );
  NAND2_X1 U27658 ( .A1(n34693), .A2(n34679), .ZN(n33484) );
  NAND2_X1 U27659 ( .A1(n34693), .A2(n34675), .ZN(n33483) );
  NAND2_X1 U27660 ( .A1(n34693), .A2(n34676), .ZN(n33482) );
  NAND2_X1 U27661 ( .A1(n35967), .A2(n35947), .ZN(n34752) );
  NAND2_X1 U27662 ( .A1(n35967), .A2(n35953), .ZN(n34758) );
  NAND2_X1 U27663 ( .A1(n35967), .A2(n35949), .ZN(n34757) );
  NAND2_X1 U27664 ( .A1(n35967), .A2(n35950), .ZN(n34756) );
  BUF_X1 U27665 ( .A(n33273), .Z(n40517) );
  BUF_X1 U27666 ( .A(n33273), .Z(n40518) );
  BUF_X1 U27667 ( .A(n33273), .Z(n40519) );
  BUF_X1 U27668 ( .A(n33273), .Z(n40520) );
  BUF_X1 U27669 ( .A(n33273), .Z(n40516) );
  BUF_X1 U27670 ( .A(n33263), .Z(n40556) );
  BUF_X1 U27671 ( .A(n33263), .Z(n40557) );
  BUF_X1 U27672 ( .A(n33263), .Z(n40558) );
  BUF_X1 U27673 ( .A(n33263), .Z(n40559) );
  BUF_X1 U27674 ( .A(n33263), .Z(n40560) );
  BUF_X1 U27675 ( .A(n33268), .Z(n40536) );
  BUF_X1 U27676 ( .A(n33268), .Z(n40537) );
  BUF_X1 U27677 ( .A(n33268), .Z(n40538) );
  BUF_X1 U27678 ( .A(n33268), .Z(n40539) );
  BUF_X1 U27679 ( .A(n33268), .Z(n40540) );
  BUF_X1 U27680 ( .A(n33278), .Z(n40497) );
  BUF_X1 U27681 ( .A(n33278), .Z(n40498) );
  BUF_X1 U27682 ( .A(n33278), .Z(n40499) );
  BUF_X1 U27683 ( .A(n33278), .Z(n40500) );
  BUF_X1 U27684 ( .A(n33278), .Z(n40496) );
  BUF_X1 U27685 ( .A(n33254), .Z(n40579) );
  BUF_X1 U27686 ( .A(n33254), .Z(n40580) );
  BUF_X1 U27687 ( .A(n33254), .Z(n40576) );
  BUF_X1 U27688 ( .A(n33254), .Z(n40578) );
  BUF_X1 U27689 ( .A(n33254), .Z(n40577) );
  BUF_X1 U27690 ( .A(n33283), .Z(n40476) );
  BUF_X1 U27691 ( .A(n33283), .Z(n40477) );
  BUF_X1 U27692 ( .A(n33283), .Z(n40478) );
  BUF_X1 U27693 ( .A(n33283), .Z(n40479) );
  BUF_X1 U27694 ( .A(n33283), .Z(n40480) );
  BUF_X1 U27695 ( .A(n33288), .Z(n40456) );
  BUF_X1 U27696 ( .A(n33288), .Z(n40457) );
  BUF_X1 U27697 ( .A(n33288), .Z(n40458) );
  BUF_X1 U27698 ( .A(n33288), .Z(n40459) );
  BUF_X1 U27699 ( .A(n33288), .Z(n40460) );
  BUF_X1 U27700 ( .A(n33293), .Z(n40436) );
  BUF_X1 U27701 ( .A(n33293), .Z(n40437) );
  BUF_X1 U27702 ( .A(n33293), .Z(n40438) );
  BUF_X1 U27703 ( .A(n33293), .Z(n40439) );
  BUF_X1 U27704 ( .A(n33293), .Z(n40440) );
  BUF_X1 U27705 ( .A(n40582), .Z(n40585) );
  BUF_X1 U27706 ( .A(n40582), .Z(n40584) );
  BUF_X1 U27707 ( .A(n40582), .Z(n40587) );
  BUF_X1 U27708 ( .A(n40582), .Z(n40586) );
  BUF_X1 U27709 ( .A(n40582), .Z(n40583) );
  NAND2_X1 U27710 ( .A1(n37226), .A2(n37227), .ZN(n35993) );
  NAND2_X1 U27711 ( .A1(n37226), .A2(n37228), .ZN(n35992) );
  NAND2_X1 U27712 ( .A1(n37226), .A2(n37229), .ZN(n35991) );
  NAND2_X1 U27713 ( .A1(n37226), .A2(n37233), .ZN(n35999) );
  NAND2_X1 U27714 ( .A1(n37226), .A2(n37234), .ZN(n35998) );
  NAND2_X1 U27715 ( .A1(n37226), .A2(n37235), .ZN(n35997) );
  BUF_X1 U27716 ( .A(n40522), .Z(n40523) );
  BUF_X1 U27717 ( .A(n40522), .Z(n40527) );
  BUF_X1 U27718 ( .A(n40522), .Z(n40526) );
  BUF_X1 U27719 ( .A(n40522), .Z(n40525) );
  BUF_X1 U27720 ( .A(n40522), .Z(n40524) );
  BUF_X1 U27721 ( .A(n40502), .Z(n40503) );
  BUF_X1 U27722 ( .A(n40502), .Z(n40507) );
  BUF_X1 U27723 ( .A(n40502), .Z(n40506) );
  BUF_X1 U27724 ( .A(n40502), .Z(n40505) );
  BUF_X1 U27725 ( .A(n40502), .Z(n40504) );
  BUF_X1 U27726 ( .A(n40562), .Z(n40567) );
  BUF_X1 U27727 ( .A(n40562), .Z(n40566) );
  BUF_X1 U27728 ( .A(n40562), .Z(n40565) );
  BUF_X1 U27729 ( .A(n40562), .Z(n40564) );
  BUF_X1 U27730 ( .A(n40562), .Z(n40563) );
  BUF_X1 U27731 ( .A(n40542), .Z(n40547) );
  BUF_X1 U27732 ( .A(n40542), .Z(n40546) );
  BUF_X1 U27733 ( .A(n40542), .Z(n40545) );
  BUF_X1 U27734 ( .A(n40542), .Z(n40544) );
  BUF_X1 U27735 ( .A(n40542), .Z(n40543) );
  BUF_X1 U27736 ( .A(n40482), .Z(n40487) );
  BUF_X1 U27737 ( .A(n40482), .Z(n40486) );
  BUF_X1 U27738 ( .A(n40482), .Z(n40485) );
  BUF_X1 U27739 ( .A(n40482), .Z(n40484) );
  BUF_X1 U27740 ( .A(n40482), .Z(n40483) );
  BUF_X1 U27741 ( .A(n40462), .Z(n40467) );
  BUF_X1 U27742 ( .A(n40462), .Z(n40466) );
  BUF_X1 U27743 ( .A(n40462), .Z(n40465) );
  BUF_X1 U27744 ( .A(n40462), .Z(n40464) );
  BUF_X1 U27745 ( .A(n40462), .Z(n40463) );
  BUF_X1 U27746 ( .A(n40442), .Z(n40447) );
  BUF_X1 U27747 ( .A(n40442), .Z(n40446) );
  BUF_X1 U27748 ( .A(n40442), .Z(n40445) );
  BUF_X1 U27749 ( .A(n40442), .Z(n40444) );
  BUF_X1 U27750 ( .A(n40442), .Z(n40443) );
  NAND2_X1 U27751 ( .A1(n37235), .A2(n37239), .ZN(n36021) );
  NAND2_X1 U27752 ( .A1(n37234), .A2(n37239), .ZN(n36019) );
  NAND2_X1 U27753 ( .A1(n37228), .A2(n37239), .ZN(n36009) );
  NAND2_X1 U27754 ( .A1(n37233), .A2(n37246), .ZN(n36031) );
  NAND2_X1 U27755 ( .A1(n37230), .A2(n37246), .ZN(n36027) );
  NAND2_X1 U27756 ( .A1(n37227), .A2(n37246), .ZN(n36025) );
  NAND2_X1 U27757 ( .A1(n34675), .A2(n34690), .ZN(n33472) );
  NAND2_X1 U27758 ( .A1(n35949), .A2(n35964), .ZN(n34746) );
  NAND2_X1 U27759 ( .A1(n37229), .A2(n37246), .ZN(n36026) );
  NAND2_X1 U27760 ( .A1(n37229), .A2(n37239), .ZN(n36011) );
  NAND2_X1 U27761 ( .A1(n34680), .A2(n34684), .ZN(n33466) );
  NAND2_X1 U27762 ( .A1(n34679), .A2(n34684), .ZN(n33464) );
  NAND2_X1 U27763 ( .A1(n34679), .A2(n34672), .ZN(n33443) );
  NAND2_X1 U27764 ( .A1(n34680), .A2(n34672), .ZN(n33442) );
  NAND2_X1 U27765 ( .A1(n35954), .A2(n35958), .ZN(n34740) );
  NAND2_X1 U27766 ( .A1(n35953), .A2(n35958), .ZN(n34738) );
  NAND2_X1 U27767 ( .A1(n35953), .A2(n35946), .ZN(n34717) );
  NAND2_X1 U27768 ( .A1(n35954), .A2(n35946), .ZN(n34716) );
  NAND2_X1 U27769 ( .A1(n34678), .A2(n34690), .ZN(n33476) );
  NAND2_X1 U27770 ( .A1(n34671), .A2(n34690), .ZN(n33470) );
  NAND2_X1 U27771 ( .A1(n34671), .A2(n34672), .ZN(n33438) );
  NAND2_X1 U27772 ( .A1(n34673), .A2(n34672), .ZN(n33437) );
  NAND2_X1 U27773 ( .A1(n34678), .A2(n34672), .ZN(n33444) );
  NAND2_X1 U27774 ( .A1(n34673), .A2(n34684), .ZN(n33454) );
  NAND2_X1 U27775 ( .A1(n35952), .A2(n35964), .ZN(n34750) );
  NAND2_X1 U27776 ( .A1(n35945), .A2(n35964), .ZN(n34744) );
  NAND2_X1 U27777 ( .A1(n35945), .A2(n35946), .ZN(n34712) );
  NAND2_X1 U27778 ( .A1(n35947), .A2(n35946), .ZN(n34711) );
  NAND2_X1 U27779 ( .A1(n35952), .A2(n35946), .ZN(n34718) );
  NAND2_X1 U27780 ( .A1(n35947), .A2(n35958), .ZN(n34728) );
  NAND2_X1 U27781 ( .A1(n37239), .A2(n37231), .ZN(n36020) );
  NAND2_X1 U27782 ( .A1(n34690), .A2(n34680), .ZN(n33477) );
  NAND2_X1 U27783 ( .A1(n35964), .A2(n35954), .ZN(n34751) );
  NAND2_X1 U27784 ( .A1(n37246), .A2(n37235), .ZN(n36032) );
  NAND2_X1 U27785 ( .A1(n34674), .A2(n34690), .ZN(n33471) );
  NAND2_X1 U27786 ( .A1(n34674), .A2(n34672), .ZN(n33436) );
  NAND2_X1 U27787 ( .A1(n34674), .A2(n34684), .ZN(n33456) );
  NAND2_X1 U27788 ( .A1(n35948), .A2(n35964), .ZN(n34745) );
  NAND2_X1 U27789 ( .A1(n35948), .A2(n35946), .ZN(n34710) );
  NAND2_X1 U27790 ( .A1(n35948), .A2(n35958), .ZN(n34730) );
  AND2_X1 U27791 ( .A1(n33331), .A2(n33294), .ZN(n33395) );
  INV_X1 U27792 ( .A(n33255), .ZN(n32153) );
  NAND2_X1 U27793 ( .A1(n37236), .A2(n37233), .ZN(n36010) );
  NAND2_X1 U27794 ( .A1(n37236), .A2(n37231), .ZN(n36005) );
  NAND2_X1 U27795 ( .A1(n37236), .A2(n37227), .ZN(n36004) );
  NAND2_X1 U27796 ( .A1(n37236), .A2(n37230), .ZN(n36003) );
  NAND2_X1 U27797 ( .A1(n34684), .A2(n34676), .ZN(n33465) );
  NAND2_X1 U27798 ( .A1(n34681), .A2(n34676), .ZN(n33450) );
  NAND2_X1 U27799 ( .A1(n35958), .A2(n35950), .ZN(n34739) );
  NAND2_X1 U27800 ( .A1(n35955), .A2(n35950), .ZN(n34724) );
  NAND2_X1 U27801 ( .A1(n34681), .A2(n34671), .ZN(n33449) );
  NAND2_X1 U27802 ( .A1(n35955), .A2(n35945), .ZN(n34723) );
  NAND2_X1 U27803 ( .A1(n34681), .A2(n34675), .ZN(n33448) );
  NAND2_X1 U27804 ( .A1(n35955), .A2(n35949), .ZN(n34722) );
  NAND2_X1 U27805 ( .A1(n34681), .A2(n34678), .ZN(n33455) );
  NAND2_X1 U27806 ( .A1(n35955), .A2(n35952), .ZN(n34729) );
  BUF_X1 U27807 ( .A(n33310), .Z(n40402) );
  OAI211_X1 U27808 ( .C1(n33264), .C2(n33305), .A(n40401), .B(n41367), .ZN(
        n33310) );
  BUF_X1 U27809 ( .A(n33400), .Z(n39925) );
  OAI211_X1 U27810 ( .C1(n33264), .C2(n33394), .A(n39920), .B(n41369), .ZN(
        n33400) );
  BUF_X1 U27811 ( .A(n33348), .Z(n40202) );
  OAI211_X1 U27812 ( .C1(n33274), .C2(n33337), .A(n40201), .B(n41368), .ZN(
        n33348) );
  BUF_X1 U27813 ( .A(n33316), .Z(n40362) );
  OAI211_X1 U27814 ( .C1(n33274), .C2(n33305), .A(n40361), .B(n41368), .ZN(
        n33316) );
  BUF_X1 U27815 ( .A(n33342), .Z(n40242) );
  OAI211_X1 U27816 ( .C1(n33264), .C2(n33337), .A(n40241), .B(n41368), .ZN(
        n33342) );
  BUF_X1 U27817 ( .A(n33371), .Z(n40083) );
  OAI211_X1 U27818 ( .C1(n33264), .C2(n33366), .A(n40082), .B(n41369), .ZN(
        n33371) );
  BUF_X1 U27819 ( .A(n33377), .Z(n40043) );
  OAI211_X1 U27820 ( .C1(n33274), .C2(n33366), .A(n40042), .B(n41369), .ZN(
        n33377) );
  BUF_X1 U27821 ( .A(n33407), .Z(n39887) );
  OAI211_X1 U27822 ( .C1(n33274), .C2(n33394), .A(n39886), .B(n41369), .ZN(
        n33407) );
  BUF_X1 U27823 ( .A(n33404), .Z(n39906) );
  OAI211_X1 U27824 ( .C1(n33269), .C2(n33394), .A(n39901), .B(n41369), .ZN(
        n33404) );
  BUF_X1 U27825 ( .A(n33345), .Z(n40222) );
  OAI211_X1 U27826 ( .C1(n33269), .C2(n33337), .A(n40221), .B(n41368), .ZN(
        n33345) );
  BUF_X1 U27827 ( .A(n33313), .Z(n40382) );
  OAI211_X1 U27828 ( .C1(n33269), .C2(n33305), .A(n40381), .B(n41367), .ZN(
        n33313) );
  BUF_X1 U27829 ( .A(n33374), .Z(n40063) );
  OAI211_X1 U27830 ( .C1(n33269), .C2(n33366), .A(n40062), .B(n41369), .ZN(
        n33374) );
  BUF_X1 U27831 ( .A(n33303), .Z(n40422) );
  OAI211_X1 U27832 ( .C1(n33255), .C2(n33305), .A(n40421), .B(n41368), .ZN(
        n33303) );
  BUF_X1 U27833 ( .A(n33383), .Z(n40004) );
  OAI211_X1 U27834 ( .C1(n32158), .C2(n33366), .A(n39999), .B(n41369), .ZN(
        n33383) );
  BUF_X1 U27835 ( .A(n33380), .Z(n40023) );
  OAI211_X1 U27836 ( .C1(n32157), .C2(n33366), .A(n40018), .B(n41369), .ZN(
        n33380) );
  BUF_X1 U27837 ( .A(n33325), .Z(n40302) );
  OAI211_X1 U27838 ( .C1(n32159), .C2(n33305), .A(n40301), .B(n41368), .ZN(
        n33325) );
  BUF_X1 U27839 ( .A(n33322), .Z(n40322) );
  OAI211_X1 U27840 ( .C1(n32158), .C2(n33305), .A(n40321), .B(n41367), .ZN(
        n33322) );
  BUF_X1 U27841 ( .A(n33319), .Z(n40342) );
  OAI211_X1 U27842 ( .C1(n32157), .C2(n33305), .A(n40341), .B(n41368), .ZN(
        n33319) );
  BUF_X1 U27843 ( .A(n33328), .Z(n40282) );
  OAI211_X1 U27844 ( .C1(n32160), .C2(n33305), .A(n40281), .B(n41368), .ZN(
        n33328) );
  BUF_X1 U27845 ( .A(n33335), .Z(n40262) );
  OAI211_X1 U27846 ( .C1(n33255), .C2(n33337), .A(n40261), .B(n41368), .ZN(
        n33335) );
  BUF_X1 U27847 ( .A(n33351), .Z(n40182) );
  OAI211_X1 U27848 ( .C1(n32157), .C2(n33337), .A(n40181), .B(n41368), .ZN(
        n33351) );
  BUF_X1 U27849 ( .A(n33354), .Z(n40162) );
  OAI211_X1 U27850 ( .C1(n32158), .C2(n33337), .A(n40161), .B(n41368), .ZN(
        n33354) );
  BUF_X1 U27851 ( .A(n33357), .Z(n40142) );
  OAI211_X1 U27852 ( .C1(n32159), .C2(n33337), .A(n40141), .B(n41369), .ZN(
        n33357) );
  BUF_X1 U27853 ( .A(n33360), .Z(n40122) );
  OAI211_X1 U27854 ( .C1(n32160), .C2(n33337), .A(n40116), .B(n41369), .ZN(
        n33360) );
  BUF_X1 U27855 ( .A(n33364), .Z(n40102) );
  OAI211_X1 U27856 ( .C1(n33255), .C2(n33366), .A(n40097), .B(n41369), .ZN(
        n33364) );
  BUF_X1 U27857 ( .A(n33386), .Z(n39985) );
  OAI211_X1 U27858 ( .C1(n32159), .C2(n33366), .A(n39984), .B(n41369), .ZN(
        n33386) );
  BUF_X1 U27859 ( .A(n33389), .Z(n39965) );
  OAI211_X1 U27860 ( .C1(n32160), .C2(n33366), .A(n39964), .B(n41369), .ZN(
        n33389) );
  BUF_X1 U27861 ( .A(n33392), .Z(n39945) );
  OAI211_X1 U27862 ( .C1(n33255), .C2(n33394), .A(n39944), .B(n41369), .ZN(
        n33392) );
  BUF_X1 U27863 ( .A(n33416), .Z(n39827) );
  OAI211_X1 U27864 ( .C1(n32159), .C2(n33394), .A(n39826), .B(n41370), .ZN(
        n33416) );
  BUF_X1 U27865 ( .A(n33410), .Z(n39867) );
  OAI211_X1 U27866 ( .C1(n32157), .C2(n33394), .A(n39866), .B(n41370), .ZN(
        n33410) );
  BUF_X1 U27867 ( .A(n33413), .Z(n39847) );
  OAI211_X1 U27868 ( .C1(n32158), .C2(n33394), .A(n39846), .B(n41370), .ZN(
        n33413) );
  BUF_X1 U27869 ( .A(n33419), .Z(n39807) );
  OAI211_X1 U27870 ( .C1(n32160), .C2(n33394), .A(n39802), .B(n41370), .ZN(
        n33419) );
  BUF_X1 U27871 ( .A(n33302), .Z(n40429) );
  BUF_X1 U27872 ( .A(n33309), .Z(n40409) );
  BUF_X1 U27873 ( .A(n33347), .Z(n40209) );
  BUF_X1 U27874 ( .A(n33344), .Z(n40229) );
  BUF_X1 U27875 ( .A(n33324), .Z(n40309) );
  BUF_X1 U27876 ( .A(n33321), .Z(n40329) );
  BUF_X1 U27877 ( .A(n33415), .Z(n39834) );
  BUF_X1 U27878 ( .A(n33271), .Z(n40529) );
  BUF_X1 U27879 ( .A(n33276), .Z(n40509) );
  BUF_X1 U27880 ( .A(n33252), .Z(n40589) );
  BUF_X1 U27881 ( .A(n33261), .Z(n40569) );
  BUF_X1 U27882 ( .A(n33266), .Z(n40549) );
  BUF_X1 U27883 ( .A(n33281), .Z(n40489) );
  BUF_X1 U27884 ( .A(n33286), .Z(n40469) );
  BUF_X1 U27885 ( .A(n33291), .Z(n40449) );
  BUF_X1 U27886 ( .A(n33312), .Z(n40389) );
  BUF_X1 U27887 ( .A(n33315), .Z(n40369) );
  BUF_X1 U27888 ( .A(n33318), .Z(n40349) );
  BUF_X1 U27889 ( .A(n33327), .Z(n40289) );
  BUF_X1 U27890 ( .A(n33334), .Z(n40269) );
  BUF_X1 U27891 ( .A(n33341), .Z(n40249) );
  BUF_X1 U27892 ( .A(n33350), .Z(n40189) );
  BUF_X1 U27893 ( .A(n33353), .Z(n40169) );
  BUF_X1 U27894 ( .A(n33356), .Z(n40149) );
  BUF_X1 U27895 ( .A(n33370), .Z(n40090) );
  BUF_X1 U27896 ( .A(n33373), .Z(n40070) );
  BUF_X1 U27897 ( .A(n33376), .Z(n40050) );
  BUF_X1 U27898 ( .A(n33385), .Z(n39992) );
  BUF_X1 U27899 ( .A(n33388), .Z(n39972) );
  BUF_X1 U27900 ( .A(n33409), .Z(n39874) );
  BUF_X1 U27901 ( .A(n33412), .Z(n39854) );
  BUF_X1 U27902 ( .A(n33379), .Z(n40030) );
  BUF_X1 U27903 ( .A(n33382), .Z(n40011) );
  BUF_X1 U27904 ( .A(n33359), .Z(n40129) );
  BUF_X1 U27905 ( .A(n33363), .Z(n40109) );
  BUF_X1 U27906 ( .A(n33418), .Z(n39814) );
  AND2_X1 U27907 ( .A1(n37249), .A2(n37227), .ZN(n36028) );
  AND2_X1 U27908 ( .A1(n37249), .A2(n37229), .ZN(n36029) );
  AND2_X1 U27909 ( .A1(n37249), .A2(n37233), .ZN(n36034) );
  AND2_X1 U27910 ( .A1(n37249), .A2(n37235), .ZN(n36035) );
  AND2_X1 U27911 ( .A1(n34693), .A2(n34671), .ZN(n33473) );
  AND2_X1 U27912 ( .A1(n34693), .A2(n34674), .ZN(n33474) );
  AND2_X1 U27913 ( .A1(n34693), .A2(n34678), .ZN(n33479) );
  AND2_X1 U27914 ( .A1(n34693), .A2(n34680), .ZN(n33480) );
  AND2_X1 U27915 ( .A1(n35967), .A2(n35945), .ZN(n34747) );
  AND2_X1 U27916 ( .A1(n35967), .A2(n35948), .ZN(n34748) );
  AND2_X1 U27917 ( .A1(n35967), .A2(n35952), .ZN(n34753) );
  AND2_X1 U27918 ( .A1(n35967), .A2(n35954), .ZN(n34754) );
  AND2_X1 U27919 ( .A1(n37226), .A2(n37231), .ZN(n35988) );
  AND2_X1 U27920 ( .A1(n37226), .A2(n37230), .ZN(n35989) );
  AND2_X1 U27921 ( .A1(n34676), .A2(n34672), .ZN(n33433) );
  AND2_X1 U27922 ( .A1(n35950), .A2(n35946), .ZN(n34707) );
  AND2_X1 U27923 ( .A1(n37233), .A2(n37239), .ZN(n36017) );
  AND2_X1 U27924 ( .A1(n37230), .A2(n37239), .ZN(n36006) );
  AND2_X1 U27925 ( .A1(n37227), .A2(n37239), .ZN(n36007) );
  AND2_X1 U27926 ( .A1(n34675), .A2(n34672), .ZN(n33434) );
  AND2_X1 U27927 ( .A1(n34675), .A2(n34684), .ZN(n33451) );
  AND2_X1 U27928 ( .A1(n35949), .A2(n35946), .ZN(n34708) );
  AND2_X1 U27929 ( .A1(n35949), .A2(n35958), .ZN(n34725) );
  AND2_X1 U27930 ( .A1(n34673), .A2(n34690), .ZN(n33461) );
  AND2_X1 U27931 ( .A1(n34678), .A2(n34684), .ZN(n33462) );
  AND2_X1 U27932 ( .A1(n34671), .A2(n34684), .ZN(n33452) );
  AND2_X1 U27933 ( .A1(n35947), .A2(n35964), .ZN(n34735) );
  AND2_X1 U27934 ( .A1(n35952), .A2(n35958), .ZN(n34736) );
  AND2_X1 U27935 ( .A1(n35945), .A2(n35958), .ZN(n34726) );
  AND2_X1 U27936 ( .A1(n37246), .A2(n37234), .ZN(n36022) );
  AND2_X1 U27937 ( .A1(n37246), .A2(n37231), .ZN(n36023) );
  AND2_X1 U27938 ( .A1(n34690), .A2(n34679), .ZN(n33467) );
  AND2_X1 U27939 ( .A1(n34690), .A2(n34676), .ZN(n33468) );
  AND2_X1 U27940 ( .A1(n35964), .A2(n35953), .ZN(n34741) );
  AND2_X1 U27941 ( .A1(n35964), .A2(n35950), .ZN(n34742) );
  AND2_X1 U27942 ( .A1(n37236), .A2(n37235), .ZN(n36000) );
  AND2_X1 U27943 ( .A1(n37236), .A2(n37234), .ZN(n36001) );
  AND2_X1 U27944 ( .A1(n37236), .A2(n37229), .ZN(n35994) );
  AND2_X1 U27945 ( .A1(n37236), .A2(n37228), .ZN(n35995) );
  AND2_X1 U27946 ( .A1(n34681), .A2(n34680), .ZN(n33445) );
  AND2_X1 U27947 ( .A1(n34681), .A2(n34679), .ZN(n33446) );
  AND2_X1 U27948 ( .A1(n35955), .A2(n35954), .ZN(n34719) );
  AND2_X1 U27949 ( .A1(n35955), .A2(n35953), .ZN(n34720) );
  AND2_X1 U27950 ( .A1(n34681), .A2(n34673), .ZN(n33440) );
  AND2_X1 U27951 ( .A1(n35955), .A2(n35947), .ZN(n34714) );
  AND2_X1 U27952 ( .A1(n34681), .A2(n34674), .ZN(n33439) );
  AND2_X1 U27953 ( .A1(n35955), .A2(n35948), .ZN(n34713) );
  INV_X1 U27954 ( .A(n33301), .ZN(n32150) );
  NAND2_X1 U27955 ( .A1(n41370), .A2(n35972), .ZN(n35981) );
  INV_X1 U27956 ( .A(n33225), .ZN(n32075) );
  NAND2_X1 U27957 ( .A1(n41370), .A2(n39796), .ZN(n33426) );
  NAND2_X1 U27958 ( .A1(n41370), .A2(n39544), .ZN(n34700) );
  BUF_X1 U27959 ( .A(n40981), .Z(n40984) );
  BUF_X1 U27960 ( .A(n40987), .Z(n40990) );
  BUF_X1 U27961 ( .A(n40993), .Z(n40996) );
  BUF_X1 U27962 ( .A(n40999), .Z(n41002) );
  BUF_X1 U27963 ( .A(n41005), .Z(n41008) );
  BUF_X1 U27964 ( .A(n41011), .Z(n41014) );
  BUF_X1 U27965 ( .A(n41017), .Z(n41020) );
  BUF_X1 U27966 ( .A(n41023), .Z(n41026) );
  BUF_X1 U27967 ( .A(n41029), .Z(n41032) );
  BUF_X1 U27968 ( .A(n41035), .Z(n41038) );
  BUF_X1 U27969 ( .A(n41041), .Z(n41044) );
  BUF_X1 U27970 ( .A(n41047), .Z(n41050) );
  BUF_X1 U27971 ( .A(n41053), .Z(n41056) );
  BUF_X1 U27972 ( .A(n41059), .Z(n41062) );
  BUF_X1 U27973 ( .A(n41065), .Z(n41068) );
  BUF_X1 U27974 ( .A(n41071), .Z(n41074) );
  BUF_X1 U27975 ( .A(n41077), .Z(n41080) );
  BUF_X1 U27976 ( .A(n41083), .Z(n41086) );
  BUF_X1 U27977 ( .A(n41089), .Z(n41092) );
  BUF_X1 U27978 ( .A(n41095), .Z(n41098) );
  BUF_X1 U27979 ( .A(n41101), .Z(n41104) );
  BUF_X1 U27980 ( .A(n41107), .Z(n41110) );
  BUF_X1 U27981 ( .A(n41113), .Z(n41116) );
  BUF_X1 U27982 ( .A(n41119), .Z(n41122) );
  BUF_X1 U27983 ( .A(n41125), .Z(n41128) );
  BUF_X1 U27984 ( .A(n41131), .Z(n41134) );
  BUF_X1 U27985 ( .A(n41137), .Z(n41140) );
  BUF_X1 U27986 ( .A(n41143), .Z(n41146) );
  BUF_X1 U27987 ( .A(n41149), .Z(n41152) );
  BUF_X1 U27988 ( .A(n41155), .Z(n41158) );
  BUF_X1 U27989 ( .A(n41161), .Z(n41164) );
  BUF_X1 U27990 ( .A(n41167), .Z(n41170) );
  BUF_X1 U27991 ( .A(n41173), .Z(n41176) );
  BUF_X1 U27992 ( .A(n41179), .Z(n41182) );
  BUF_X1 U27993 ( .A(n41185), .Z(n41188) );
  BUF_X1 U27994 ( .A(n41191), .Z(n41194) );
  BUF_X1 U27995 ( .A(n41197), .Z(n41200) );
  BUF_X1 U27996 ( .A(n41203), .Z(n41206) );
  BUF_X1 U27997 ( .A(n41209), .Z(n41212) );
  BUF_X1 U27998 ( .A(n41215), .Z(n41218) );
  BUF_X1 U27999 ( .A(n41221), .Z(n41224) );
  BUF_X1 U28000 ( .A(n41227), .Z(n41230) );
  BUF_X1 U28001 ( .A(n41233), .Z(n41236) );
  BUF_X1 U28002 ( .A(n41239), .Z(n41242) );
  BUF_X1 U28003 ( .A(n41245), .Z(n41248) );
  BUF_X1 U28004 ( .A(n41251), .Z(n41254) );
  BUF_X1 U28005 ( .A(n41257), .Z(n41260) );
  BUF_X1 U28006 ( .A(n41263), .Z(n41266) );
  BUF_X1 U28007 ( .A(n41269), .Z(n41272) );
  BUF_X1 U28008 ( .A(n41275), .Z(n41278) );
  BUF_X1 U28009 ( .A(n41281), .Z(n41284) );
  BUF_X1 U28010 ( .A(n41287), .Z(n41290) );
  BUF_X1 U28011 ( .A(n41293), .Z(n41296) );
  BUF_X1 U28012 ( .A(n41299), .Z(n41302) );
  BUF_X1 U28013 ( .A(n41305), .Z(n41308) );
  BUF_X1 U28014 ( .A(n41311), .Z(n41314) );
  BUF_X1 U28015 ( .A(n41317), .Z(n41320) );
  BUF_X1 U28016 ( .A(n41323), .Z(n41326) );
  BUF_X1 U28017 ( .A(n41329), .Z(n41332) );
  BUF_X1 U28018 ( .A(n41335), .Z(n41338) );
  BUF_X1 U28019 ( .A(n41341), .Z(n41344) );
  BUF_X1 U28020 ( .A(n41347), .Z(n41350) );
  BUF_X1 U28021 ( .A(n41353), .Z(n41356) );
  BUF_X1 U28022 ( .A(n41359), .Z(n41362) );
  BUF_X1 U28023 ( .A(n40980), .Z(n40983) );
  BUF_X1 U28024 ( .A(n40986), .Z(n40989) );
  BUF_X1 U28025 ( .A(n40992), .Z(n40995) );
  BUF_X1 U28026 ( .A(n40998), .Z(n41001) );
  BUF_X1 U28027 ( .A(n41004), .Z(n41007) );
  BUF_X1 U28028 ( .A(n41010), .Z(n41013) );
  BUF_X1 U28029 ( .A(n41016), .Z(n41019) );
  BUF_X1 U28030 ( .A(n41022), .Z(n41025) );
  BUF_X1 U28031 ( .A(n41028), .Z(n41031) );
  BUF_X1 U28032 ( .A(n41034), .Z(n41037) );
  BUF_X1 U28033 ( .A(n41040), .Z(n41043) );
  BUF_X1 U28034 ( .A(n41046), .Z(n41049) );
  BUF_X1 U28035 ( .A(n41052), .Z(n41055) );
  BUF_X1 U28036 ( .A(n41058), .Z(n41061) );
  BUF_X1 U28037 ( .A(n41064), .Z(n41067) );
  BUF_X1 U28038 ( .A(n41070), .Z(n41073) );
  BUF_X1 U28039 ( .A(n41076), .Z(n41079) );
  BUF_X1 U28040 ( .A(n41082), .Z(n41085) );
  BUF_X1 U28041 ( .A(n41088), .Z(n41091) );
  BUF_X1 U28042 ( .A(n41094), .Z(n41097) );
  BUF_X1 U28043 ( .A(n41100), .Z(n41103) );
  BUF_X1 U28044 ( .A(n41106), .Z(n41109) );
  BUF_X1 U28045 ( .A(n41112), .Z(n41115) );
  BUF_X1 U28046 ( .A(n41118), .Z(n41121) );
  BUF_X1 U28047 ( .A(n41124), .Z(n41127) );
  BUF_X1 U28048 ( .A(n41130), .Z(n41133) );
  BUF_X1 U28049 ( .A(n41136), .Z(n41139) );
  BUF_X1 U28050 ( .A(n41142), .Z(n41145) );
  BUF_X1 U28051 ( .A(n41148), .Z(n41151) );
  BUF_X1 U28052 ( .A(n41154), .Z(n41157) );
  BUF_X1 U28053 ( .A(n41160), .Z(n41163) );
  BUF_X1 U28054 ( .A(n41166), .Z(n41169) );
  BUF_X1 U28055 ( .A(n41172), .Z(n41175) );
  BUF_X1 U28056 ( .A(n41178), .Z(n41181) );
  BUF_X1 U28057 ( .A(n41184), .Z(n41187) );
  BUF_X1 U28058 ( .A(n41190), .Z(n41193) );
  BUF_X1 U28059 ( .A(n41196), .Z(n41199) );
  BUF_X1 U28060 ( .A(n41202), .Z(n41205) );
  BUF_X1 U28061 ( .A(n41208), .Z(n41211) );
  BUF_X1 U28062 ( .A(n41214), .Z(n41217) );
  BUF_X1 U28063 ( .A(n41220), .Z(n41223) );
  BUF_X1 U28064 ( .A(n41226), .Z(n41229) );
  BUF_X1 U28065 ( .A(n41232), .Z(n41235) );
  BUF_X1 U28066 ( .A(n41238), .Z(n41241) );
  BUF_X1 U28067 ( .A(n41244), .Z(n41247) );
  BUF_X1 U28068 ( .A(n41250), .Z(n41253) );
  BUF_X1 U28069 ( .A(n41256), .Z(n41259) );
  BUF_X1 U28070 ( .A(n41262), .Z(n41265) );
  BUF_X1 U28071 ( .A(n41268), .Z(n41271) );
  BUF_X1 U28072 ( .A(n41274), .Z(n41277) );
  BUF_X1 U28073 ( .A(n41280), .Z(n41283) );
  BUF_X1 U28074 ( .A(n41286), .Z(n41289) );
  BUF_X1 U28075 ( .A(n41292), .Z(n41295) );
  BUF_X1 U28076 ( .A(n41298), .Z(n41301) );
  BUF_X1 U28077 ( .A(n41304), .Z(n41307) );
  BUF_X1 U28078 ( .A(n41310), .Z(n41313) );
  BUF_X1 U28079 ( .A(n41316), .Z(n41319) );
  BUF_X1 U28080 ( .A(n41322), .Z(n41325) );
  BUF_X1 U28081 ( .A(n41328), .Z(n41331) );
  BUF_X1 U28082 ( .A(n41334), .Z(n41337) );
  BUF_X1 U28083 ( .A(n41340), .Z(n41343) );
  BUF_X1 U28084 ( .A(n41346), .Z(n41349) );
  BUF_X1 U28085 ( .A(n41352), .Z(n41355) );
  BUF_X1 U28086 ( .A(n41358), .Z(n41361) );
  BUF_X1 U28087 ( .A(n41118), .Z(n41120) );
  BUF_X1 U28088 ( .A(n41124), .Z(n41126) );
  BUF_X1 U28089 ( .A(n41130), .Z(n41132) );
  BUF_X1 U28090 ( .A(n41136), .Z(n41138) );
  BUF_X1 U28091 ( .A(n41142), .Z(n41144) );
  BUF_X1 U28092 ( .A(n41148), .Z(n41150) );
  BUF_X1 U28093 ( .A(n41154), .Z(n41156) );
  BUF_X1 U28094 ( .A(n41160), .Z(n41162) );
  BUF_X1 U28095 ( .A(n41166), .Z(n41168) );
  BUF_X1 U28096 ( .A(n41172), .Z(n41174) );
  BUF_X1 U28097 ( .A(n41178), .Z(n41180) );
  BUF_X1 U28098 ( .A(n41184), .Z(n41186) );
  BUF_X1 U28099 ( .A(n41190), .Z(n41192) );
  BUF_X1 U28100 ( .A(n41196), .Z(n41198) );
  BUF_X1 U28101 ( .A(n41202), .Z(n41204) );
  BUF_X1 U28102 ( .A(n41208), .Z(n41210) );
  BUF_X1 U28103 ( .A(n41214), .Z(n41216) );
  BUF_X1 U28104 ( .A(n41220), .Z(n41222) );
  BUF_X1 U28105 ( .A(n41226), .Z(n41228) );
  BUF_X1 U28106 ( .A(n41232), .Z(n41234) );
  BUF_X1 U28107 ( .A(n41238), .Z(n41240) );
  BUF_X1 U28108 ( .A(n41244), .Z(n41246) );
  BUF_X1 U28109 ( .A(n41250), .Z(n41252) );
  BUF_X1 U28110 ( .A(n41256), .Z(n41258) );
  BUF_X1 U28111 ( .A(n41262), .Z(n41264) );
  BUF_X1 U28112 ( .A(n41268), .Z(n41270) );
  BUF_X1 U28113 ( .A(n41274), .Z(n41276) );
  BUF_X1 U28114 ( .A(n41280), .Z(n41282) );
  BUF_X1 U28115 ( .A(n41286), .Z(n41288) );
  BUF_X1 U28116 ( .A(n41292), .Z(n41294) );
  BUF_X1 U28117 ( .A(n41298), .Z(n41300) );
  BUF_X1 U28118 ( .A(n41304), .Z(n41306) );
  BUF_X1 U28119 ( .A(n41310), .Z(n41312) );
  BUF_X1 U28120 ( .A(n41316), .Z(n41318) );
  BUF_X1 U28121 ( .A(n41322), .Z(n41324) );
  BUF_X1 U28122 ( .A(n41328), .Z(n41330) );
  BUF_X1 U28123 ( .A(n41334), .Z(n41336) );
  BUF_X1 U28124 ( .A(n41340), .Z(n41342) );
  BUF_X1 U28125 ( .A(n41346), .Z(n41348) );
  BUF_X1 U28126 ( .A(n41352), .Z(n41354) );
  BUF_X1 U28127 ( .A(n41358), .Z(n41360) );
  BUF_X1 U28128 ( .A(n40980), .Z(n40982) );
  BUF_X1 U28129 ( .A(n40986), .Z(n40988) );
  BUF_X1 U28130 ( .A(n40992), .Z(n40994) );
  BUF_X1 U28131 ( .A(n40998), .Z(n41000) );
  BUF_X1 U28132 ( .A(n41004), .Z(n41006) );
  BUF_X1 U28133 ( .A(n41010), .Z(n41012) );
  BUF_X1 U28134 ( .A(n41016), .Z(n41018) );
  BUF_X1 U28135 ( .A(n41022), .Z(n41024) );
  BUF_X1 U28136 ( .A(n41028), .Z(n41030) );
  BUF_X1 U28137 ( .A(n41034), .Z(n41036) );
  BUF_X1 U28138 ( .A(n41040), .Z(n41042) );
  BUF_X1 U28139 ( .A(n41046), .Z(n41048) );
  BUF_X1 U28140 ( .A(n41052), .Z(n41054) );
  BUF_X1 U28141 ( .A(n41058), .Z(n41060) );
  BUF_X1 U28142 ( .A(n41064), .Z(n41066) );
  BUF_X1 U28143 ( .A(n41070), .Z(n41072) );
  BUF_X1 U28144 ( .A(n41076), .Z(n41078) );
  BUF_X1 U28145 ( .A(n41082), .Z(n41084) );
  BUF_X1 U28146 ( .A(n41088), .Z(n41090) );
  BUF_X1 U28147 ( .A(n41094), .Z(n41096) );
  BUF_X1 U28148 ( .A(n41100), .Z(n41102) );
  BUF_X1 U28149 ( .A(n41106), .Z(n41108) );
  BUF_X1 U28150 ( .A(n41112), .Z(n41114) );
  BUF_X1 U28151 ( .A(n40597), .Z(n40600) );
  BUF_X1 U28152 ( .A(n40603), .Z(n40606) );
  BUF_X1 U28153 ( .A(n40609), .Z(n40612) );
  BUF_X1 U28154 ( .A(n40615), .Z(n40618) );
  BUF_X1 U28155 ( .A(n40621), .Z(n40624) );
  BUF_X1 U28156 ( .A(n40627), .Z(n40630) );
  BUF_X1 U28157 ( .A(n40633), .Z(n40636) );
  BUF_X1 U28158 ( .A(n40639), .Z(n40642) );
  BUF_X1 U28159 ( .A(n40645), .Z(n40648) );
  BUF_X1 U28160 ( .A(n40651), .Z(n40654) );
  BUF_X1 U28161 ( .A(n40657), .Z(n40660) );
  BUF_X1 U28162 ( .A(n40663), .Z(n40666) );
  BUF_X1 U28163 ( .A(n40669), .Z(n40672) );
  BUF_X1 U28164 ( .A(n40675), .Z(n40678) );
  BUF_X1 U28165 ( .A(n40681), .Z(n40684) );
  BUF_X1 U28166 ( .A(n40687), .Z(n40690) );
  BUF_X1 U28167 ( .A(n40693), .Z(n40696) );
  BUF_X1 U28168 ( .A(n40699), .Z(n40702) );
  BUF_X1 U28169 ( .A(n40705), .Z(n40708) );
  BUF_X1 U28170 ( .A(n40711), .Z(n40714) );
  BUF_X1 U28171 ( .A(n40717), .Z(n40720) );
  BUF_X1 U28172 ( .A(n40723), .Z(n40726) );
  BUF_X1 U28173 ( .A(n40729), .Z(n40732) );
  BUF_X1 U28174 ( .A(n40735), .Z(n40738) );
  BUF_X1 U28175 ( .A(n40741), .Z(n40744) );
  BUF_X1 U28176 ( .A(n40747), .Z(n40750) );
  BUF_X1 U28177 ( .A(n40753), .Z(n40756) );
  BUF_X1 U28178 ( .A(n40759), .Z(n40762) );
  BUF_X1 U28179 ( .A(n40765), .Z(n40768) );
  BUF_X1 U28180 ( .A(n40771), .Z(n40774) );
  BUF_X1 U28181 ( .A(n40777), .Z(n40780) );
  BUF_X1 U28182 ( .A(n40783), .Z(n40786) );
  BUF_X1 U28183 ( .A(n40789), .Z(n40792) );
  BUF_X1 U28184 ( .A(n40795), .Z(n40798) );
  BUF_X1 U28185 ( .A(n40801), .Z(n40804) );
  BUF_X1 U28186 ( .A(n40807), .Z(n40810) );
  BUF_X1 U28187 ( .A(n40813), .Z(n40816) );
  BUF_X1 U28188 ( .A(n40819), .Z(n40822) );
  BUF_X1 U28189 ( .A(n40825), .Z(n40828) );
  BUF_X1 U28190 ( .A(n40831), .Z(n40834) );
  BUF_X1 U28191 ( .A(n40837), .Z(n40840) );
  BUF_X1 U28192 ( .A(n40843), .Z(n40846) );
  BUF_X1 U28193 ( .A(n40849), .Z(n40852) );
  BUF_X1 U28194 ( .A(n40855), .Z(n40858) );
  BUF_X1 U28195 ( .A(n40861), .Z(n40864) );
  BUF_X1 U28196 ( .A(n40867), .Z(n40870) );
  BUF_X1 U28197 ( .A(n40873), .Z(n40876) );
  BUF_X1 U28198 ( .A(n40879), .Z(n40882) );
  BUF_X1 U28199 ( .A(n40885), .Z(n40888) );
  BUF_X1 U28200 ( .A(n40891), .Z(n40894) );
  BUF_X1 U28201 ( .A(n40897), .Z(n40900) );
  BUF_X1 U28202 ( .A(n40903), .Z(n40906) );
  BUF_X1 U28203 ( .A(n40909), .Z(n40912) );
  BUF_X1 U28204 ( .A(n40915), .Z(n40918) );
  BUF_X1 U28205 ( .A(n40921), .Z(n40924) );
  BUF_X1 U28206 ( .A(n40927), .Z(n40930) );
  BUF_X1 U28207 ( .A(n40933), .Z(n40936) );
  BUF_X1 U28208 ( .A(n40939), .Z(n40942) );
  BUF_X1 U28209 ( .A(n40945), .Z(n40948) );
  BUF_X1 U28210 ( .A(n40951), .Z(n40954) );
  BUF_X1 U28211 ( .A(n40957), .Z(n40960) );
  BUF_X1 U28212 ( .A(n40963), .Z(n40966) );
  BUF_X1 U28213 ( .A(n40969), .Z(n40972) );
  BUF_X1 U28214 ( .A(n40975), .Z(n40978) );
  BUF_X1 U28215 ( .A(n40596), .Z(n40599) );
  BUF_X1 U28216 ( .A(n40602), .Z(n40605) );
  BUF_X1 U28217 ( .A(n40608), .Z(n40611) );
  BUF_X1 U28218 ( .A(n40614), .Z(n40617) );
  BUF_X1 U28219 ( .A(n40620), .Z(n40623) );
  BUF_X1 U28220 ( .A(n40626), .Z(n40629) );
  BUF_X1 U28221 ( .A(n40632), .Z(n40635) );
  BUF_X1 U28222 ( .A(n40638), .Z(n40641) );
  BUF_X1 U28223 ( .A(n40644), .Z(n40647) );
  BUF_X1 U28224 ( .A(n40650), .Z(n40653) );
  BUF_X1 U28225 ( .A(n40656), .Z(n40659) );
  BUF_X1 U28226 ( .A(n40662), .Z(n40665) );
  BUF_X1 U28227 ( .A(n40668), .Z(n40671) );
  BUF_X1 U28228 ( .A(n40674), .Z(n40677) );
  BUF_X1 U28229 ( .A(n40680), .Z(n40683) );
  BUF_X1 U28230 ( .A(n40686), .Z(n40689) );
  BUF_X1 U28231 ( .A(n40692), .Z(n40695) );
  BUF_X1 U28232 ( .A(n40698), .Z(n40701) );
  BUF_X1 U28233 ( .A(n40704), .Z(n40707) );
  BUF_X1 U28234 ( .A(n40710), .Z(n40713) );
  BUF_X1 U28235 ( .A(n40716), .Z(n40719) );
  BUF_X1 U28236 ( .A(n40722), .Z(n40725) );
  BUF_X1 U28237 ( .A(n40728), .Z(n40731) );
  BUF_X1 U28238 ( .A(n40734), .Z(n40737) );
  BUF_X1 U28239 ( .A(n40740), .Z(n40743) );
  BUF_X1 U28240 ( .A(n40746), .Z(n40749) );
  BUF_X1 U28241 ( .A(n40752), .Z(n40755) );
  BUF_X1 U28242 ( .A(n40758), .Z(n40761) );
  BUF_X1 U28243 ( .A(n40764), .Z(n40767) );
  BUF_X1 U28244 ( .A(n40770), .Z(n40773) );
  BUF_X1 U28245 ( .A(n40776), .Z(n40779) );
  BUF_X1 U28246 ( .A(n40782), .Z(n40785) );
  BUF_X1 U28247 ( .A(n40788), .Z(n40791) );
  BUF_X1 U28248 ( .A(n40794), .Z(n40797) );
  BUF_X1 U28249 ( .A(n40800), .Z(n40803) );
  BUF_X1 U28250 ( .A(n40806), .Z(n40809) );
  BUF_X1 U28251 ( .A(n40812), .Z(n40815) );
  BUF_X1 U28252 ( .A(n40818), .Z(n40821) );
  BUF_X1 U28253 ( .A(n40824), .Z(n40827) );
  BUF_X1 U28254 ( .A(n40830), .Z(n40833) );
  BUF_X1 U28255 ( .A(n40836), .Z(n40839) );
  BUF_X1 U28256 ( .A(n40842), .Z(n40845) );
  BUF_X1 U28257 ( .A(n40848), .Z(n40851) );
  BUF_X1 U28258 ( .A(n40854), .Z(n40857) );
  BUF_X1 U28259 ( .A(n40860), .Z(n40863) );
  BUF_X1 U28260 ( .A(n40866), .Z(n40869) );
  BUF_X1 U28261 ( .A(n40872), .Z(n40875) );
  BUF_X1 U28262 ( .A(n40878), .Z(n40881) );
  BUF_X1 U28263 ( .A(n40884), .Z(n40887) );
  BUF_X1 U28264 ( .A(n40890), .Z(n40893) );
  BUF_X1 U28265 ( .A(n40896), .Z(n40899) );
  BUF_X1 U28266 ( .A(n40902), .Z(n40905) );
  BUF_X1 U28267 ( .A(n40908), .Z(n40911) );
  BUF_X1 U28268 ( .A(n40914), .Z(n40917) );
  BUF_X1 U28269 ( .A(n40920), .Z(n40923) );
  BUF_X1 U28270 ( .A(n40926), .Z(n40929) );
  BUF_X1 U28271 ( .A(n40932), .Z(n40935) );
  BUF_X1 U28272 ( .A(n40938), .Z(n40941) );
  BUF_X1 U28273 ( .A(n40944), .Z(n40947) );
  BUF_X1 U28274 ( .A(n40950), .Z(n40953) );
  BUF_X1 U28275 ( .A(n40956), .Z(n40959) );
  BUF_X1 U28276 ( .A(n40962), .Z(n40965) );
  BUF_X1 U28277 ( .A(n40968), .Z(n40971) );
  BUF_X1 U28278 ( .A(n40974), .Z(n40977) );
  BUF_X1 U28279 ( .A(n40734), .Z(n40736) );
  BUF_X1 U28280 ( .A(n40740), .Z(n40742) );
  BUF_X1 U28281 ( .A(n40746), .Z(n40748) );
  BUF_X1 U28282 ( .A(n40752), .Z(n40754) );
  BUF_X1 U28283 ( .A(n40758), .Z(n40760) );
  BUF_X1 U28284 ( .A(n40764), .Z(n40766) );
  BUF_X1 U28285 ( .A(n40770), .Z(n40772) );
  BUF_X1 U28286 ( .A(n40776), .Z(n40778) );
  BUF_X1 U28287 ( .A(n40782), .Z(n40784) );
  BUF_X1 U28288 ( .A(n40788), .Z(n40790) );
  BUF_X1 U28289 ( .A(n40794), .Z(n40796) );
  BUF_X1 U28290 ( .A(n40800), .Z(n40802) );
  BUF_X1 U28291 ( .A(n40806), .Z(n40808) );
  BUF_X1 U28292 ( .A(n40812), .Z(n40814) );
  BUF_X1 U28293 ( .A(n40818), .Z(n40820) );
  BUF_X1 U28294 ( .A(n40824), .Z(n40826) );
  BUF_X1 U28295 ( .A(n40830), .Z(n40832) );
  BUF_X1 U28296 ( .A(n40836), .Z(n40838) );
  BUF_X1 U28297 ( .A(n40842), .Z(n40844) );
  BUF_X1 U28298 ( .A(n40848), .Z(n40850) );
  BUF_X1 U28299 ( .A(n40854), .Z(n40856) );
  BUF_X1 U28300 ( .A(n40860), .Z(n40862) );
  BUF_X1 U28301 ( .A(n40866), .Z(n40868) );
  BUF_X1 U28302 ( .A(n40872), .Z(n40874) );
  BUF_X1 U28303 ( .A(n40878), .Z(n40880) );
  BUF_X1 U28304 ( .A(n40884), .Z(n40886) );
  BUF_X1 U28305 ( .A(n40890), .Z(n40892) );
  BUF_X1 U28306 ( .A(n40896), .Z(n40898) );
  BUF_X1 U28307 ( .A(n40902), .Z(n40904) );
  BUF_X1 U28308 ( .A(n40908), .Z(n40910) );
  BUF_X1 U28309 ( .A(n40914), .Z(n40916) );
  BUF_X1 U28310 ( .A(n40920), .Z(n40922) );
  BUF_X1 U28311 ( .A(n40926), .Z(n40928) );
  BUF_X1 U28312 ( .A(n40932), .Z(n40934) );
  BUF_X1 U28313 ( .A(n40938), .Z(n40940) );
  BUF_X1 U28314 ( .A(n40944), .Z(n40946) );
  BUF_X1 U28315 ( .A(n40950), .Z(n40952) );
  BUF_X1 U28316 ( .A(n40956), .Z(n40958) );
  BUF_X1 U28317 ( .A(n40962), .Z(n40964) );
  BUF_X1 U28318 ( .A(n40968), .Z(n40970) );
  BUF_X1 U28319 ( .A(n40974), .Z(n40976) );
  BUF_X1 U28320 ( .A(n40596), .Z(n40598) );
  BUF_X1 U28321 ( .A(n40602), .Z(n40604) );
  BUF_X1 U28322 ( .A(n40608), .Z(n40610) );
  BUF_X1 U28323 ( .A(n40614), .Z(n40616) );
  BUF_X1 U28324 ( .A(n40620), .Z(n40622) );
  BUF_X1 U28325 ( .A(n40626), .Z(n40628) );
  BUF_X1 U28326 ( .A(n40632), .Z(n40634) );
  BUF_X1 U28327 ( .A(n40638), .Z(n40640) );
  BUF_X1 U28328 ( .A(n40644), .Z(n40646) );
  BUF_X1 U28329 ( .A(n40650), .Z(n40652) );
  BUF_X1 U28330 ( .A(n40656), .Z(n40658) );
  BUF_X1 U28331 ( .A(n40662), .Z(n40664) );
  BUF_X1 U28332 ( .A(n40668), .Z(n40670) );
  BUF_X1 U28333 ( .A(n40674), .Z(n40676) );
  BUF_X1 U28334 ( .A(n40680), .Z(n40682) );
  BUF_X1 U28335 ( .A(n40686), .Z(n40688) );
  BUF_X1 U28336 ( .A(n40692), .Z(n40694) );
  BUF_X1 U28337 ( .A(n40698), .Z(n40700) );
  BUF_X1 U28338 ( .A(n40704), .Z(n40706) );
  BUF_X1 U28339 ( .A(n40710), .Z(n40712) );
  BUF_X1 U28340 ( .A(n40716), .Z(n40718) );
  BUF_X1 U28341 ( .A(n40722), .Z(n40724) );
  BUF_X1 U28342 ( .A(n40728), .Z(n40730) );
  BUF_X1 U28343 ( .A(n40981), .Z(n40985) );
  BUF_X1 U28344 ( .A(n40987), .Z(n40991) );
  BUF_X1 U28345 ( .A(n40993), .Z(n40997) );
  BUF_X1 U28346 ( .A(n40999), .Z(n41003) );
  BUF_X1 U28347 ( .A(n41005), .Z(n41009) );
  BUF_X1 U28348 ( .A(n41011), .Z(n41015) );
  BUF_X1 U28349 ( .A(n41017), .Z(n41021) );
  BUF_X1 U28350 ( .A(n41023), .Z(n41027) );
  BUF_X1 U28351 ( .A(n41029), .Z(n41033) );
  BUF_X1 U28352 ( .A(n41035), .Z(n41039) );
  BUF_X1 U28353 ( .A(n41041), .Z(n41045) );
  BUF_X1 U28354 ( .A(n41047), .Z(n41051) );
  BUF_X1 U28355 ( .A(n41053), .Z(n41057) );
  BUF_X1 U28356 ( .A(n41059), .Z(n41063) );
  BUF_X1 U28357 ( .A(n41065), .Z(n41069) );
  BUF_X1 U28358 ( .A(n41071), .Z(n41075) );
  BUF_X1 U28359 ( .A(n41077), .Z(n41081) );
  BUF_X1 U28360 ( .A(n41083), .Z(n41087) );
  BUF_X1 U28361 ( .A(n41089), .Z(n41093) );
  BUF_X1 U28362 ( .A(n41095), .Z(n41099) );
  BUF_X1 U28363 ( .A(n41101), .Z(n41105) );
  BUF_X1 U28364 ( .A(n41107), .Z(n41111) );
  BUF_X1 U28365 ( .A(n41113), .Z(n41117) );
  BUF_X1 U28366 ( .A(n41119), .Z(n41123) );
  BUF_X1 U28367 ( .A(n41125), .Z(n41129) );
  BUF_X1 U28368 ( .A(n41131), .Z(n41135) );
  BUF_X1 U28369 ( .A(n41137), .Z(n41141) );
  BUF_X1 U28370 ( .A(n41143), .Z(n41147) );
  BUF_X1 U28371 ( .A(n41149), .Z(n41153) );
  BUF_X1 U28372 ( .A(n41155), .Z(n41159) );
  BUF_X1 U28373 ( .A(n41161), .Z(n41165) );
  BUF_X1 U28374 ( .A(n41167), .Z(n41171) );
  BUF_X1 U28375 ( .A(n41173), .Z(n41177) );
  BUF_X1 U28376 ( .A(n41179), .Z(n41183) );
  BUF_X1 U28377 ( .A(n41185), .Z(n41189) );
  BUF_X1 U28378 ( .A(n41191), .Z(n41195) );
  BUF_X1 U28379 ( .A(n41197), .Z(n41201) );
  BUF_X1 U28380 ( .A(n41203), .Z(n41207) );
  BUF_X1 U28381 ( .A(n41209), .Z(n41213) );
  BUF_X1 U28382 ( .A(n41215), .Z(n41219) );
  BUF_X1 U28383 ( .A(n41221), .Z(n41225) );
  BUF_X1 U28384 ( .A(n41227), .Z(n41231) );
  BUF_X1 U28385 ( .A(n41233), .Z(n41237) );
  BUF_X1 U28386 ( .A(n41239), .Z(n41243) );
  BUF_X1 U28387 ( .A(n41245), .Z(n41249) );
  BUF_X1 U28388 ( .A(n41251), .Z(n41255) );
  BUF_X1 U28389 ( .A(n41257), .Z(n41261) );
  BUF_X1 U28390 ( .A(n41263), .Z(n41267) );
  BUF_X1 U28391 ( .A(n41269), .Z(n41273) );
  BUF_X1 U28392 ( .A(n41275), .Z(n41279) );
  BUF_X1 U28393 ( .A(n41281), .Z(n41285) );
  BUF_X1 U28394 ( .A(n41287), .Z(n41291) );
  BUF_X1 U28395 ( .A(n41293), .Z(n41297) );
  BUF_X1 U28396 ( .A(n41299), .Z(n41303) );
  BUF_X1 U28397 ( .A(n41305), .Z(n41309) );
  BUF_X1 U28398 ( .A(n41311), .Z(n41315) );
  BUF_X1 U28399 ( .A(n41317), .Z(n41321) );
  BUF_X1 U28400 ( .A(n41323), .Z(n41327) );
  BUF_X1 U28401 ( .A(n41329), .Z(n41333) );
  BUF_X1 U28402 ( .A(n41335), .Z(n41339) );
  BUF_X1 U28403 ( .A(n41341), .Z(n41345) );
  BUF_X1 U28404 ( .A(n41347), .Z(n41351) );
  BUF_X1 U28405 ( .A(n41353), .Z(n41357) );
  BUF_X1 U28406 ( .A(n41359), .Z(n41363) );
  BUF_X1 U28407 ( .A(n40597), .Z(n40601) );
  BUF_X1 U28408 ( .A(n40603), .Z(n40607) );
  BUF_X1 U28409 ( .A(n40609), .Z(n40613) );
  BUF_X1 U28410 ( .A(n40615), .Z(n40619) );
  BUF_X1 U28411 ( .A(n40621), .Z(n40625) );
  BUF_X1 U28412 ( .A(n40627), .Z(n40631) );
  BUF_X1 U28413 ( .A(n40633), .Z(n40637) );
  BUF_X1 U28414 ( .A(n40639), .Z(n40643) );
  BUF_X1 U28415 ( .A(n40645), .Z(n40649) );
  BUF_X1 U28416 ( .A(n40651), .Z(n40655) );
  BUF_X1 U28417 ( .A(n40657), .Z(n40661) );
  BUF_X1 U28418 ( .A(n40663), .Z(n40667) );
  BUF_X1 U28419 ( .A(n40669), .Z(n40673) );
  BUF_X1 U28420 ( .A(n40675), .Z(n40679) );
  BUF_X1 U28421 ( .A(n40681), .Z(n40685) );
  BUF_X1 U28422 ( .A(n40687), .Z(n40691) );
  BUF_X1 U28423 ( .A(n40693), .Z(n40697) );
  BUF_X1 U28424 ( .A(n40699), .Z(n40703) );
  BUF_X1 U28425 ( .A(n40705), .Z(n40709) );
  BUF_X1 U28426 ( .A(n40711), .Z(n40715) );
  BUF_X1 U28427 ( .A(n40717), .Z(n40721) );
  BUF_X1 U28428 ( .A(n40723), .Z(n40727) );
  BUF_X1 U28429 ( .A(n40729), .Z(n40733) );
  BUF_X1 U28430 ( .A(n40735), .Z(n40739) );
  BUF_X1 U28431 ( .A(n40741), .Z(n40745) );
  BUF_X1 U28432 ( .A(n40747), .Z(n40751) );
  BUF_X1 U28433 ( .A(n40753), .Z(n40757) );
  BUF_X1 U28434 ( .A(n40759), .Z(n40763) );
  BUF_X1 U28435 ( .A(n40765), .Z(n40769) );
  BUF_X1 U28436 ( .A(n40771), .Z(n40775) );
  BUF_X1 U28437 ( .A(n40777), .Z(n40781) );
  BUF_X1 U28438 ( .A(n40783), .Z(n40787) );
  BUF_X1 U28439 ( .A(n40789), .Z(n40793) );
  BUF_X1 U28440 ( .A(n40795), .Z(n40799) );
  BUF_X1 U28441 ( .A(n40801), .Z(n40805) );
  BUF_X1 U28442 ( .A(n40807), .Z(n40811) );
  BUF_X1 U28443 ( .A(n40813), .Z(n40817) );
  BUF_X1 U28444 ( .A(n40819), .Z(n40823) );
  BUF_X1 U28445 ( .A(n40825), .Z(n40829) );
  BUF_X1 U28446 ( .A(n40831), .Z(n40835) );
  BUF_X1 U28447 ( .A(n40837), .Z(n40841) );
  BUF_X1 U28448 ( .A(n40843), .Z(n40847) );
  BUF_X1 U28449 ( .A(n40849), .Z(n40853) );
  BUF_X1 U28450 ( .A(n40855), .Z(n40859) );
  BUF_X1 U28451 ( .A(n40861), .Z(n40865) );
  BUF_X1 U28452 ( .A(n40867), .Z(n40871) );
  BUF_X1 U28453 ( .A(n40873), .Z(n40877) );
  BUF_X1 U28454 ( .A(n40879), .Z(n40883) );
  BUF_X1 U28455 ( .A(n40885), .Z(n40889) );
  BUF_X1 U28456 ( .A(n40891), .Z(n40895) );
  BUF_X1 U28457 ( .A(n40897), .Z(n40901) );
  BUF_X1 U28458 ( .A(n40903), .Z(n40907) );
  BUF_X1 U28459 ( .A(n40909), .Z(n40913) );
  BUF_X1 U28460 ( .A(n40915), .Z(n40919) );
  BUF_X1 U28461 ( .A(n40921), .Z(n40925) );
  BUF_X1 U28462 ( .A(n40927), .Z(n40931) );
  BUF_X1 U28463 ( .A(n40933), .Z(n40937) );
  BUF_X1 U28464 ( .A(n40939), .Z(n40943) );
  BUF_X1 U28465 ( .A(n40945), .Z(n40949) );
  BUF_X1 U28466 ( .A(n40951), .Z(n40955) );
  BUF_X1 U28467 ( .A(n40957), .Z(n40961) );
  BUF_X1 U28468 ( .A(n40963), .Z(n40967) );
  BUF_X1 U28469 ( .A(n40969), .Z(n40973) );
  BUF_X1 U28470 ( .A(n40975), .Z(n40979) );
  NAND2_X1 U28471 ( .A1(n32244), .A2(n33208), .ZN(n34697) );
  NAND2_X1 U28472 ( .A1(n32244), .A2(n33207), .ZN(n35971) );
  OAI221_X1 U28473 ( .B1(n33258), .B2(n33274), .C1(n33259), .C2(n33275), .A(
        n41364), .ZN(n33273) );
  OAI221_X1 U28474 ( .B1(n33258), .B2(n33264), .C1(n33259), .C2(n33265), .A(
        n41364), .ZN(n33263) );
  OAI221_X1 U28475 ( .B1(n33258), .B2(n33269), .C1(n33259), .C2(n33270), .A(
        n41364), .ZN(n33268) );
  OAI221_X1 U28476 ( .B1(n33258), .B2(n32157), .C1(n33259), .C2(n33280), .A(
        n41365), .ZN(n33278) );
  OAI221_X1 U28477 ( .B1(n33258), .B2(n33255), .C1(n33259), .C2(n33260), .A(
        n41364), .ZN(n33254) );
  OAI221_X1 U28478 ( .B1(n33258), .B2(n32158), .C1(n33259), .C2(n33285), .A(
        n41364), .ZN(n33283) );
  OAI221_X1 U28479 ( .B1(n33258), .B2(n32159), .C1(n33259), .C2(n33290), .A(
        n41365), .ZN(n33288) );
  OAI221_X1 U28480 ( .B1(n33258), .B2(n32160), .C1(n33259), .C2(n33296), .A(
        n41365), .ZN(n33293) );
  NOR3_X1 U28481 ( .A1(n32254), .A2(N689), .A3(n32251), .ZN(n37231) );
  NOR3_X1 U28482 ( .A1(n34694), .A2(N6271), .A3(n32166), .ZN(n34676) );
  NOR3_X1 U28483 ( .A1(n35968), .A2(N6396), .A3(n32171), .ZN(n35950) );
  NOR3_X1 U28484 ( .A1(n33398), .A2(N689), .A3(n32251), .ZN(n37234) );
  NOR3_X1 U28485 ( .A1(N688), .A2(N689), .A3(n32254), .ZN(n37235) );
  NOR3_X1 U28486 ( .A1(n33398), .A2(N688), .A3(n32248), .ZN(n37230) );
  NOR3_X1 U28487 ( .A1(N688), .A2(N689), .A3(n33398), .ZN(n37233) );
  NOR3_X1 U28488 ( .A1(n32254), .A2(N688), .A3(n32248), .ZN(n37227) );
  NOR3_X1 U28489 ( .A1(n32168), .A2(N6270), .A3(n32165), .ZN(n34675) );
  NOR3_X1 U28490 ( .A1(n32173), .A2(N6395), .A3(n32170), .ZN(n35949) );
  NOR3_X1 U28491 ( .A1(n33398), .A2(n32251), .A3(n32248), .ZN(n37229) );
  NOR3_X1 U28492 ( .A1(n32166), .A2(N6271), .A3(n32168), .ZN(n34679) );
  NOR3_X1 U28493 ( .A1(n32171), .A2(N6396), .A3(n32173), .ZN(n35953) );
  NOR3_X1 U28494 ( .A1(N6270), .A2(N6271), .A3(n34694), .ZN(n34680) );
  NOR3_X1 U28495 ( .A1(N6395), .A2(N6396), .A3(n35968), .ZN(n35954) );
  NOR3_X1 U28496 ( .A1(N6270), .A2(N6271), .A3(n32168), .ZN(n34678) );
  NOR3_X1 U28497 ( .A1(n34694), .A2(N6270), .A3(n32165), .ZN(n34671) );
  NOR3_X1 U28498 ( .A1(N6395), .A2(N6396), .A3(n32173), .ZN(n35952) );
  NOR3_X1 U28499 ( .A1(n35968), .A2(N6395), .A3(n32170), .ZN(n35945) );
  NOR3_X1 U28500 ( .A1(n32166), .A2(n34694), .A3(n32165), .ZN(n34673) );
  NOR3_X1 U28501 ( .A1(n32171), .A2(n35968), .A3(n32170), .ZN(n35947) );
  NOR2_X1 U28502 ( .A1(n37240), .A2(N690), .ZN(n37239) );
  NOR2_X1 U28503 ( .A1(n32164), .A2(N6273), .ZN(n34690) );
  NOR2_X1 U28504 ( .A1(n32169), .A2(N6398), .ZN(n35964) );
  NOR3_X1 U28505 ( .A1(N929), .A2(N930), .A3(n33402), .ZN(n33289) );
  NOR3_X1 U28506 ( .A1(n33402), .A2(N930), .A3(n32161), .ZN(n33279) );
  NOR3_X1 U28507 ( .A1(n32161), .A2(N930), .A3(n32163), .ZN(n33284) );
  NOR3_X1 U28508 ( .A1(N929), .A2(N930), .A3(n32163), .ZN(n33295) );
  NOR2_X1 U28509 ( .A1(n32246), .A2(n37240), .ZN(n37236) );
  NAND2_X1 U28510 ( .A1(n32244), .A2(n33209), .ZN(n33422) );
  NAND3_X1 U28511 ( .A1(N929), .A2(n32163), .A3(N930), .ZN(n33255) );
  AOI221_X1 U28512 ( .B1(n39638), .B2(n32822), .C1(n39632), .C2(n32774), .A(
        n33558), .ZN(n33555) );
  OAI222_X1 U28513 ( .A1(n30988), .A2(n39626), .B1(n31052), .B2(n39620), .C1(
        n30924), .C2(n39614), .ZN(n33558) );
  AOI221_X1 U28514 ( .B1(n39386), .B2(n32822), .C1(n39380), .C2(n32774), .A(
        n34832), .ZN(n34829) );
  OAI222_X1 U28515 ( .A1(n30988), .A2(n39374), .B1(n31052), .B2(n39368), .C1(
        n30924), .C2(n39362), .ZN(n34832) );
  AOI221_X1 U28516 ( .B1(n39638), .B2(n32821), .C1(n39632), .C2(n32773), .A(
        n33577), .ZN(n33574) );
  OAI222_X1 U28517 ( .A1(n30987), .A2(n39626), .B1(n31051), .B2(n39620), .C1(
        n30923), .C2(n39614), .ZN(n33577) );
  AOI221_X1 U28518 ( .B1(n39386), .B2(n32821), .C1(n39380), .C2(n32773), .A(
        n34851), .ZN(n34848) );
  OAI222_X1 U28519 ( .A1(n30987), .A2(n39374), .B1(n31051), .B2(n39368), .C1(
        n30923), .C2(n39362), .ZN(n34851) );
  AOI221_X1 U28520 ( .B1(n39638), .B2(n32820), .C1(n39632), .C2(n32772), .A(
        n33596), .ZN(n33593) );
  OAI222_X1 U28521 ( .A1(n30986), .A2(n39626), .B1(n31050), .B2(n39620), .C1(
        n30922), .C2(n39614), .ZN(n33596) );
  AOI221_X1 U28522 ( .B1(n39386), .B2(n32820), .C1(n39380), .C2(n32772), .A(
        n34870), .ZN(n34867) );
  OAI222_X1 U28523 ( .A1(n30986), .A2(n39374), .B1(n31050), .B2(n39368), .C1(
        n30922), .C2(n39362), .ZN(n34870) );
  AOI221_X1 U28524 ( .B1(n39638), .B2(n32819), .C1(n39632), .C2(n32771), .A(
        n33615), .ZN(n33612) );
  OAI222_X1 U28525 ( .A1(n30985), .A2(n39626), .B1(n31049), .B2(n39620), .C1(
        n30921), .C2(n39614), .ZN(n33615) );
  AOI221_X1 U28526 ( .B1(n39386), .B2(n32819), .C1(n39380), .C2(n32771), .A(
        n34889), .ZN(n34886) );
  OAI222_X1 U28527 ( .A1(n30985), .A2(n39374), .B1(n31049), .B2(n39368), .C1(
        n30921), .C2(n39362), .ZN(n34889) );
  AOI221_X1 U28528 ( .B1(n39638), .B2(n32818), .C1(n39632), .C2(n32770), .A(
        n33634), .ZN(n33631) );
  OAI222_X1 U28529 ( .A1(n30984), .A2(n39626), .B1(n31048), .B2(n39620), .C1(
        n30920), .C2(n39614), .ZN(n33634) );
  AOI221_X1 U28530 ( .B1(n39386), .B2(n32818), .C1(n39380), .C2(n32770), .A(
        n34908), .ZN(n34905) );
  OAI222_X1 U28531 ( .A1(n30984), .A2(n39374), .B1(n31048), .B2(n39368), .C1(
        n30920), .C2(n39362), .ZN(n34908) );
  AOI221_X1 U28532 ( .B1(n39638), .B2(n32817), .C1(n39632), .C2(n32769), .A(
        n33653), .ZN(n33650) );
  OAI222_X1 U28533 ( .A1(n30983), .A2(n39626), .B1(n31047), .B2(n39620), .C1(
        n30919), .C2(n39614), .ZN(n33653) );
  AOI221_X1 U28534 ( .B1(n39386), .B2(n32817), .C1(n39380), .C2(n32769), .A(
        n34927), .ZN(n34924) );
  OAI222_X1 U28535 ( .A1(n30983), .A2(n39374), .B1(n31047), .B2(n39368), .C1(
        n30919), .C2(n39362), .ZN(n34927) );
  AOI221_X1 U28536 ( .B1(n39638), .B2(n32816), .C1(n39632), .C2(n32768), .A(
        n33672), .ZN(n33669) );
  OAI222_X1 U28537 ( .A1(n30982), .A2(n39626), .B1(n31046), .B2(n39620), .C1(
        n30918), .C2(n39614), .ZN(n33672) );
  AOI221_X1 U28538 ( .B1(n39386), .B2(n32816), .C1(n39380), .C2(n32768), .A(
        n34946), .ZN(n34943) );
  OAI222_X1 U28539 ( .A1(n30982), .A2(n39374), .B1(n31046), .B2(n39368), .C1(
        n30918), .C2(n39362), .ZN(n34946) );
  AOI221_X1 U28540 ( .B1(n39638), .B2(n32815), .C1(n39632), .C2(n32767), .A(
        n33691), .ZN(n33688) );
  OAI222_X1 U28541 ( .A1(n30981), .A2(n39626), .B1(n31045), .B2(n39620), .C1(
        n30917), .C2(n39614), .ZN(n33691) );
  AOI221_X1 U28542 ( .B1(n39386), .B2(n32815), .C1(n39380), .C2(n32767), .A(
        n34965), .ZN(n34962) );
  OAI222_X1 U28543 ( .A1(n30981), .A2(n39374), .B1(n31045), .B2(n39368), .C1(
        n30917), .C2(n39362), .ZN(n34965) );
  AOI221_X1 U28544 ( .B1(n39638), .B2(n32814), .C1(n39632), .C2(n32766), .A(
        n33710), .ZN(n33707) );
  OAI222_X1 U28545 ( .A1(n30980), .A2(n39626), .B1(n31044), .B2(n39620), .C1(
        n30916), .C2(n39614), .ZN(n33710) );
  AOI221_X1 U28546 ( .B1(n39386), .B2(n32814), .C1(n39380), .C2(n32766), .A(
        n34984), .ZN(n34981) );
  OAI222_X1 U28547 ( .A1(n30980), .A2(n39374), .B1(n31044), .B2(n39368), .C1(
        n30916), .C2(n39362), .ZN(n34984) );
  AOI221_X1 U28548 ( .B1(n39638), .B2(n32813), .C1(n39632), .C2(n32765), .A(
        n33729), .ZN(n33726) );
  OAI222_X1 U28549 ( .A1(n30979), .A2(n39626), .B1(n31043), .B2(n39620), .C1(
        n30915), .C2(n39614), .ZN(n33729) );
  AOI221_X1 U28550 ( .B1(n39386), .B2(n32813), .C1(n39380), .C2(n32765), .A(
        n35003), .ZN(n35000) );
  OAI222_X1 U28551 ( .A1(n30979), .A2(n39374), .B1(n31043), .B2(n39368), .C1(
        n30915), .C2(n39362), .ZN(n35003) );
  AOI221_X1 U28552 ( .B1(n39638), .B2(n32812), .C1(n39632), .C2(n32764), .A(
        n33748), .ZN(n33745) );
  OAI222_X1 U28553 ( .A1(n30978), .A2(n39626), .B1(n31042), .B2(n39620), .C1(
        n30914), .C2(n39614), .ZN(n33748) );
  AOI221_X1 U28554 ( .B1(n39386), .B2(n32812), .C1(n39380), .C2(n32764), .A(
        n35022), .ZN(n35019) );
  OAI222_X1 U28555 ( .A1(n30978), .A2(n39374), .B1(n31042), .B2(n39368), .C1(
        n30914), .C2(n39362), .ZN(n35022) );
  AOI221_X1 U28556 ( .B1(n39638), .B2(n32811), .C1(n39632), .C2(n32763), .A(
        n33767), .ZN(n33764) );
  OAI222_X1 U28557 ( .A1(n30977), .A2(n39626), .B1(n31041), .B2(n39620), .C1(
        n30913), .C2(n39614), .ZN(n33767) );
  AOI221_X1 U28558 ( .B1(n39386), .B2(n32811), .C1(n39380), .C2(n32763), .A(
        n35041), .ZN(n35038) );
  OAI222_X1 U28559 ( .A1(n30977), .A2(n39374), .B1(n31041), .B2(n39368), .C1(
        n30913), .C2(n39362), .ZN(n35041) );
  AOI221_X1 U28560 ( .B1(n39637), .B2(n32810), .C1(n39631), .C2(n32762), .A(
        n33786), .ZN(n33783) );
  OAI222_X1 U28561 ( .A1(n30976), .A2(n39625), .B1(n31040), .B2(n39619), .C1(
        n30912), .C2(n39613), .ZN(n33786) );
  AOI221_X1 U28562 ( .B1(n39385), .B2(n32810), .C1(n39379), .C2(n32762), .A(
        n35060), .ZN(n35057) );
  OAI222_X1 U28563 ( .A1(n30976), .A2(n39373), .B1(n31040), .B2(n39367), .C1(
        n30912), .C2(n39361), .ZN(n35060) );
  AOI221_X1 U28564 ( .B1(n39637), .B2(n32809), .C1(n39631), .C2(n32761), .A(
        n33805), .ZN(n33802) );
  OAI222_X1 U28565 ( .A1(n30975), .A2(n39625), .B1(n31039), .B2(n39619), .C1(
        n30911), .C2(n39613), .ZN(n33805) );
  AOI221_X1 U28566 ( .B1(n39385), .B2(n32809), .C1(n39379), .C2(n32761), .A(
        n35079), .ZN(n35076) );
  OAI222_X1 U28567 ( .A1(n30975), .A2(n39373), .B1(n31039), .B2(n39367), .C1(
        n30911), .C2(n39361), .ZN(n35079) );
  AOI221_X1 U28568 ( .B1(n39637), .B2(n32808), .C1(n39631), .C2(n32760), .A(
        n33824), .ZN(n33821) );
  OAI222_X1 U28569 ( .A1(n30974), .A2(n39625), .B1(n31038), .B2(n39619), .C1(
        n30910), .C2(n39613), .ZN(n33824) );
  AOI221_X1 U28570 ( .B1(n39385), .B2(n32808), .C1(n39379), .C2(n32760), .A(
        n35098), .ZN(n35095) );
  OAI222_X1 U28571 ( .A1(n30974), .A2(n39373), .B1(n31038), .B2(n39367), .C1(
        n30910), .C2(n39361), .ZN(n35098) );
  AOI221_X1 U28572 ( .B1(n39637), .B2(n32807), .C1(n39631), .C2(n32759), .A(
        n33843), .ZN(n33840) );
  OAI222_X1 U28573 ( .A1(n30973), .A2(n39625), .B1(n31037), .B2(n39619), .C1(
        n30909), .C2(n39613), .ZN(n33843) );
  AOI221_X1 U28574 ( .B1(n39385), .B2(n32807), .C1(n39379), .C2(n32759), .A(
        n35117), .ZN(n35114) );
  OAI222_X1 U28575 ( .A1(n30973), .A2(n39373), .B1(n31037), .B2(n39367), .C1(
        n30909), .C2(n39361), .ZN(n35117) );
  AOI221_X1 U28576 ( .B1(n39637), .B2(n32806), .C1(n39631), .C2(n32758), .A(
        n33862), .ZN(n33859) );
  OAI222_X1 U28577 ( .A1(n30972), .A2(n39625), .B1(n31036), .B2(n39619), .C1(
        n30908), .C2(n39613), .ZN(n33862) );
  AOI221_X1 U28578 ( .B1(n39385), .B2(n32806), .C1(n39379), .C2(n32758), .A(
        n35136), .ZN(n35133) );
  OAI222_X1 U28579 ( .A1(n30972), .A2(n39373), .B1(n31036), .B2(n39367), .C1(
        n30908), .C2(n39361), .ZN(n35136) );
  AOI221_X1 U28580 ( .B1(n39637), .B2(n32805), .C1(n39631), .C2(n32757), .A(
        n33881), .ZN(n33878) );
  OAI222_X1 U28581 ( .A1(n30971), .A2(n39625), .B1(n31035), .B2(n39619), .C1(
        n30907), .C2(n39613), .ZN(n33881) );
  AOI221_X1 U28582 ( .B1(n39385), .B2(n32805), .C1(n39379), .C2(n32757), .A(
        n35155), .ZN(n35152) );
  OAI222_X1 U28583 ( .A1(n30971), .A2(n39373), .B1(n31035), .B2(n39367), .C1(
        n30907), .C2(n39361), .ZN(n35155) );
  AOI221_X1 U28584 ( .B1(n39637), .B2(n32804), .C1(n39631), .C2(n32756), .A(
        n33900), .ZN(n33897) );
  OAI222_X1 U28585 ( .A1(n30970), .A2(n39625), .B1(n31034), .B2(n39619), .C1(
        n30906), .C2(n39613), .ZN(n33900) );
  AOI221_X1 U28586 ( .B1(n39385), .B2(n32804), .C1(n39379), .C2(n32756), .A(
        n35174), .ZN(n35171) );
  OAI222_X1 U28587 ( .A1(n30970), .A2(n39373), .B1(n31034), .B2(n39367), .C1(
        n30906), .C2(n39361), .ZN(n35174) );
  AOI221_X1 U28588 ( .B1(n39637), .B2(n32803), .C1(n39631), .C2(n32755), .A(
        n33919), .ZN(n33916) );
  OAI222_X1 U28589 ( .A1(n30969), .A2(n39625), .B1(n31033), .B2(n39619), .C1(
        n30905), .C2(n39613), .ZN(n33919) );
  AOI221_X1 U28590 ( .B1(n39385), .B2(n32803), .C1(n39379), .C2(n32755), .A(
        n35193), .ZN(n35190) );
  OAI222_X1 U28591 ( .A1(n30969), .A2(n39373), .B1(n31033), .B2(n39367), .C1(
        n30905), .C2(n39361), .ZN(n35193) );
  AOI221_X1 U28592 ( .B1(n39637), .B2(n32802), .C1(n39631), .C2(n32754), .A(
        n33938), .ZN(n33935) );
  OAI222_X1 U28593 ( .A1(n30968), .A2(n39625), .B1(n31032), .B2(n39619), .C1(
        n30904), .C2(n39613), .ZN(n33938) );
  AOI221_X1 U28594 ( .B1(n39385), .B2(n32802), .C1(n39379), .C2(n32754), .A(
        n35212), .ZN(n35209) );
  OAI222_X1 U28595 ( .A1(n30968), .A2(n39373), .B1(n31032), .B2(n39367), .C1(
        n30904), .C2(n39361), .ZN(n35212) );
  AOI221_X1 U28596 ( .B1(n39637), .B2(n32801), .C1(n39631), .C2(n32753), .A(
        n33957), .ZN(n33954) );
  OAI222_X1 U28597 ( .A1(n30967), .A2(n39625), .B1(n31031), .B2(n39619), .C1(
        n30903), .C2(n39613), .ZN(n33957) );
  AOI221_X1 U28598 ( .B1(n39385), .B2(n32801), .C1(n39379), .C2(n32753), .A(
        n35231), .ZN(n35228) );
  OAI222_X1 U28599 ( .A1(n30967), .A2(n39373), .B1(n31031), .B2(n39367), .C1(
        n30903), .C2(n39361), .ZN(n35231) );
  AOI221_X1 U28600 ( .B1(n39637), .B2(n32800), .C1(n39631), .C2(n32752), .A(
        n33976), .ZN(n33973) );
  OAI222_X1 U28601 ( .A1(n30966), .A2(n39625), .B1(n31030), .B2(n39619), .C1(
        n30902), .C2(n39613), .ZN(n33976) );
  AOI221_X1 U28602 ( .B1(n39385), .B2(n32800), .C1(n39379), .C2(n32752), .A(
        n35250), .ZN(n35247) );
  OAI222_X1 U28603 ( .A1(n30966), .A2(n39373), .B1(n31030), .B2(n39367), .C1(
        n30902), .C2(n39361), .ZN(n35250) );
  AOI221_X1 U28604 ( .B1(n39637), .B2(n32799), .C1(n39631), .C2(n32751), .A(
        n33995), .ZN(n33992) );
  OAI222_X1 U28605 ( .A1(n30965), .A2(n39625), .B1(n31029), .B2(n39619), .C1(
        n30901), .C2(n39613), .ZN(n33995) );
  AOI221_X1 U28606 ( .B1(n39385), .B2(n32799), .C1(n39379), .C2(n32751), .A(
        n35269), .ZN(n35266) );
  OAI222_X1 U28607 ( .A1(n30965), .A2(n39373), .B1(n31029), .B2(n39367), .C1(
        n30901), .C2(n39361), .ZN(n35269) );
  AOI221_X1 U28608 ( .B1(n39636), .B2(n32798), .C1(n39630), .C2(n32750), .A(
        n34014), .ZN(n34011) );
  OAI222_X1 U28609 ( .A1(n30964), .A2(n39624), .B1(n31028), .B2(n39618), .C1(
        n30900), .C2(n39612), .ZN(n34014) );
  AOI221_X1 U28610 ( .B1(n39384), .B2(n32798), .C1(n39378), .C2(n32750), .A(
        n35288), .ZN(n35285) );
  OAI222_X1 U28611 ( .A1(n30964), .A2(n39372), .B1(n31028), .B2(n39366), .C1(
        n30900), .C2(n39360), .ZN(n35288) );
  AOI221_X1 U28612 ( .B1(n39636), .B2(n32797), .C1(n39630), .C2(n32749), .A(
        n34033), .ZN(n34030) );
  OAI222_X1 U28613 ( .A1(n30963), .A2(n39624), .B1(n31027), .B2(n39618), .C1(
        n30899), .C2(n39612), .ZN(n34033) );
  AOI221_X1 U28614 ( .B1(n39384), .B2(n32797), .C1(n39378), .C2(n32749), .A(
        n35307), .ZN(n35304) );
  OAI222_X1 U28615 ( .A1(n30963), .A2(n39372), .B1(n31027), .B2(n39366), .C1(
        n30899), .C2(n39360), .ZN(n35307) );
  AOI221_X1 U28616 ( .B1(n39636), .B2(n32796), .C1(n39630), .C2(n32748), .A(
        n34052), .ZN(n34049) );
  OAI222_X1 U28617 ( .A1(n30962), .A2(n39624), .B1(n31026), .B2(n39618), .C1(
        n30898), .C2(n39612), .ZN(n34052) );
  AOI221_X1 U28618 ( .B1(n39384), .B2(n32796), .C1(n39378), .C2(n32748), .A(
        n35326), .ZN(n35323) );
  OAI222_X1 U28619 ( .A1(n30962), .A2(n39372), .B1(n31026), .B2(n39366), .C1(
        n30898), .C2(n39360), .ZN(n35326) );
  AOI221_X1 U28620 ( .B1(n39636), .B2(n32795), .C1(n39630), .C2(n32747), .A(
        n34071), .ZN(n34068) );
  OAI222_X1 U28621 ( .A1(n30961), .A2(n39624), .B1(n31025), .B2(n39618), .C1(
        n30897), .C2(n39612), .ZN(n34071) );
  AOI221_X1 U28622 ( .B1(n39384), .B2(n32795), .C1(n39378), .C2(n32747), .A(
        n35345), .ZN(n35342) );
  OAI222_X1 U28623 ( .A1(n30961), .A2(n39372), .B1(n31025), .B2(n39366), .C1(
        n30897), .C2(n39360), .ZN(n35345) );
  AOI221_X1 U28624 ( .B1(n39636), .B2(n32794), .C1(n39630), .C2(n32746), .A(
        n34090), .ZN(n34087) );
  OAI222_X1 U28625 ( .A1(n30960), .A2(n39624), .B1(n31024), .B2(n39618), .C1(
        n30896), .C2(n39612), .ZN(n34090) );
  AOI221_X1 U28626 ( .B1(n39384), .B2(n32794), .C1(n39378), .C2(n32746), .A(
        n35364), .ZN(n35361) );
  OAI222_X1 U28627 ( .A1(n30960), .A2(n39372), .B1(n31024), .B2(n39366), .C1(
        n30896), .C2(n39360), .ZN(n35364) );
  AOI221_X1 U28628 ( .B1(n39636), .B2(n32793), .C1(n39630), .C2(n32745), .A(
        n34109), .ZN(n34106) );
  OAI222_X1 U28629 ( .A1(n30959), .A2(n39624), .B1(n31023), .B2(n39618), .C1(
        n30895), .C2(n39612), .ZN(n34109) );
  AOI221_X1 U28630 ( .B1(n39384), .B2(n32793), .C1(n39378), .C2(n32745), .A(
        n35383), .ZN(n35380) );
  OAI222_X1 U28631 ( .A1(n30959), .A2(n39372), .B1(n31023), .B2(n39366), .C1(
        n30895), .C2(n39360), .ZN(n35383) );
  AOI221_X1 U28632 ( .B1(n39636), .B2(n32792), .C1(n39630), .C2(n32744), .A(
        n34128), .ZN(n34125) );
  OAI222_X1 U28633 ( .A1(n30958), .A2(n39624), .B1(n31022), .B2(n39618), .C1(
        n30894), .C2(n39612), .ZN(n34128) );
  AOI221_X1 U28634 ( .B1(n39384), .B2(n32792), .C1(n39378), .C2(n32744), .A(
        n35402), .ZN(n35399) );
  OAI222_X1 U28635 ( .A1(n30958), .A2(n39372), .B1(n31022), .B2(n39366), .C1(
        n30894), .C2(n39360), .ZN(n35402) );
  AOI221_X1 U28636 ( .B1(n39636), .B2(n32791), .C1(n39630), .C2(n32743), .A(
        n34147), .ZN(n34144) );
  OAI222_X1 U28637 ( .A1(n30957), .A2(n39624), .B1(n31021), .B2(n39618), .C1(
        n30893), .C2(n39612), .ZN(n34147) );
  AOI221_X1 U28638 ( .B1(n39384), .B2(n32791), .C1(n39378), .C2(n32743), .A(
        n35421), .ZN(n35418) );
  OAI222_X1 U28639 ( .A1(n30957), .A2(n39372), .B1(n31021), .B2(n39366), .C1(
        n30893), .C2(n39360), .ZN(n35421) );
  AOI221_X1 U28640 ( .B1(n39636), .B2(n32790), .C1(n39630), .C2(n32742), .A(
        n34166), .ZN(n34163) );
  OAI222_X1 U28641 ( .A1(n30956), .A2(n39624), .B1(n31020), .B2(n39618), .C1(
        n30892), .C2(n39612), .ZN(n34166) );
  AOI221_X1 U28642 ( .B1(n39384), .B2(n32790), .C1(n39378), .C2(n32742), .A(
        n35440), .ZN(n35437) );
  OAI222_X1 U28643 ( .A1(n30956), .A2(n39372), .B1(n31020), .B2(n39366), .C1(
        n30892), .C2(n39360), .ZN(n35440) );
  AOI221_X1 U28644 ( .B1(n39636), .B2(n32789), .C1(n39630), .C2(n32741), .A(
        n34185), .ZN(n34182) );
  OAI222_X1 U28645 ( .A1(n30955), .A2(n39624), .B1(n31019), .B2(n39618), .C1(
        n30891), .C2(n39612), .ZN(n34185) );
  AOI221_X1 U28646 ( .B1(n39384), .B2(n32789), .C1(n39378), .C2(n32741), .A(
        n35459), .ZN(n35456) );
  OAI222_X1 U28647 ( .A1(n30955), .A2(n39372), .B1(n31019), .B2(n39366), .C1(
        n30891), .C2(n39360), .ZN(n35459) );
  AOI221_X1 U28648 ( .B1(n39636), .B2(n32788), .C1(n39630), .C2(n32740), .A(
        n34204), .ZN(n34201) );
  OAI222_X1 U28649 ( .A1(n30954), .A2(n39624), .B1(n31018), .B2(n39618), .C1(
        n30890), .C2(n39612), .ZN(n34204) );
  AOI221_X1 U28650 ( .B1(n39384), .B2(n32788), .C1(n39378), .C2(n32740), .A(
        n35478), .ZN(n35475) );
  OAI222_X1 U28651 ( .A1(n30954), .A2(n39372), .B1(n31018), .B2(n39366), .C1(
        n30890), .C2(n39360), .ZN(n35478) );
  AOI221_X1 U28652 ( .B1(n39636), .B2(n32787), .C1(n39630), .C2(n32739), .A(
        n34223), .ZN(n34220) );
  OAI222_X1 U28653 ( .A1(n30953), .A2(n39624), .B1(n31017), .B2(n39618), .C1(
        n30889), .C2(n39612), .ZN(n34223) );
  AOI221_X1 U28654 ( .B1(n39384), .B2(n32787), .C1(n39378), .C2(n32739), .A(
        n35497), .ZN(n35494) );
  OAI222_X1 U28655 ( .A1(n30953), .A2(n39372), .B1(n31017), .B2(n39366), .C1(
        n30889), .C2(n39360), .ZN(n35497) );
  AOI221_X1 U28656 ( .B1(n39635), .B2(n32786), .C1(n39629), .C2(n32738), .A(
        n34242), .ZN(n34239) );
  OAI222_X1 U28657 ( .A1(n30952), .A2(n39623), .B1(n31016), .B2(n39617), .C1(
        n30888), .C2(n39611), .ZN(n34242) );
  AOI221_X1 U28658 ( .B1(n39383), .B2(n32786), .C1(n39377), .C2(n32738), .A(
        n35516), .ZN(n35513) );
  OAI222_X1 U28659 ( .A1(n30952), .A2(n39371), .B1(n31016), .B2(n39365), .C1(
        n30888), .C2(n39359), .ZN(n35516) );
  AOI221_X1 U28660 ( .B1(n39635), .B2(n32785), .C1(n39629), .C2(n32737), .A(
        n34261), .ZN(n34258) );
  OAI222_X1 U28661 ( .A1(n30951), .A2(n39623), .B1(n31015), .B2(n39617), .C1(
        n30887), .C2(n39611), .ZN(n34261) );
  AOI221_X1 U28662 ( .B1(n39383), .B2(n32785), .C1(n39377), .C2(n32737), .A(
        n35535), .ZN(n35532) );
  OAI222_X1 U28663 ( .A1(n30951), .A2(n39371), .B1(n31015), .B2(n39365), .C1(
        n30887), .C2(n39359), .ZN(n35535) );
  AOI221_X1 U28664 ( .B1(n39635), .B2(n32784), .C1(n39629), .C2(n32736), .A(
        n34280), .ZN(n34277) );
  OAI222_X1 U28665 ( .A1(n30950), .A2(n39623), .B1(n31014), .B2(n39617), .C1(
        n30886), .C2(n39611), .ZN(n34280) );
  AOI221_X1 U28666 ( .B1(n39383), .B2(n32784), .C1(n39377), .C2(n32736), .A(
        n35554), .ZN(n35551) );
  OAI222_X1 U28667 ( .A1(n30950), .A2(n39371), .B1(n31014), .B2(n39365), .C1(
        n30886), .C2(n39359), .ZN(n35554) );
  AOI221_X1 U28668 ( .B1(n39635), .B2(n32783), .C1(n39629), .C2(n32735), .A(
        n34299), .ZN(n34296) );
  OAI222_X1 U28669 ( .A1(n30949), .A2(n39623), .B1(n31013), .B2(n39617), .C1(
        n30885), .C2(n39611), .ZN(n34299) );
  AOI221_X1 U28670 ( .B1(n39383), .B2(n32783), .C1(n39377), .C2(n32735), .A(
        n35573), .ZN(n35570) );
  OAI222_X1 U28671 ( .A1(n30949), .A2(n39371), .B1(n31013), .B2(n39365), .C1(
        n30885), .C2(n39359), .ZN(n35573) );
  AOI221_X1 U28672 ( .B1(n39635), .B2(n32782), .C1(n39629), .C2(n32734), .A(
        n34318), .ZN(n34315) );
  OAI222_X1 U28673 ( .A1(n30948), .A2(n39623), .B1(n31012), .B2(n39617), .C1(
        n30884), .C2(n39611), .ZN(n34318) );
  AOI221_X1 U28674 ( .B1(n39383), .B2(n32782), .C1(n39377), .C2(n32734), .A(
        n35592), .ZN(n35589) );
  OAI222_X1 U28675 ( .A1(n30948), .A2(n39371), .B1(n31012), .B2(n39365), .C1(
        n30884), .C2(n39359), .ZN(n35592) );
  AOI221_X1 U28676 ( .B1(n39635), .B2(n32781), .C1(n39629), .C2(n32733), .A(
        n34337), .ZN(n34334) );
  OAI222_X1 U28677 ( .A1(n30947), .A2(n39623), .B1(n31011), .B2(n39617), .C1(
        n30883), .C2(n39611), .ZN(n34337) );
  AOI221_X1 U28678 ( .B1(n39383), .B2(n32781), .C1(n39377), .C2(n32733), .A(
        n35611), .ZN(n35608) );
  OAI222_X1 U28679 ( .A1(n30947), .A2(n39371), .B1(n31011), .B2(n39365), .C1(
        n30883), .C2(n39359), .ZN(n35611) );
  AOI221_X1 U28680 ( .B1(n39635), .B2(n32780), .C1(n39629), .C2(n32732), .A(
        n34356), .ZN(n34353) );
  OAI222_X1 U28681 ( .A1(n30946), .A2(n39623), .B1(n31010), .B2(n39617), .C1(
        n30882), .C2(n39611), .ZN(n34356) );
  AOI221_X1 U28682 ( .B1(n39383), .B2(n32780), .C1(n39377), .C2(n32732), .A(
        n35630), .ZN(n35627) );
  OAI222_X1 U28683 ( .A1(n30946), .A2(n39371), .B1(n31010), .B2(n39365), .C1(
        n30882), .C2(n39359), .ZN(n35630) );
  AOI221_X1 U28684 ( .B1(n39635), .B2(n32779), .C1(n39629), .C2(n32731), .A(
        n34375), .ZN(n34372) );
  OAI222_X1 U28685 ( .A1(n30945), .A2(n39623), .B1(n31009), .B2(n39617), .C1(
        n30881), .C2(n39611), .ZN(n34375) );
  AOI221_X1 U28686 ( .B1(n39383), .B2(n32779), .C1(n39377), .C2(n32731), .A(
        n35649), .ZN(n35646) );
  OAI222_X1 U28687 ( .A1(n30945), .A2(n39371), .B1(n31009), .B2(n39365), .C1(
        n30881), .C2(n39359), .ZN(n35649) );
  AOI221_X1 U28688 ( .B1(n39635), .B2(n32778), .C1(n39629), .C2(n32730), .A(
        n34394), .ZN(n34391) );
  OAI222_X1 U28689 ( .A1(n30944), .A2(n39623), .B1(n31008), .B2(n39617), .C1(
        n30880), .C2(n39611), .ZN(n34394) );
  AOI221_X1 U28690 ( .B1(n39383), .B2(n32778), .C1(n39377), .C2(n32730), .A(
        n35668), .ZN(n35665) );
  OAI222_X1 U28691 ( .A1(n30944), .A2(n39371), .B1(n31008), .B2(n39365), .C1(
        n30880), .C2(n39359), .ZN(n35668) );
  AOI221_X1 U28692 ( .B1(n39635), .B2(n32777), .C1(n39629), .C2(n32729), .A(
        n34413), .ZN(n34410) );
  OAI222_X1 U28693 ( .A1(n30943), .A2(n39623), .B1(n31007), .B2(n39617), .C1(
        n30879), .C2(n39611), .ZN(n34413) );
  AOI221_X1 U28694 ( .B1(n39383), .B2(n32777), .C1(n39377), .C2(n32729), .A(
        n35687), .ZN(n35684) );
  OAI222_X1 U28695 ( .A1(n30943), .A2(n39371), .B1(n31007), .B2(n39365), .C1(
        n30879), .C2(n39359), .ZN(n35687) );
  AOI221_X1 U28696 ( .B1(n39635), .B2(n32776), .C1(n39629), .C2(n32728), .A(
        n34432), .ZN(n34429) );
  OAI222_X1 U28697 ( .A1(n30942), .A2(n39623), .B1(n31006), .B2(n39617), .C1(
        n30878), .C2(n39611), .ZN(n34432) );
  AOI221_X1 U28698 ( .B1(n39383), .B2(n32776), .C1(n39377), .C2(n32728), .A(
        n35706), .ZN(n35703) );
  OAI222_X1 U28699 ( .A1(n30942), .A2(n39371), .B1(n31006), .B2(n39365), .C1(
        n30878), .C2(n39359), .ZN(n35706) );
  AOI221_X1 U28700 ( .B1(n39635), .B2(n32775), .C1(n39629), .C2(n32727), .A(
        n34451), .ZN(n34448) );
  OAI222_X1 U28701 ( .A1(n30941), .A2(n39623), .B1(n31005), .B2(n39617), .C1(
        n30877), .C2(n39611), .ZN(n34451) );
  AOI221_X1 U28702 ( .B1(n39383), .B2(n32775), .C1(n39377), .C2(n32727), .A(
        n35725), .ZN(n35722) );
  OAI222_X1 U28703 ( .A1(n30941), .A2(n39371), .B1(n31005), .B2(n39365), .C1(
        n30877), .C2(n39359), .ZN(n35725) );
  AOI221_X1 U28704 ( .B1(n39634), .B2(n32846), .C1(n39628), .C2(n32834), .A(
        n34470), .ZN(n34467) );
  OAI222_X1 U28705 ( .A1(n30940), .A2(n39622), .B1(n31004), .B2(n39616), .C1(
        n30876), .C2(n39610), .ZN(n34470) );
  AOI221_X1 U28706 ( .B1(n39382), .B2(n32846), .C1(n39376), .C2(n32834), .A(
        n35744), .ZN(n35741) );
  OAI222_X1 U28707 ( .A1(n30940), .A2(n39370), .B1(n31004), .B2(n39364), .C1(
        n30876), .C2(n39358), .ZN(n35744) );
  AOI221_X1 U28708 ( .B1(n39634), .B2(n32845), .C1(n39628), .C2(n32833), .A(
        n34489), .ZN(n34486) );
  OAI222_X1 U28709 ( .A1(n30939), .A2(n39622), .B1(n31003), .B2(n39616), .C1(
        n30875), .C2(n39610), .ZN(n34489) );
  AOI221_X1 U28710 ( .B1(n39382), .B2(n32845), .C1(n39376), .C2(n32833), .A(
        n35763), .ZN(n35760) );
  OAI222_X1 U28711 ( .A1(n30939), .A2(n39370), .B1(n31003), .B2(n39364), .C1(
        n30875), .C2(n39358), .ZN(n35763) );
  AOI221_X1 U28712 ( .B1(n39634), .B2(n32844), .C1(n39628), .C2(n32832), .A(
        n34508), .ZN(n34505) );
  OAI222_X1 U28713 ( .A1(n30938), .A2(n39622), .B1(n31002), .B2(n39616), .C1(
        n30874), .C2(n39610), .ZN(n34508) );
  AOI221_X1 U28714 ( .B1(n39382), .B2(n32844), .C1(n39376), .C2(n32832), .A(
        n35782), .ZN(n35779) );
  OAI222_X1 U28715 ( .A1(n30938), .A2(n39370), .B1(n31002), .B2(n39364), .C1(
        n30874), .C2(n39358), .ZN(n35782) );
  AOI221_X1 U28716 ( .B1(n39634), .B2(n32843), .C1(n39628), .C2(n32831), .A(
        n34527), .ZN(n34524) );
  OAI222_X1 U28717 ( .A1(n30937), .A2(n39622), .B1(n31001), .B2(n39616), .C1(
        n30873), .C2(n39610), .ZN(n34527) );
  AOI221_X1 U28718 ( .B1(n39382), .B2(n32843), .C1(n39376), .C2(n32831), .A(
        n35801), .ZN(n35798) );
  OAI222_X1 U28719 ( .A1(n30937), .A2(n39370), .B1(n31001), .B2(n39364), .C1(
        n30873), .C2(n39358), .ZN(n35801) );
  AOI221_X1 U28720 ( .B1(n39634), .B2(n32842), .C1(n39628), .C2(n32830), .A(
        n34546), .ZN(n34543) );
  OAI222_X1 U28721 ( .A1(n30936), .A2(n39622), .B1(n31000), .B2(n39616), .C1(
        n30872), .C2(n39610), .ZN(n34546) );
  AOI221_X1 U28722 ( .B1(n39382), .B2(n32842), .C1(n39376), .C2(n32830), .A(
        n35820), .ZN(n35817) );
  OAI222_X1 U28723 ( .A1(n30936), .A2(n39370), .B1(n31000), .B2(n39364), .C1(
        n30872), .C2(n39358), .ZN(n35820) );
  AOI221_X1 U28724 ( .B1(n39634), .B2(n32841), .C1(n39628), .C2(n32829), .A(
        n34565), .ZN(n34562) );
  OAI222_X1 U28725 ( .A1(n30935), .A2(n39622), .B1(n30999), .B2(n39616), .C1(
        n30871), .C2(n39610), .ZN(n34565) );
  AOI221_X1 U28726 ( .B1(n39382), .B2(n32841), .C1(n39376), .C2(n32829), .A(
        n35839), .ZN(n35836) );
  OAI222_X1 U28727 ( .A1(n30935), .A2(n39370), .B1(n30999), .B2(n39364), .C1(
        n30871), .C2(n39358), .ZN(n35839) );
  AOI221_X1 U28728 ( .B1(n39634), .B2(n32840), .C1(n39628), .C2(n32828), .A(
        n34584), .ZN(n34581) );
  OAI222_X1 U28729 ( .A1(n30934), .A2(n39622), .B1(n30998), .B2(n39616), .C1(
        n30870), .C2(n39610), .ZN(n34584) );
  AOI221_X1 U28730 ( .B1(n39382), .B2(n32840), .C1(n39376), .C2(n32828), .A(
        n35858), .ZN(n35855) );
  OAI222_X1 U28731 ( .A1(n30934), .A2(n39370), .B1(n30998), .B2(n39364), .C1(
        n30870), .C2(n39358), .ZN(n35858) );
  AOI221_X1 U28732 ( .B1(n39634), .B2(n32839), .C1(n39628), .C2(n32827), .A(
        n34603), .ZN(n34600) );
  OAI222_X1 U28733 ( .A1(n30933), .A2(n39622), .B1(n30997), .B2(n39616), .C1(
        n30869), .C2(n39610), .ZN(n34603) );
  AOI221_X1 U28734 ( .B1(n39382), .B2(n32839), .C1(n39376), .C2(n32827), .A(
        n35877), .ZN(n35874) );
  OAI222_X1 U28735 ( .A1(n30933), .A2(n39370), .B1(n30997), .B2(n39364), .C1(
        n30869), .C2(n39358), .ZN(n35877) );
  AOI221_X1 U28736 ( .B1(n39634), .B2(n32838), .C1(n39628), .C2(n32826), .A(
        n34622), .ZN(n34619) );
  OAI222_X1 U28737 ( .A1(n30932), .A2(n39622), .B1(n30996), .B2(n39616), .C1(
        n30868), .C2(n39610), .ZN(n34622) );
  AOI221_X1 U28738 ( .B1(n39382), .B2(n32838), .C1(n39376), .C2(n32826), .A(
        n35896), .ZN(n35893) );
  OAI222_X1 U28739 ( .A1(n30932), .A2(n39370), .B1(n30996), .B2(n39364), .C1(
        n30868), .C2(n39358), .ZN(n35896) );
  AOI221_X1 U28740 ( .B1(n39634), .B2(n32837), .C1(n39628), .C2(n32825), .A(
        n34641), .ZN(n34638) );
  OAI222_X1 U28741 ( .A1(n30931), .A2(n39622), .B1(n30995), .B2(n39616), .C1(
        n30867), .C2(n39610), .ZN(n34641) );
  AOI221_X1 U28742 ( .B1(n39382), .B2(n32837), .C1(n39376), .C2(n32825), .A(
        n35915), .ZN(n35912) );
  OAI222_X1 U28743 ( .A1(n30931), .A2(n39370), .B1(n30995), .B2(n39364), .C1(
        n30867), .C2(n39358), .ZN(n35915) );
  AOI221_X1 U28744 ( .B1(n39634), .B2(n32836), .C1(n39628), .C2(n32824), .A(
        n34660), .ZN(n34657) );
  OAI222_X1 U28745 ( .A1(n30930), .A2(n39622), .B1(n30994), .B2(n39616), .C1(
        n30866), .C2(n39610), .ZN(n34660) );
  AOI221_X1 U28746 ( .B1(n39382), .B2(n32836), .C1(n39376), .C2(n32824), .A(
        n35934), .ZN(n35931) );
  OAI222_X1 U28747 ( .A1(n30930), .A2(n39370), .B1(n30994), .B2(n39364), .C1(
        n30866), .C2(n39358), .ZN(n35934) );
  AOI221_X1 U28748 ( .B1(n39634), .B2(n32835), .C1(n39628), .C2(n32823), .A(
        n34691), .ZN(n34687) );
  OAI222_X1 U28749 ( .A1(n30929), .A2(n39622), .B1(n30993), .B2(n39616), .C1(
        n30865), .C2(n39610), .ZN(n34691) );
  AOI221_X1 U28750 ( .B1(n39382), .B2(n32835), .C1(n39376), .C2(n32823), .A(
        n35965), .ZN(n35961) );
  OAI222_X1 U28751 ( .A1(n30929), .A2(n39370), .B1(n30993), .B2(n39364), .C1(
        n30865), .C2(n39358), .ZN(n35965) );
  NOR2_X1 U28752 ( .A1(N932), .A2(N931), .ZN(n33294) );
  OAI222_X1 U28753 ( .A1(n40952), .A2(n39895), .B1(n41336), .B2(n39888), .C1(
        n39886), .C2(n30613), .ZN(n7591) );
  OAI222_X1 U28754 ( .A1(n40964), .A2(n39895), .B1(n41348), .B2(n39888), .C1(
        n39886), .C2(n30611), .ZN(n7589) );
  OAI222_X1 U28755 ( .A1(n40970), .A2(n39895), .B1(n41354), .B2(n39888), .C1(
        n39886), .C2(n30610), .ZN(n7588) );
  OAI222_X1 U28756 ( .A1(n40976), .A2(n39895), .B1(n41360), .B2(n39888), .C1(
        n39886), .C2(n30609), .ZN(n7587) );
  OAI222_X1 U28757 ( .A1(n40954), .A2(n40390), .B1(n41338), .B2(n40383), .C1(
        n40381), .C2(n31691), .ZN(n9191) );
  OAI222_X1 U28758 ( .A1(n40966), .A2(n40390), .B1(n41350), .B2(n40383), .C1(
        n40381), .C2(n31689), .ZN(n9189) );
  OAI222_X1 U28759 ( .A1(n40972), .A2(n40390), .B1(n41356), .B2(n40383), .C1(
        n40381), .C2(n31688), .ZN(n9188) );
  OAI222_X1 U28760 ( .A1(n40978), .A2(n40390), .B1(n41362), .B2(n40383), .C1(
        n40381), .C2(n31687), .ZN(n9187) );
  OAI222_X1 U28761 ( .A1(n40954), .A2(n40370), .B1(n41338), .B2(n40363), .C1(
        n40361), .C2(n31627), .ZN(n9127) );
  OAI222_X1 U28762 ( .A1(n40966), .A2(n40370), .B1(n41350), .B2(n40363), .C1(
        n40361), .C2(n31625), .ZN(n9125) );
  OAI222_X1 U28763 ( .A1(n40972), .A2(n40370), .B1(n41356), .B2(n40363), .C1(
        n40361), .C2(n31624), .ZN(n9124) );
  OAI222_X1 U28764 ( .A1(n40978), .A2(n40370), .B1(n41362), .B2(n40363), .C1(
        n40361), .C2(n31623), .ZN(n9123) );
  OAI222_X1 U28765 ( .A1(n40954), .A2(n40350), .B1(n41338), .B2(n40343), .C1(
        n40341), .C2(n31563), .ZN(n9063) );
  OAI222_X1 U28766 ( .A1(n40966), .A2(n40350), .B1(n41350), .B2(n40343), .C1(
        n40341), .C2(n31561), .ZN(n9061) );
  OAI222_X1 U28767 ( .A1(n40972), .A2(n40350), .B1(n41356), .B2(n40343), .C1(
        n40341), .C2(n31560), .ZN(n9060) );
  OAI222_X1 U28768 ( .A1(n40978), .A2(n40350), .B1(n41362), .B2(n40343), .C1(
        n40341), .C2(n31559), .ZN(n9059) );
  OAI222_X1 U28769 ( .A1(n40954), .A2(n40290), .B1(n41338), .B2(n40283), .C1(
        n40281), .C2(n31499), .ZN(n8871) );
  OAI222_X1 U28770 ( .A1(n40966), .A2(n40290), .B1(n41350), .B2(n40283), .C1(
        n40281), .C2(n31497), .ZN(n8869) );
  OAI222_X1 U28771 ( .A1(n40972), .A2(n40290), .B1(n41356), .B2(n40283), .C1(
        n40281), .C2(n31496), .ZN(n8868) );
  OAI222_X1 U28772 ( .A1(n40978), .A2(n40290), .B1(n41362), .B2(n40283), .C1(
        n40281), .C2(n31495), .ZN(n8867) );
  OAI222_X1 U28773 ( .A1(n40953), .A2(n40270), .B1(n41337), .B2(n40263), .C1(
        n40261), .C2(n31435), .ZN(n8807) );
  OAI222_X1 U28774 ( .A1(n40965), .A2(n40270), .B1(n41349), .B2(n40263), .C1(
        n40261), .C2(n31433), .ZN(n8805) );
  OAI222_X1 U28775 ( .A1(n40971), .A2(n40270), .B1(n41355), .B2(n40263), .C1(
        n40261), .C2(n31432), .ZN(n8804) );
  OAI222_X1 U28776 ( .A1(n40977), .A2(n40270), .B1(n41361), .B2(n40263), .C1(
        n40261), .C2(n31431), .ZN(n8803) );
  OAI222_X1 U28777 ( .A1(n40953), .A2(n40250), .B1(n41337), .B2(n40243), .C1(
        n40241), .C2(n31371), .ZN(n8743) );
  OAI222_X1 U28778 ( .A1(n40965), .A2(n40250), .B1(n41349), .B2(n40243), .C1(
        n40241), .C2(n31369), .ZN(n8741) );
  OAI222_X1 U28779 ( .A1(n40971), .A2(n40250), .B1(n41355), .B2(n40243), .C1(
        n40241), .C2(n31368), .ZN(n8740) );
  OAI222_X1 U28780 ( .A1(n40977), .A2(n40250), .B1(n41361), .B2(n40243), .C1(
        n40241), .C2(n31367), .ZN(n8739) );
  OAI222_X1 U28781 ( .A1(n40953), .A2(n40190), .B1(n41337), .B2(n40183), .C1(
        n40181), .C2(n31307), .ZN(n8551) );
  OAI222_X1 U28782 ( .A1(n40965), .A2(n40190), .B1(n41349), .B2(n40183), .C1(
        n40181), .C2(n31305), .ZN(n8549) );
  OAI222_X1 U28783 ( .A1(n40971), .A2(n40190), .B1(n41355), .B2(n40183), .C1(
        n40181), .C2(n31304), .ZN(n8548) );
  OAI222_X1 U28784 ( .A1(n40977), .A2(n40190), .B1(n41361), .B2(n40183), .C1(
        n40181), .C2(n31303), .ZN(n8547) );
  OAI222_X1 U28785 ( .A1(n40953), .A2(n40170), .B1(n41337), .B2(n40163), .C1(
        n40161), .C2(n31243), .ZN(n8487) );
  OAI222_X1 U28786 ( .A1(n40965), .A2(n40170), .B1(n41349), .B2(n40163), .C1(
        n40161), .C2(n31241), .ZN(n8485) );
  OAI222_X1 U28787 ( .A1(n40971), .A2(n40170), .B1(n41355), .B2(n40163), .C1(
        n40161), .C2(n31240), .ZN(n8484) );
  OAI222_X1 U28788 ( .A1(n40977), .A2(n40170), .B1(n41361), .B2(n40163), .C1(
        n40161), .C2(n31239), .ZN(n8483) );
  OAI222_X1 U28789 ( .A1(n40953), .A2(n40150), .B1(n41337), .B2(n40143), .C1(
        n40141), .C2(n31179), .ZN(n8423) );
  OAI222_X1 U28790 ( .A1(n40965), .A2(n40150), .B1(n41349), .B2(n40143), .C1(
        n40141), .C2(n31177), .ZN(n8421) );
  OAI222_X1 U28791 ( .A1(n40971), .A2(n40150), .B1(n41355), .B2(n40143), .C1(
        n40141), .C2(n31176), .ZN(n8420) );
  OAI222_X1 U28792 ( .A1(n40977), .A2(n40150), .B1(n41361), .B2(n40143), .C1(
        n40141), .C2(n31175), .ZN(n8419) );
  OAI222_X1 U28793 ( .A1(n40953), .A2(n40091), .B1(n41337), .B2(n40084), .C1(
        n40082), .C2(n30997), .ZN(n8231) );
  OAI222_X1 U28794 ( .A1(n40965), .A2(n40091), .B1(n41349), .B2(n40084), .C1(
        n40082), .C2(n30995), .ZN(n8229) );
  OAI222_X1 U28795 ( .A1(n40971), .A2(n40091), .B1(n41355), .B2(n40084), .C1(
        n40082), .C2(n30994), .ZN(n8228) );
  OAI222_X1 U28796 ( .A1(n40977), .A2(n40091), .B1(n41361), .B2(n40084), .C1(
        n40082), .C2(n30993), .ZN(n8227) );
  OAI222_X1 U28797 ( .A1(n40953), .A2(n40071), .B1(n41337), .B2(n40064), .C1(
        n40062), .C2(n30933), .ZN(n8167) );
  OAI222_X1 U28798 ( .A1(n40965), .A2(n40071), .B1(n41349), .B2(n40064), .C1(
        n40062), .C2(n30931), .ZN(n8165) );
  OAI222_X1 U28799 ( .A1(n40971), .A2(n40071), .B1(n41355), .B2(n40064), .C1(
        n40062), .C2(n30930), .ZN(n8164) );
  OAI222_X1 U28800 ( .A1(n40977), .A2(n40071), .B1(n41361), .B2(n40064), .C1(
        n40062), .C2(n30929), .ZN(n8163) );
  OAI222_X1 U28801 ( .A1(n40953), .A2(n40051), .B1(n41337), .B2(n40044), .C1(
        n40042), .C2(n30869), .ZN(n8103) );
  OAI222_X1 U28802 ( .A1(n40965), .A2(n40051), .B1(n41349), .B2(n40044), .C1(
        n40042), .C2(n30867), .ZN(n8101) );
  OAI222_X1 U28803 ( .A1(n40971), .A2(n40051), .B1(n41355), .B2(n40044), .C1(
        n40042), .C2(n30866), .ZN(n8100) );
  OAI222_X1 U28804 ( .A1(n40977), .A2(n40051), .B1(n41361), .B2(n40044), .C1(
        n40042), .C2(n30865), .ZN(n8099) );
  OAI222_X1 U28805 ( .A1(n40952), .A2(n39993), .B1(n41336), .B2(n39986), .C1(
        n39984), .C2(n30805), .ZN(n7911) );
  OAI222_X1 U28806 ( .A1(n40964), .A2(n39993), .B1(n41348), .B2(n39986), .C1(
        n39984), .C2(n30803), .ZN(n7909) );
  OAI222_X1 U28807 ( .A1(n40970), .A2(n39993), .B1(n41354), .B2(n39986), .C1(
        n39984), .C2(n30802), .ZN(n7908) );
  OAI222_X1 U28808 ( .A1(n40976), .A2(n39993), .B1(n41360), .B2(n39986), .C1(
        n39984), .C2(n30801), .ZN(n7907) );
  OAI222_X1 U28809 ( .A1(n40952), .A2(n39973), .B1(n41336), .B2(n39966), .C1(
        n39964), .C2(n30741), .ZN(n7847) );
  OAI222_X1 U28810 ( .A1(n40964), .A2(n39973), .B1(n41348), .B2(n39966), .C1(
        n39964), .C2(n30739), .ZN(n7845) );
  OAI222_X1 U28811 ( .A1(n40970), .A2(n39973), .B1(n41354), .B2(n39966), .C1(
        n39964), .C2(n30738), .ZN(n7844) );
  OAI222_X1 U28812 ( .A1(n40976), .A2(n39973), .B1(n41360), .B2(n39966), .C1(
        n39964), .C2(n30737), .ZN(n7843) );
  OAI222_X1 U28813 ( .A1(n40590), .A2(n40955), .B1(n40583), .B2(n41339), .C1(
        n40581), .C2(n32054), .ZN(n9831) );
  OAI222_X1 U28814 ( .A1(n40590), .A2(n40967), .B1(n40583), .B2(n41351), .C1(
        n40581), .C2(n32053), .ZN(n9829) );
  OAI222_X1 U28815 ( .A1(n40590), .A2(n40973), .B1(n40583), .B2(n41357), .C1(
        n40581), .C2(n32052), .ZN(n9828) );
  OAI222_X1 U28816 ( .A1(n40590), .A2(n40979), .B1(n40583), .B2(n41363), .C1(
        n40581), .C2(n32051), .ZN(n9827) );
  OAI222_X1 U28817 ( .A1(n40955), .A2(n40570), .B1(n41339), .B2(n40563), .C1(
        n40561), .C2(n31995), .ZN(n9767) );
  OAI222_X1 U28818 ( .A1(n40967), .A2(n40570), .B1(n41351), .B2(n40563), .C1(
        n40561), .C2(n31993), .ZN(n9765) );
  OAI222_X1 U28819 ( .A1(n40973), .A2(n40570), .B1(n41357), .B2(n40563), .C1(
        n40561), .C2(n31992), .ZN(n9764) );
  OAI222_X1 U28820 ( .A1(n40979), .A2(n40570), .B1(n41363), .B2(n40563), .C1(
        n40561), .C2(n31991), .ZN(n9763) );
  OAI222_X1 U28821 ( .A1(n40955), .A2(n40550), .B1(n41339), .B2(n40543), .C1(
        n40541), .C2(n31935), .ZN(n9703) );
  OAI222_X1 U28822 ( .A1(n40967), .A2(n40550), .B1(n41351), .B2(n40543), .C1(
        n40541), .C2(n31933), .ZN(n9701) );
  OAI222_X1 U28823 ( .A1(n40973), .A2(n40550), .B1(n41357), .B2(n40543), .C1(
        n40541), .C2(n31932), .ZN(n9700) );
  OAI222_X1 U28824 ( .A1(n40979), .A2(n40550), .B1(n41363), .B2(n40543), .C1(
        n40541), .C2(n31931), .ZN(n9699) );
  OAI222_X1 U28825 ( .A1(n40954), .A2(n40490), .B1(n41338), .B2(n40483), .C1(
        n40481), .C2(n31875), .ZN(n9511) );
  OAI222_X1 U28826 ( .A1(n40966), .A2(n40490), .B1(n41350), .B2(n40483), .C1(
        n40481), .C2(n31873), .ZN(n9509) );
  OAI222_X1 U28827 ( .A1(n40972), .A2(n40490), .B1(n41356), .B2(n40483), .C1(
        n40481), .C2(n31872), .ZN(n9508) );
  OAI222_X1 U28828 ( .A1(n40978), .A2(n40490), .B1(n41362), .B2(n40483), .C1(
        n40481), .C2(n31871), .ZN(n9507) );
  OAI222_X1 U28829 ( .A1(n40954), .A2(n40470), .B1(n41338), .B2(n40463), .C1(
        n40461), .C2(n31815), .ZN(n9447) );
  OAI222_X1 U28830 ( .A1(n40966), .A2(n40470), .B1(n41350), .B2(n40463), .C1(
        n40461), .C2(n31813), .ZN(n9445) );
  OAI222_X1 U28831 ( .A1(n40972), .A2(n40470), .B1(n41356), .B2(n40463), .C1(
        n40461), .C2(n31812), .ZN(n9444) );
  OAI222_X1 U28832 ( .A1(n40978), .A2(n40470), .B1(n41362), .B2(n40463), .C1(
        n40461), .C2(n31811), .ZN(n9443) );
  OAI222_X1 U28833 ( .A1(n40954), .A2(n40450), .B1(n41338), .B2(n40443), .C1(
        n40441), .C2(n31755), .ZN(n9383) );
  OAI222_X1 U28834 ( .A1(n40966), .A2(n40450), .B1(n41350), .B2(n40443), .C1(
        n40441), .C2(n31753), .ZN(n9381) );
  OAI222_X1 U28835 ( .A1(n40972), .A2(n40450), .B1(n41356), .B2(n40443), .C1(
        n40441), .C2(n31752), .ZN(n9380) );
  OAI222_X1 U28836 ( .A1(n40978), .A2(n40450), .B1(n41362), .B2(n40443), .C1(
        n40441), .C2(n31751), .ZN(n9379) );
  OAI222_X1 U28837 ( .A1(n40952), .A2(n39953), .B1(n41336), .B2(n39946), .C1(
        n39944), .C2(n30677), .ZN(n7783) );
  OAI222_X1 U28838 ( .A1(n40964), .A2(n39953), .B1(n41348), .B2(n39946), .C1(
        n39944), .C2(n30675), .ZN(n7781) );
  OAI222_X1 U28839 ( .A1(n40970), .A2(n39953), .B1(n41354), .B2(n39946), .C1(
        n39944), .C2(n30674), .ZN(n7780) );
  OAI222_X1 U28840 ( .A1(n40976), .A2(n39953), .B1(n41360), .B2(n39946), .C1(
        n39944), .C2(n30673), .ZN(n7779) );
  OAI222_X1 U28841 ( .A1(n40952), .A2(n39875), .B1(n41336), .B2(n39868), .C1(
        n39866), .C2(n30549), .ZN(n7527) );
  OAI222_X1 U28842 ( .A1(n40964), .A2(n39875), .B1(n41348), .B2(n39868), .C1(
        n39866), .C2(n30547), .ZN(n7525) );
  OAI222_X1 U28843 ( .A1(n40970), .A2(n39875), .B1(n41354), .B2(n39868), .C1(
        n39866), .C2(n30546), .ZN(n7524) );
  OAI222_X1 U28844 ( .A1(n40976), .A2(n39875), .B1(n41360), .B2(n39868), .C1(
        n39866), .C2(n30545), .ZN(n7523) );
  OAI222_X1 U28845 ( .A1(n40952), .A2(n39855), .B1(n41336), .B2(n39848), .C1(
        n39846), .C2(n30485), .ZN(n7463) );
  OAI222_X1 U28846 ( .A1(n40964), .A2(n39855), .B1(n41348), .B2(n39848), .C1(
        n39846), .C2(n30483), .ZN(n7461) );
  OAI222_X1 U28847 ( .A1(n40970), .A2(n39855), .B1(n41354), .B2(n39848), .C1(
        n39846), .C2(n30482), .ZN(n7460) );
  OAI222_X1 U28848 ( .A1(n40976), .A2(n39855), .B1(n41360), .B2(n39848), .C1(
        n39846), .C2(n30481), .ZN(n7459) );
  AOI221_X1 U28849 ( .B1(n39162), .B2(n31109), .C1(n39156), .C2(n31173), .A(
        n37024), .ZN(n37023) );
  OAI222_X1 U28850 ( .A1(n31291), .A2(n39150), .B1(n31355), .B2(n39144), .C1(
        n31227), .C2(n39138), .ZN(n37024) );
  AOI221_X1 U28851 ( .B1(n39163), .B2(n31108), .C1(n39157), .C2(n31172), .A(
        n37005), .ZN(n37004) );
  OAI222_X1 U28852 ( .A1(n31290), .A2(n39151), .B1(n31354), .B2(n39145), .C1(
        n31226), .C2(n39139), .ZN(n37005) );
  AOI221_X1 U28853 ( .B1(n39163), .B2(n31107), .C1(n39157), .C2(n31171), .A(
        n36986), .ZN(n36985) );
  OAI222_X1 U28854 ( .A1(n31289), .A2(n39151), .B1(n31353), .B2(n39145), .C1(
        n31225), .C2(n39139), .ZN(n36986) );
  AOI221_X1 U28855 ( .B1(n39163), .B2(n31106), .C1(n39157), .C2(n31170), .A(
        n36967), .ZN(n36966) );
  OAI222_X1 U28856 ( .A1(n31288), .A2(n39151), .B1(n31352), .B2(n39145), .C1(
        n31224), .C2(n39139), .ZN(n36967) );
  AOI221_X1 U28857 ( .B1(n39163), .B2(n31105), .C1(n39157), .C2(n31169), .A(
        n36948), .ZN(n36947) );
  OAI222_X1 U28858 ( .A1(n31287), .A2(n39151), .B1(n31351), .B2(n39145), .C1(
        n31223), .C2(n39139), .ZN(n36948) );
  AOI221_X1 U28859 ( .B1(n39163), .B2(n31104), .C1(n39157), .C2(n31168), .A(
        n36929), .ZN(n36928) );
  OAI222_X1 U28860 ( .A1(n31286), .A2(n39151), .B1(n31350), .B2(n39145), .C1(
        n31222), .C2(n39139), .ZN(n36929) );
  AOI221_X1 U28861 ( .B1(n39163), .B2(n31103), .C1(n39157), .C2(n31167), .A(
        n36910), .ZN(n36909) );
  OAI222_X1 U28862 ( .A1(n31285), .A2(n39151), .B1(n31349), .B2(n39145), .C1(
        n31221), .C2(n39139), .ZN(n36910) );
  AOI221_X1 U28863 ( .B1(n39163), .B2(n31102), .C1(n39157), .C2(n31166), .A(
        n36891), .ZN(n36890) );
  OAI222_X1 U28864 ( .A1(n31284), .A2(n39151), .B1(n31348), .B2(n39145), .C1(
        n31220), .C2(n39139), .ZN(n36891) );
  AOI221_X1 U28865 ( .B1(n39163), .B2(n31101), .C1(n39157), .C2(n31165), .A(
        n36872), .ZN(n36871) );
  OAI222_X1 U28866 ( .A1(n31283), .A2(n39151), .B1(n31347), .B2(n39145), .C1(
        n31219), .C2(n39139), .ZN(n36872) );
  AOI221_X1 U28867 ( .B1(n39163), .B2(n31100), .C1(n39157), .C2(n31164), .A(
        n36853), .ZN(n36852) );
  OAI222_X1 U28868 ( .A1(n31282), .A2(n39151), .B1(n31346), .B2(n39145), .C1(
        n31218), .C2(n39139), .ZN(n36853) );
  AOI221_X1 U28869 ( .B1(n39163), .B2(n31099), .C1(n39157), .C2(n31163), .A(
        n36834), .ZN(n36833) );
  OAI222_X1 U28870 ( .A1(n31281), .A2(n39151), .B1(n31345), .B2(n39145), .C1(
        n31217), .C2(n39139), .ZN(n36834) );
  AOI221_X1 U28871 ( .B1(n39163), .B2(n31098), .C1(n39157), .C2(n31162), .A(
        n36815), .ZN(n36814) );
  OAI222_X1 U28872 ( .A1(n31280), .A2(n39151), .B1(n31344), .B2(n39145), .C1(
        n31216), .C2(n39139), .ZN(n36815) );
  AOI221_X1 U28873 ( .B1(n39163), .B2(n31097), .C1(n39157), .C2(n31161), .A(
        n36796), .ZN(n36795) );
  OAI222_X1 U28874 ( .A1(n31279), .A2(n39151), .B1(n31343), .B2(n39145), .C1(
        n31215), .C2(n39139), .ZN(n36796) );
  AOI221_X1 U28875 ( .B1(n39164), .B2(n31096), .C1(n39158), .C2(n31160), .A(
        n36777), .ZN(n36776) );
  OAI222_X1 U28876 ( .A1(n31278), .A2(n39152), .B1(n31342), .B2(n39146), .C1(
        n31214), .C2(n39140), .ZN(n36777) );
  AOI221_X1 U28877 ( .B1(n39164), .B2(n31095), .C1(n39158), .C2(n31159), .A(
        n36758), .ZN(n36757) );
  OAI222_X1 U28878 ( .A1(n31277), .A2(n39152), .B1(n31341), .B2(n39146), .C1(
        n31213), .C2(n39140), .ZN(n36758) );
  AOI221_X1 U28879 ( .B1(n39164), .B2(n31094), .C1(n39158), .C2(n31158), .A(
        n36739), .ZN(n36738) );
  OAI222_X1 U28880 ( .A1(n31276), .A2(n39152), .B1(n31340), .B2(n39146), .C1(
        n31212), .C2(n39140), .ZN(n36739) );
  AOI221_X1 U28881 ( .B1(n39164), .B2(n31093), .C1(n39158), .C2(n31157), .A(
        n36720), .ZN(n36719) );
  OAI222_X1 U28882 ( .A1(n31275), .A2(n39152), .B1(n31339), .B2(n39146), .C1(
        n31211), .C2(n39140), .ZN(n36720) );
  AOI221_X1 U28883 ( .B1(n39164), .B2(n31092), .C1(n39158), .C2(n31156), .A(
        n36701), .ZN(n36700) );
  OAI222_X1 U28884 ( .A1(n31274), .A2(n39152), .B1(n31338), .B2(n39146), .C1(
        n31210), .C2(n39140), .ZN(n36701) );
  AOI221_X1 U28885 ( .B1(n39164), .B2(n31091), .C1(n39158), .C2(n31155), .A(
        n36682), .ZN(n36681) );
  OAI222_X1 U28886 ( .A1(n31273), .A2(n39152), .B1(n31337), .B2(n39146), .C1(
        n31209), .C2(n39140), .ZN(n36682) );
  AOI221_X1 U28887 ( .B1(n39164), .B2(n31090), .C1(n39158), .C2(n31154), .A(
        n36663), .ZN(n36662) );
  OAI222_X1 U28888 ( .A1(n31272), .A2(n39152), .B1(n31336), .B2(n39146), .C1(
        n31208), .C2(n39140), .ZN(n36663) );
  AOI221_X1 U28889 ( .B1(n39164), .B2(n31089), .C1(n39158), .C2(n31153), .A(
        n36644), .ZN(n36643) );
  OAI222_X1 U28890 ( .A1(n31271), .A2(n39152), .B1(n31335), .B2(n39146), .C1(
        n31207), .C2(n39140), .ZN(n36644) );
  AOI221_X1 U28891 ( .B1(n39164), .B2(n31088), .C1(n39158), .C2(n31152), .A(
        n36625), .ZN(n36624) );
  OAI222_X1 U28892 ( .A1(n31270), .A2(n39152), .B1(n31334), .B2(n39146), .C1(
        n31206), .C2(n39140), .ZN(n36625) );
  AOI221_X1 U28893 ( .B1(n39164), .B2(n31087), .C1(n39158), .C2(n31151), .A(
        n36606), .ZN(n36605) );
  OAI222_X1 U28894 ( .A1(n31269), .A2(n39152), .B1(n31333), .B2(n39146), .C1(
        n31205), .C2(n39140), .ZN(n36606) );
  AOI221_X1 U28895 ( .B1(n39164), .B2(n31086), .C1(n39158), .C2(n31150), .A(
        n36587), .ZN(n36586) );
  OAI222_X1 U28896 ( .A1(n31268), .A2(n39152), .B1(n31332), .B2(n39146), .C1(
        n31204), .C2(n39140), .ZN(n36587) );
  AOI221_X1 U28897 ( .B1(n39164), .B2(n31085), .C1(n39158), .C2(n31149), .A(
        n36568), .ZN(n36567) );
  OAI222_X1 U28898 ( .A1(n31267), .A2(n39152), .B1(n31331), .B2(n39146), .C1(
        n31203), .C2(n39140), .ZN(n36568) );
  AOI221_X1 U28899 ( .B1(n39165), .B2(n31084), .C1(n39159), .C2(n31148), .A(
        n36549), .ZN(n36548) );
  OAI222_X1 U28900 ( .A1(n31266), .A2(n39153), .B1(n31330), .B2(n39147), .C1(
        n31202), .C2(n39141), .ZN(n36549) );
  AOI221_X1 U28901 ( .B1(n39165), .B2(n31083), .C1(n39159), .C2(n31147), .A(
        n36530), .ZN(n36529) );
  OAI222_X1 U28902 ( .A1(n31265), .A2(n39153), .B1(n31329), .B2(n39147), .C1(
        n31201), .C2(n39141), .ZN(n36530) );
  AOI221_X1 U28903 ( .B1(n39165), .B2(n31082), .C1(n39159), .C2(n31146), .A(
        n36511), .ZN(n36510) );
  OAI222_X1 U28904 ( .A1(n31264), .A2(n39153), .B1(n31328), .B2(n39147), .C1(
        n31200), .C2(n39141), .ZN(n36511) );
  AOI221_X1 U28905 ( .B1(n39165), .B2(n31081), .C1(n39159), .C2(n31145), .A(
        n36492), .ZN(n36491) );
  OAI222_X1 U28906 ( .A1(n31263), .A2(n39153), .B1(n31327), .B2(n39147), .C1(
        n31199), .C2(n39141), .ZN(n36492) );
  AOI221_X1 U28907 ( .B1(n39165), .B2(n31080), .C1(n39159), .C2(n31144), .A(
        n36473), .ZN(n36472) );
  OAI222_X1 U28908 ( .A1(n31262), .A2(n39153), .B1(n31326), .B2(n39147), .C1(
        n31198), .C2(n39141), .ZN(n36473) );
  AOI221_X1 U28909 ( .B1(n39165), .B2(n31079), .C1(n39159), .C2(n31143), .A(
        n36454), .ZN(n36453) );
  OAI222_X1 U28910 ( .A1(n31261), .A2(n39153), .B1(n31325), .B2(n39147), .C1(
        n31197), .C2(n39141), .ZN(n36454) );
  AOI221_X1 U28911 ( .B1(n39165), .B2(n31078), .C1(n39159), .C2(n31142), .A(
        n36435), .ZN(n36434) );
  OAI222_X1 U28912 ( .A1(n31260), .A2(n39153), .B1(n31324), .B2(n39147), .C1(
        n31196), .C2(n39141), .ZN(n36435) );
  AOI221_X1 U28913 ( .B1(n39165), .B2(n31077), .C1(n39159), .C2(n31141), .A(
        n36416), .ZN(n36415) );
  OAI222_X1 U28914 ( .A1(n31259), .A2(n39153), .B1(n31323), .B2(n39147), .C1(
        n31195), .C2(n39141), .ZN(n36416) );
  AOI221_X1 U28915 ( .B1(n39165), .B2(n31076), .C1(n39159), .C2(n31140), .A(
        n36397), .ZN(n36396) );
  OAI222_X1 U28916 ( .A1(n31258), .A2(n39153), .B1(n31322), .B2(n39147), .C1(
        n31194), .C2(n39141), .ZN(n36397) );
  AOI221_X1 U28917 ( .B1(n39165), .B2(n31075), .C1(n39159), .C2(n31139), .A(
        n36378), .ZN(n36377) );
  OAI222_X1 U28918 ( .A1(n31257), .A2(n39153), .B1(n31321), .B2(n39147), .C1(
        n31193), .C2(n39141), .ZN(n36378) );
  AOI221_X1 U28919 ( .B1(n39165), .B2(n31074), .C1(n39159), .C2(n31138), .A(
        n36359), .ZN(n36358) );
  OAI222_X1 U28920 ( .A1(n31256), .A2(n39153), .B1(n31320), .B2(n39147), .C1(
        n31192), .C2(n39141), .ZN(n36359) );
  AOI221_X1 U28921 ( .B1(n39165), .B2(n31073), .C1(n39159), .C2(n31137), .A(
        n36340), .ZN(n36339) );
  OAI222_X1 U28922 ( .A1(n31255), .A2(n39153), .B1(n31319), .B2(n39147), .C1(
        n31191), .C2(n39141), .ZN(n36340) );
  AOI221_X1 U28923 ( .B1(n39166), .B2(n31072), .C1(n39160), .C2(n31136), .A(
        n36321), .ZN(n36320) );
  OAI222_X1 U28924 ( .A1(n31254), .A2(n39154), .B1(n31318), .B2(n39148), .C1(
        n31190), .C2(n39142), .ZN(n36321) );
  AOI221_X1 U28925 ( .B1(n39166), .B2(n31071), .C1(n39160), .C2(n31135), .A(
        n36302), .ZN(n36301) );
  OAI222_X1 U28926 ( .A1(n31253), .A2(n39154), .B1(n31317), .B2(n39148), .C1(
        n31189), .C2(n39142), .ZN(n36302) );
  AOI221_X1 U28927 ( .B1(n39166), .B2(n31070), .C1(n39160), .C2(n31134), .A(
        n36283), .ZN(n36282) );
  OAI222_X1 U28928 ( .A1(n31252), .A2(n39154), .B1(n31316), .B2(n39148), .C1(
        n31188), .C2(n39142), .ZN(n36283) );
  AOI221_X1 U28929 ( .B1(n39166), .B2(n31069), .C1(n39160), .C2(n31133), .A(
        n36264), .ZN(n36263) );
  OAI222_X1 U28930 ( .A1(n31251), .A2(n39154), .B1(n31315), .B2(n39148), .C1(
        n31187), .C2(n39142), .ZN(n36264) );
  AOI221_X1 U28931 ( .B1(n39166), .B2(n31068), .C1(n39160), .C2(n31132), .A(
        n36245), .ZN(n36244) );
  OAI222_X1 U28932 ( .A1(n31250), .A2(n39154), .B1(n31314), .B2(n39148), .C1(
        n31186), .C2(n39142), .ZN(n36245) );
  AOI221_X1 U28933 ( .B1(n39166), .B2(n31067), .C1(n39160), .C2(n31131), .A(
        n36226), .ZN(n36225) );
  OAI222_X1 U28934 ( .A1(n31249), .A2(n39154), .B1(n31313), .B2(n39148), .C1(
        n31185), .C2(n39142), .ZN(n36226) );
  AOI221_X1 U28935 ( .B1(n39167), .B2(n31060), .C1(n39161), .C2(n31124), .A(
        n36093), .ZN(n36092) );
  OAI222_X1 U28936 ( .A1(n31242), .A2(n39155), .B1(n31306), .B2(n39149), .C1(
        n31178), .C2(n39143), .ZN(n36093) );
  AOI221_X1 U28937 ( .B1(n39167), .B2(n31059), .C1(n39161), .C2(n31123), .A(
        n36074), .ZN(n36073) );
  OAI222_X1 U28938 ( .A1(n31241), .A2(n39155), .B1(n31305), .B2(n39149), .C1(
        n31177), .C2(n39143), .ZN(n36074) );
  AOI221_X1 U28939 ( .B1(n39167), .B2(n31058), .C1(n39161), .C2(n31122), .A(
        n36055), .ZN(n36054) );
  OAI222_X1 U28940 ( .A1(n31240), .A2(n39155), .B1(n31304), .B2(n39149), .C1(
        n31176), .C2(n39143), .ZN(n36055) );
  AOI221_X1 U28941 ( .B1(n39167), .B2(n31057), .C1(n39161), .C2(n31121), .A(
        n36018), .ZN(n36015) );
  OAI222_X1 U28942 ( .A1(n31239), .A2(n39155), .B1(n31303), .B2(n39149), .C1(
        n31175), .C2(n39143), .ZN(n36018) );
  AOI221_X1 U28943 ( .B1(n39162), .B2(n31110), .C1(n39156), .C2(n31174), .A(
        n37043), .ZN(n37042) );
  OAI222_X1 U28944 ( .A1(n31292), .A2(n39150), .B1(n31356), .B2(n39144), .C1(
        n31228), .C2(n39138), .ZN(n37043) );
  AOI221_X1 U28945 ( .B1(n39166), .B2(n31066), .C1(n39160), .C2(n31130), .A(
        n36207), .ZN(n36206) );
  OAI222_X1 U28946 ( .A1(n31248), .A2(n39154), .B1(n31312), .B2(n39148), .C1(
        n31184), .C2(n39142), .ZN(n36207) );
  AOI221_X1 U28947 ( .B1(n39166), .B2(n31065), .C1(n39160), .C2(n31129), .A(
        n36188), .ZN(n36187) );
  OAI222_X1 U28948 ( .A1(n31247), .A2(n39154), .B1(n31311), .B2(n39148), .C1(
        n31183), .C2(n39142), .ZN(n36188) );
  AOI221_X1 U28949 ( .B1(n39166), .B2(n31064), .C1(n39160), .C2(n31128), .A(
        n36169), .ZN(n36168) );
  OAI222_X1 U28950 ( .A1(n31246), .A2(n39154), .B1(n31310), .B2(n39148), .C1(
        n31182), .C2(n39142), .ZN(n36169) );
  AOI221_X1 U28951 ( .B1(n39166), .B2(n31063), .C1(n39160), .C2(n31127), .A(
        n36150), .ZN(n36149) );
  OAI222_X1 U28952 ( .A1(n31245), .A2(n39154), .B1(n31309), .B2(n39148), .C1(
        n31181), .C2(n39142), .ZN(n36150) );
  AOI221_X1 U28953 ( .B1(n39166), .B2(n31062), .C1(n39160), .C2(n31126), .A(
        n36131), .ZN(n36130) );
  OAI222_X1 U28954 ( .A1(n31244), .A2(n39154), .B1(n31308), .B2(n39148), .C1(
        n31180), .C2(n39142), .ZN(n36131) );
  AOI221_X1 U28955 ( .B1(n39166), .B2(n31061), .C1(n39160), .C2(n31125), .A(
        n36112), .ZN(n36111) );
  OAI222_X1 U28956 ( .A1(n31243), .A2(n39154), .B1(n31307), .B2(n39148), .C1(
        n31179), .C2(n39142), .ZN(n36112) );
  AOI221_X1 U28957 ( .B1(n39668), .B2(n31110), .C1(n39662), .C2(n31174), .A(
        n33671), .ZN(n33670) );
  OAI222_X1 U28958 ( .A1(n31292), .A2(n39656), .B1(n31356), .B2(n39650), .C1(
        n31228), .C2(n39644), .ZN(n33671) );
  AOI221_X1 U28959 ( .B1(n39416), .B2(n31110), .C1(n39410), .C2(n31174), .A(
        n34945), .ZN(n34944) );
  OAI222_X1 U28960 ( .A1(n31292), .A2(n39404), .B1(n31356), .B2(n39398), .C1(
        n31228), .C2(n39392), .ZN(n34945) );
  AOI221_X1 U28961 ( .B1(n39668), .B2(n31109), .C1(n39662), .C2(n31173), .A(
        n33690), .ZN(n33689) );
  OAI222_X1 U28962 ( .A1(n31291), .A2(n39656), .B1(n31355), .B2(n39650), .C1(
        n31227), .C2(n39644), .ZN(n33690) );
  AOI221_X1 U28963 ( .B1(n39416), .B2(n31109), .C1(n39410), .C2(n31173), .A(
        n34964), .ZN(n34963) );
  OAI222_X1 U28964 ( .A1(n31291), .A2(n39404), .B1(n31355), .B2(n39398), .C1(
        n31227), .C2(n39392), .ZN(n34964) );
  AOI221_X1 U28965 ( .B1(n39668), .B2(n31108), .C1(n39662), .C2(n31172), .A(
        n33709), .ZN(n33708) );
  OAI222_X1 U28966 ( .A1(n31290), .A2(n39656), .B1(n31354), .B2(n39650), .C1(
        n31226), .C2(n39644), .ZN(n33709) );
  AOI221_X1 U28967 ( .B1(n39416), .B2(n31108), .C1(n39410), .C2(n31172), .A(
        n34983), .ZN(n34982) );
  OAI222_X1 U28968 ( .A1(n31290), .A2(n39404), .B1(n31354), .B2(n39398), .C1(
        n31226), .C2(n39392), .ZN(n34983) );
  AOI221_X1 U28969 ( .B1(n39668), .B2(n31107), .C1(n39662), .C2(n31171), .A(
        n33728), .ZN(n33727) );
  OAI222_X1 U28970 ( .A1(n31289), .A2(n39656), .B1(n31353), .B2(n39650), .C1(
        n31225), .C2(n39644), .ZN(n33728) );
  AOI221_X1 U28971 ( .B1(n39416), .B2(n31107), .C1(n39410), .C2(n31171), .A(
        n35002), .ZN(n35001) );
  OAI222_X1 U28972 ( .A1(n31289), .A2(n39404), .B1(n31353), .B2(n39398), .C1(
        n31225), .C2(n39392), .ZN(n35002) );
  AOI221_X1 U28973 ( .B1(n39668), .B2(n31106), .C1(n39662), .C2(n31170), .A(
        n33747), .ZN(n33746) );
  OAI222_X1 U28974 ( .A1(n31288), .A2(n39656), .B1(n31352), .B2(n39650), .C1(
        n31224), .C2(n39644), .ZN(n33747) );
  AOI221_X1 U28975 ( .B1(n39416), .B2(n31106), .C1(n39410), .C2(n31170), .A(
        n35021), .ZN(n35020) );
  OAI222_X1 U28976 ( .A1(n31288), .A2(n39404), .B1(n31352), .B2(n39398), .C1(
        n31224), .C2(n39392), .ZN(n35021) );
  AOI221_X1 U28977 ( .B1(n39668), .B2(n31105), .C1(n39662), .C2(n31169), .A(
        n33766), .ZN(n33765) );
  OAI222_X1 U28978 ( .A1(n31287), .A2(n39656), .B1(n31351), .B2(n39650), .C1(
        n31223), .C2(n39644), .ZN(n33766) );
  AOI221_X1 U28979 ( .B1(n39416), .B2(n31105), .C1(n39410), .C2(n31169), .A(
        n35040), .ZN(n35039) );
  OAI222_X1 U28980 ( .A1(n31287), .A2(n39404), .B1(n31351), .B2(n39398), .C1(
        n31223), .C2(n39392), .ZN(n35040) );
  AOI221_X1 U28981 ( .B1(n39667), .B2(n31104), .C1(n39661), .C2(n31168), .A(
        n33785), .ZN(n33784) );
  OAI222_X1 U28982 ( .A1(n31286), .A2(n39655), .B1(n31350), .B2(n39649), .C1(
        n31222), .C2(n39643), .ZN(n33785) );
  AOI221_X1 U28983 ( .B1(n39415), .B2(n31104), .C1(n39409), .C2(n31168), .A(
        n35059), .ZN(n35058) );
  OAI222_X1 U28984 ( .A1(n31286), .A2(n39403), .B1(n31350), .B2(n39397), .C1(
        n31222), .C2(n39391), .ZN(n35059) );
  AOI221_X1 U28985 ( .B1(n39667), .B2(n31103), .C1(n39661), .C2(n31167), .A(
        n33804), .ZN(n33803) );
  OAI222_X1 U28986 ( .A1(n31285), .A2(n39655), .B1(n31349), .B2(n39649), .C1(
        n31221), .C2(n39643), .ZN(n33804) );
  AOI221_X1 U28987 ( .B1(n39415), .B2(n31103), .C1(n39409), .C2(n31167), .A(
        n35078), .ZN(n35077) );
  OAI222_X1 U28988 ( .A1(n31285), .A2(n39403), .B1(n31349), .B2(n39397), .C1(
        n31221), .C2(n39391), .ZN(n35078) );
  AOI221_X1 U28989 ( .B1(n39667), .B2(n31102), .C1(n39661), .C2(n31166), .A(
        n33823), .ZN(n33822) );
  OAI222_X1 U28990 ( .A1(n31284), .A2(n39655), .B1(n31348), .B2(n39649), .C1(
        n31220), .C2(n39643), .ZN(n33823) );
  AOI221_X1 U28991 ( .B1(n39415), .B2(n31102), .C1(n39409), .C2(n31166), .A(
        n35097), .ZN(n35096) );
  OAI222_X1 U28992 ( .A1(n31284), .A2(n39403), .B1(n31348), .B2(n39397), .C1(
        n31220), .C2(n39391), .ZN(n35097) );
  AOI221_X1 U28993 ( .B1(n39667), .B2(n31101), .C1(n39661), .C2(n31165), .A(
        n33842), .ZN(n33841) );
  OAI222_X1 U28994 ( .A1(n31283), .A2(n39655), .B1(n31347), .B2(n39649), .C1(
        n31219), .C2(n39643), .ZN(n33842) );
  AOI221_X1 U28995 ( .B1(n39415), .B2(n31101), .C1(n39409), .C2(n31165), .A(
        n35116), .ZN(n35115) );
  OAI222_X1 U28996 ( .A1(n31283), .A2(n39403), .B1(n31347), .B2(n39397), .C1(
        n31219), .C2(n39391), .ZN(n35116) );
  AOI221_X1 U28997 ( .B1(n39667), .B2(n31100), .C1(n39661), .C2(n31164), .A(
        n33861), .ZN(n33860) );
  OAI222_X1 U28998 ( .A1(n31282), .A2(n39655), .B1(n31346), .B2(n39649), .C1(
        n31218), .C2(n39643), .ZN(n33861) );
  AOI221_X1 U28999 ( .B1(n39415), .B2(n31100), .C1(n39409), .C2(n31164), .A(
        n35135), .ZN(n35134) );
  OAI222_X1 U29000 ( .A1(n31282), .A2(n39403), .B1(n31346), .B2(n39397), .C1(
        n31218), .C2(n39391), .ZN(n35135) );
  AOI221_X1 U29001 ( .B1(n39667), .B2(n31099), .C1(n39661), .C2(n31163), .A(
        n33880), .ZN(n33879) );
  OAI222_X1 U29002 ( .A1(n31281), .A2(n39655), .B1(n31345), .B2(n39649), .C1(
        n31217), .C2(n39643), .ZN(n33880) );
  AOI221_X1 U29003 ( .B1(n39415), .B2(n31099), .C1(n39409), .C2(n31163), .A(
        n35154), .ZN(n35153) );
  OAI222_X1 U29004 ( .A1(n31281), .A2(n39403), .B1(n31345), .B2(n39397), .C1(
        n31217), .C2(n39391), .ZN(n35154) );
  AOI221_X1 U29005 ( .B1(n39667), .B2(n31098), .C1(n39661), .C2(n31162), .A(
        n33899), .ZN(n33898) );
  OAI222_X1 U29006 ( .A1(n31280), .A2(n39655), .B1(n31344), .B2(n39649), .C1(
        n31216), .C2(n39643), .ZN(n33899) );
  AOI221_X1 U29007 ( .B1(n39415), .B2(n31098), .C1(n39409), .C2(n31162), .A(
        n35173), .ZN(n35172) );
  OAI222_X1 U29008 ( .A1(n31280), .A2(n39403), .B1(n31344), .B2(n39397), .C1(
        n31216), .C2(n39391), .ZN(n35173) );
  AOI221_X1 U29009 ( .B1(n39667), .B2(n31097), .C1(n39661), .C2(n31161), .A(
        n33918), .ZN(n33917) );
  OAI222_X1 U29010 ( .A1(n31279), .A2(n39655), .B1(n31343), .B2(n39649), .C1(
        n31215), .C2(n39643), .ZN(n33918) );
  AOI221_X1 U29011 ( .B1(n39415), .B2(n31097), .C1(n39409), .C2(n31161), .A(
        n35192), .ZN(n35191) );
  OAI222_X1 U29012 ( .A1(n31279), .A2(n39403), .B1(n31343), .B2(n39397), .C1(
        n31215), .C2(n39391), .ZN(n35192) );
  AOI221_X1 U29013 ( .B1(n39667), .B2(n31096), .C1(n39661), .C2(n31160), .A(
        n33937), .ZN(n33936) );
  OAI222_X1 U29014 ( .A1(n31278), .A2(n39655), .B1(n31342), .B2(n39649), .C1(
        n31214), .C2(n39643), .ZN(n33937) );
  AOI221_X1 U29015 ( .B1(n39415), .B2(n31096), .C1(n39409), .C2(n31160), .A(
        n35211), .ZN(n35210) );
  OAI222_X1 U29016 ( .A1(n31278), .A2(n39403), .B1(n31342), .B2(n39397), .C1(
        n31214), .C2(n39391), .ZN(n35211) );
  AOI221_X1 U29017 ( .B1(n39667), .B2(n31095), .C1(n39661), .C2(n31159), .A(
        n33956), .ZN(n33955) );
  OAI222_X1 U29018 ( .A1(n31277), .A2(n39655), .B1(n31341), .B2(n39649), .C1(
        n31213), .C2(n39643), .ZN(n33956) );
  AOI221_X1 U29019 ( .B1(n39415), .B2(n31095), .C1(n39409), .C2(n31159), .A(
        n35230), .ZN(n35229) );
  OAI222_X1 U29020 ( .A1(n31277), .A2(n39403), .B1(n31341), .B2(n39397), .C1(
        n31213), .C2(n39391), .ZN(n35230) );
  AOI221_X1 U29021 ( .B1(n39667), .B2(n31094), .C1(n39661), .C2(n31158), .A(
        n33975), .ZN(n33974) );
  OAI222_X1 U29022 ( .A1(n31276), .A2(n39655), .B1(n31340), .B2(n39649), .C1(
        n31212), .C2(n39643), .ZN(n33975) );
  AOI221_X1 U29023 ( .B1(n39415), .B2(n31094), .C1(n39409), .C2(n31158), .A(
        n35249), .ZN(n35248) );
  OAI222_X1 U29024 ( .A1(n31276), .A2(n39403), .B1(n31340), .B2(n39397), .C1(
        n31212), .C2(n39391), .ZN(n35249) );
  AOI221_X1 U29025 ( .B1(n39667), .B2(n31093), .C1(n39661), .C2(n31157), .A(
        n33994), .ZN(n33993) );
  OAI222_X1 U29026 ( .A1(n31275), .A2(n39655), .B1(n31339), .B2(n39649), .C1(
        n31211), .C2(n39643), .ZN(n33994) );
  AOI221_X1 U29027 ( .B1(n39415), .B2(n31093), .C1(n39409), .C2(n31157), .A(
        n35268), .ZN(n35267) );
  OAI222_X1 U29028 ( .A1(n31275), .A2(n39403), .B1(n31339), .B2(n39397), .C1(
        n31211), .C2(n39391), .ZN(n35268) );
  AOI221_X1 U29029 ( .B1(n39666), .B2(n31092), .C1(n39660), .C2(n31156), .A(
        n34013), .ZN(n34012) );
  OAI222_X1 U29030 ( .A1(n31274), .A2(n39654), .B1(n31338), .B2(n39648), .C1(
        n31210), .C2(n39642), .ZN(n34013) );
  AOI221_X1 U29031 ( .B1(n39414), .B2(n31092), .C1(n39408), .C2(n31156), .A(
        n35287), .ZN(n35286) );
  OAI222_X1 U29032 ( .A1(n31274), .A2(n39402), .B1(n31338), .B2(n39396), .C1(
        n31210), .C2(n39390), .ZN(n35287) );
  AOI221_X1 U29033 ( .B1(n39666), .B2(n31091), .C1(n39660), .C2(n31155), .A(
        n34032), .ZN(n34031) );
  OAI222_X1 U29034 ( .A1(n31273), .A2(n39654), .B1(n31337), .B2(n39648), .C1(
        n31209), .C2(n39642), .ZN(n34032) );
  AOI221_X1 U29035 ( .B1(n39414), .B2(n31091), .C1(n39408), .C2(n31155), .A(
        n35306), .ZN(n35305) );
  OAI222_X1 U29036 ( .A1(n31273), .A2(n39402), .B1(n31337), .B2(n39396), .C1(
        n31209), .C2(n39390), .ZN(n35306) );
  AOI221_X1 U29037 ( .B1(n39666), .B2(n31090), .C1(n39660), .C2(n31154), .A(
        n34051), .ZN(n34050) );
  OAI222_X1 U29038 ( .A1(n31272), .A2(n39654), .B1(n31336), .B2(n39648), .C1(
        n31208), .C2(n39642), .ZN(n34051) );
  AOI221_X1 U29039 ( .B1(n39414), .B2(n31090), .C1(n39408), .C2(n31154), .A(
        n35325), .ZN(n35324) );
  OAI222_X1 U29040 ( .A1(n31272), .A2(n39402), .B1(n31336), .B2(n39396), .C1(
        n31208), .C2(n39390), .ZN(n35325) );
  AOI221_X1 U29041 ( .B1(n39666), .B2(n31089), .C1(n39660), .C2(n31153), .A(
        n34070), .ZN(n34069) );
  OAI222_X1 U29042 ( .A1(n31271), .A2(n39654), .B1(n31335), .B2(n39648), .C1(
        n31207), .C2(n39642), .ZN(n34070) );
  AOI221_X1 U29043 ( .B1(n39414), .B2(n31089), .C1(n39408), .C2(n31153), .A(
        n35344), .ZN(n35343) );
  OAI222_X1 U29044 ( .A1(n31271), .A2(n39402), .B1(n31335), .B2(n39396), .C1(
        n31207), .C2(n39390), .ZN(n35344) );
  AOI221_X1 U29045 ( .B1(n39666), .B2(n31088), .C1(n39660), .C2(n31152), .A(
        n34089), .ZN(n34088) );
  OAI222_X1 U29046 ( .A1(n31270), .A2(n39654), .B1(n31334), .B2(n39648), .C1(
        n31206), .C2(n39642), .ZN(n34089) );
  AOI221_X1 U29047 ( .B1(n39414), .B2(n31088), .C1(n39408), .C2(n31152), .A(
        n35363), .ZN(n35362) );
  OAI222_X1 U29048 ( .A1(n31270), .A2(n39402), .B1(n31334), .B2(n39396), .C1(
        n31206), .C2(n39390), .ZN(n35363) );
  AOI221_X1 U29049 ( .B1(n39666), .B2(n31087), .C1(n39660), .C2(n31151), .A(
        n34108), .ZN(n34107) );
  OAI222_X1 U29050 ( .A1(n31269), .A2(n39654), .B1(n31333), .B2(n39648), .C1(
        n31205), .C2(n39642), .ZN(n34108) );
  AOI221_X1 U29051 ( .B1(n39414), .B2(n31087), .C1(n39408), .C2(n31151), .A(
        n35382), .ZN(n35381) );
  OAI222_X1 U29052 ( .A1(n31269), .A2(n39402), .B1(n31333), .B2(n39396), .C1(
        n31205), .C2(n39390), .ZN(n35382) );
  AOI221_X1 U29053 ( .B1(n39666), .B2(n31086), .C1(n39660), .C2(n31150), .A(
        n34127), .ZN(n34126) );
  OAI222_X1 U29054 ( .A1(n31268), .A2(n39654), .B1(n31332), .B2(n39648), .C1(
        n31204), .C2(n39642), .ZN(n34127) );
  AOI221_X1 U29055 ( .B1(n39414), .B2(n31086), .C1(n39408), .C2(n31150), .A(
        n35401), .ZN(n35400) );
  OAI222_X1 U29056 ( .A1(n31268), .A2(n39402), .B1(n31332), .B2(n39396), .C1(
        n31204), .C2(n39390), .ZN(n35401) );
  AOI221_X1 U29057 ( .B1(n39666), .B2(n31085), .C1(n39660), .C2(n31149), .A(
        n34146), .ZN(n34145) );
  OAI222_X1 U29058 ( .A1(n31267), .A2(n39654), .B1(n31331), .B2(n39648), .C1(
        n31203), .C2(n39642), .ZN(n34146) );
  AOI221_X1 U29059 ( .B1(n39414), .B2(n31085), .C1(n39408), .C2(n31149), .A(
        n35420), .ZN(n35419) );
  OAI222_X1 U29060 ( .A1(n31267), .A2(n39402), .B1(n31331), .B2(n39396), .C1(
        n31203), .C2(n39390), .ZN(n35420) );
  AOI221_X1 U29061 ( .B1(n39666), .B2(n31084), .C1(n39660), .C2(n31148), .A(
        n34165), .ZN(n34164) );
  OAI222_X1 U29062 ( .A1(n31266), .A2(n39654), .B1(n31330), .B2(n39648), .C1(
        n31202), .C2(n39642), .ZN(n34165) );
  AOI221_X1 U29063 ( .B1(n39414), .B2(n31084), .C1(n39408), .C2(n31148), .A(
        n35439), .ZN(n35438) );
  OAI222_X1 U29064 ( .A1(n31266), .A2(n39402), .B1(n31330), .B2(n39396), .C1(
        n31202), .C2(n39390), .ZN(n35439) );
  AOI221_X1 U29065 ( .B1(n39666), .B2(n31083), .C1(n39660), .C2(n31147), .A(
        n34184), .ZN(n34183) );
  OAI222_X1 U29066 ( .A1(n31265), .A2(n39654), .B1(n31329), .B2(n39648), .C1(
        n31201), .C2(n39642), .ZN(n34184) );
  AOI221_X1 U29067 ( .B1(n39414), .B2(n31083), .C1(n39408), .C2(n31147), .A(
        n35458), .ZN(n35457) );
  OAI222_X1 U29068 ( .A1(n31265), .A2(n39402), .B1(n31329), .B2(n39396), .C1(
        n31201), .C2(n39390), .ZN(n35458) );
  AOI221_X1 U29069 ( .B1(n39666), .B2(n31082), .C1(n39660), .C2(n31146), .A(
        n34203), .ZN(n34202) );
  OAI222_X1 U29070 ( .A1(n31264), .A2(n39654), .B1(n31328), .B2(n39648), .C1(
        n31200), .C2(n39642), .ZN(n34203) );
  AOI221_X1 U29071 ( .B1(n39414), .B2(n31082), .C1(n39408), .C2(n31146), .A(
        n35477), .ZN(n35476) );
  OAI222_X1 U29072 ( .A1(n31264), .A2(n39402), .B1(n31328), .B2(n39396), .C1(
        n31200), .C2(n39390), .ZN(n35477) );
  AOI221_X1 U29073 ( .B1(n39666), .B2(n31081), .C1(n39660), .C2(n31145), .A(
        n34222), .ZN(n34221) );
  OAI222_X1 U29074 ( .A1(n31263), .A2(n39654), .B1(n31327), .B2(n39648), .C1(
        n31199), .C2(n39642), .ZN(n34222) );
  AOI221_X1 U29075 ( .B1(n39414), .B2(n31081), .C1(n39408), .C2(n31145), .A(
        n35496), .ZN(n35495) );
  OAI222_X1 U29076 ( .A1(n31263), .A2(n39402), .B1(n31327), .B2(n39396), .C1(
        n31199), .C2(n39390), .ZN(n35496) );
  AOI221_X1 U29077 ( .B1(n39665), .B2(n31080), .C1(n39659), .C2(n31144), .A(
        n34241), .ZN(n34240) );
  OAI222_X1 U29078 ( .A1(n31262), .A2(n39653), .B1(n31326), .B2(n39647), .C1(
        n31198), .C2(n39641), .ZN(n34241) );
  AOI221_X1 U29079 ( .B1(n39413), .B2(n31080), .C1(n39407), .C2(n31144), .A(
        n35515), .ZN(n35514) );
  OAI222_X1 U29080 ( .A1(n31262), .A2(n39401), .B1(n31326), .B2(n39395), .C1(
        n31198), .C2(n39389), .ZN(n35515) );
  AOI221_X1 U29081 ( .B1(n39665), .B2(n31079), .C1(n39659), .C2(n31143), .A(
        n34260), .ZN(n34259) );
  OAI222_X1 U29082 ( .A1(n31261), .A2(n39653), .B1(n31325), .B2(n39647), .C1(
        n31197), .C2(n39641), .ZN(n34260) );
  AOI221_X1 U29083 ( .B1(n39413), .B2(n31079), .C1(n39407), .C2(n31143), .A(
        n35534), .ZN(n35533) );
  OAI222_X1 U29084 ( .A1(n31261), .A2(n39401), .B1(n31325), .B2(n39395), .C1(
        n31197), .C2(n39389), .ZN(n35534) );
  AOI221_X1 U29085 ( .B1(n39665), .B2(n31078), .C1(n39659), .C2(n31142), .A(
        n34279), .ZN(n34278) );
  OAI222_X1 U29086 ( .A1(n31260), .A2(n39653), .B1(n31324), .B2(n39647), .C1(
        n31196), .C2(n39641), .ZN(n34279) );
  AOI221_X1 U29087 ( .B1(n39413), .B2(n31078), .C1(n39407), .C2(n31142), .A(
        n35553), .ZN(n35552) );
  OAI222_X1 U29088 ( .A1(n31260), .A2(n39401), .B1(n31324), .B2(n39395), .C1(
        n31196), .C2(n39389), .ZN(n35553) );
  AOI221_X1 U29089 ( .B1(n39665), .B2(n31077), .C1(n39659), .C2(n31141), .A(
        n34298), .ZN(n34297) );
  OAI222_X1 U29090 ( .A1(n31259), .A2(n39653), .B1(n31323), .B2(n39647), .C1(
        n31195), .C2(n39641), .ZN(n34298) );
  AOI221_X1 U29091 ( .B1(n39413), .B2(n31077), .C1(n39407), .C2(n31141), .A(
        n35572), .ZN(n35571) );
  OAI222_X1 U29092 ( .A1(n31259), .A2(n39401), .B1(n31323), .B2(n39395), .C1(
        n31195), .C2(n39389), .ZN(n35572) );
  AOI221_X1 U29093 ( .B1(n39665), .B2(n31076), .C1(n39659), .C2(n31140), .A(
        n34317), .ZN(n34316) );
  OAI222_X1 U29094 ( .A1(n31258), .A2(n39653), .B1(n31322), .B2(n39647), .C1(
        n31194), .C2(n39641), .ZN(n34317) );
  AOI221_X1 U29095 ( .B1(n39413), .B2(n31076), .C1(n39407), .C2(n31140), .A(
        n35591), .ZN(n35590) );
  OAI222_X1 U29096 ( .A1(n31258), .A2(n39401), .B1(n31322), .B2(n39395), .C1(
        n31194), .C2(n39389), .ZN(n35591) );
  AOI221_X1 U29097 ( .B1(n39665), .B2(n31075), .C1(n39659), .C2(n31139), .A(
        n34336), .ZN(n34335) );
  OAI222_X1 U29098 ( .A1(n31257), .A2(n39653), .B1(n31321), .B2(n39647), .C1(
        n31193), .C2(n39641), .ZN(n34336) );
  AOI221_X1 U29099 ( .B1(n39413), .B2(n31075), .C1(n39407), .C2(n31139), .A(
        n35610), .ZN(n35609) );
  OAI222_X1 U29100 ( .A1(n31257), .A2(n39401), .B1(n31321), .B2(n39395), .C1(
        n31193), .C2(n39389), .ZN(n35610) );
  AOI221_X1 U29101 ( .B1(n39665), .B2(n31074), .C1(n39659), .C2(n31138), .A(
        n34355), .ZN(n34354) );
  OAI222_X1 U29102 ( .A1(n31256), .A2(n39653), .B1(n31320), .B2(n39647), .C1(
        n31192), .C2(n39641), .ZN(n34355) );
  AOI221_X1 U29103 ( .B1(n39413), .B2(n31074), .C1(n39407), .C2(n31138), .A(
        n35629), .ZN(n35628) );
  OAI222_X1 U29104 ( .A1(n31256), .A2(n39401), .B1(n31320), .B2(n39395), .C1(
        n31192), .C2(n39389), .ZN(n35629) );
  AOI221_X1 U29105 ( .B1(n39665), .B2(n31073), .C1(n39659), .C2(n31137), .A(
        n34374), .ZN(n34373) );
  OAI222_X1 U29106 ( .A1(n31255), .A2(n39653), .B1(n31319), .B2(n39647), .C1(
        n31191), .C2(n39641), .ZN(n34374) );
  AOI221_X1 U29107 ( .B1(n39413), .B2(n31073), .C1(n39407), .C2(n31137), .A(
        n35648), .ZN(n35647) );
  OAI222_X1 U29108 ( .A1(n31255), .A2(n39401), .B1(n31319), .B2(n39395), .C1(
        n31191), .C2(n39389), .ZN(n35648) );
  AOI221_X1 U29109 ( .B1(n39665), .B2(n31072), .C1(n39659), .C2(n31136), .A(
        n34393), .ZN(n34392) );
  OAI222_X1 U29110 ( .A1(n31254), .A2(n39653), .B1(n31318), .B2(n39647), .C1(
        n31190), .C2(n39641), .ZN(n34393) );
  AOI221_X1 U29111 ( .B1(n39413), .B2(n31072), .C1(n39407), .C2(n31136), .A(
        n35667), .ZN(n35666) );
  OAI222_X1 U29112 ( .A1(n31254), .A2(n39401), .B1(n31318), .B2(n39395), .C1(
        n31190), .C2(n39389), .ZN(n35667) );
  AOI221_X1 U29113 ( .B1(n39665), .B2(n31071), .C1(n39659), .C2(n31135), .A(
        n34412), .ZN(n34411) );
  OAI222_X1 U29114 ( .A1(n31253), .A2(n39653), .B1(n31317), .B2(n39647), .C1(
        n31189), .C2(n39641), .ZN(n34412) );
  AOI221_X1 U29115 ( .B1(n39413), .B2(n31071), .C1(n39407), .C2(n31135), .A(
        n35686), .ZN(n35685) );
  OAI222_X1 U29116 ( .A1(n31253), .A2(n39401), .B1(n31317), .B2(n39395), .C1(
        n31189), .C2(n39389), .ZN(n35686) );
  AOI221_X1 U29117 ( .B1(n39665), .B2(n31070), .C1(n39659), .C2(n31134), .A(
        n34431), .ZN(n34430) );
  OAI222_X1 U29118 ( .A1(n31252), .A2(n39653), .B1(n31316), .B2(n39647), .C1(
        n31188), .C2(n39641), .ZN(n34431) );
  AOI221_X1 U29119 ( .B1(n39413), .B2(n31070), .C1(n39407), .C2(n31134), .A(
        n35705), .ZN(n35704) );
  OAI222_X1 U29120 ( .A1(n31252), .A2(n39401), .B1(n31316), .B2(n39395), .C1(
        n31188), .C2(n39389), .ZN(n35705) );
  AOI221_X1 U29121 ( .B1(n39665), .B2(n31069), .C1(n39659), .C2(n31133), .A(
        n34450), .ZN(n34449) );
  OAI222_X1 U29122 ( .A1(n31251), .A2(n39653), .B1(n31315), .B2(n39647), .C1(
        n31187), .C2(n39641), .ZN(n34450) );
  AOI221_X1 U29123 ( .B1(n39413), .B2(n31069), .C1(n39407), .C2(n31133), .A(
        n35724), .ZN(n35723) );
  OAI222_X1 U29124 ( .A1(n31251), .A2(n39401), .B1(n31315), .B2(n39395), .C1(
        n31187), .C2(n39389), .ZN(n35724) );
  AOI221_X1 U29125 ( .B1(n39664), .B2(n31068), .C1(n39658), .C2(n31132), .A(
        n34469), .ZN(n34468) );
  OAI222_X1 U29126 ( .A1(n31250), .A2(n39652), .B1(n31314), .B2(n39646), .C1(
        n31186), .C2(n39640), .ZN(n34469) );
  AOI221_X1 U29127 ( .B1(n39412), .B2(n31068), .C1(n39406), .C2(n31132), .A(
        n35743), .ZN(n35742) );
  OAI222_X1 U29128 ( .A1(n31250), .A2(n39400), .B1(n31314), .B2(n39394), .C1(
        n31186), .C2(n39388), .ZN(n35743) );
  AOI221_X1 U29129 ( .B1(n39664), .B2(n31067), .C1(n39658), .C2(n31131), .A(
        n34488), .ZN(n34487) );
  OAI222_X1 U29130 ( .A1(n31249), .A2(n39652), .B1(n31313), .B2(n39646), .C1(
        n31185), .C2(n39640), .ZN(n34488) );
  AOI221_X1 U29131 ( .B1(n39412), .B2(n31067), .C1(n39406), .C2(n31131), .A(
        n35762), .ZN(n35761) );
  OAI222_X1 U29132 ( .A1(n31249), .A2(n39400), .B1(n31313), .B2(n39394), .C1(
        n31185), .C2(n39388), .ZN(n35762) );
  AOI221_X1 U29133 ( .B1(n39664), .B2(n31066), .C1(n39658), .C2(n31130), .A(
        n34507), .ZN(n34506) );
  OAI222_X1 U29134 ( .A1(n31248), .A2(n39652), .B1(n31312), .B2(n39646), .C1(
        n31184), .C2(n39640), .ZN(n34507) );
  AOI221_X1 U29135 ( .B1(n39412), .B2(n31066), .C1(n39406), .C2(n31130), .A(
        n35781), .ZN(n35780) );
  OAI222_X1 U29136 ( .A1(n31248), .A2(n39400), .B1(n31312), .B2(n39394), .C1(
        n31184), .C2(n39388), .ZN(n35781) );
  AOI221_X1 U29137 ( .B1(n39664), .B2(n31065), .C1(n39658), .C2(n31129), .A(
        n34526), .ZN(n34525) );
  OAI222_X1 U29138 ( .A1(n31247), .A2(n39652), .B1(n31311), .B2(n39646), .C1(
        n31183), .C2(n39640), .ZN(n34526) );
  AOI221_X1 U29139 ( .B1(n39412), .B2(n31065), .C1(n39406), .C2(n31129), .A(
        n35800), .ZN(n35799) );
  OAI222_X1 U29140 ( .A1(n31247), .A2(n39400), .B1(n31311), .B2(n39394), .C1(
        n31183), .C2(n39388), .ZN(n35800) );
  AOI221_X1 U29141 ( .B1(n39664), .B2(n31064), .C1(n39658), .C2(n31128), .A(
        n34545), .ZN(n34544) );
  OAI222_X1 U29142 ( .A1(n31246), .A2(n39652), .B1(n31310), .B2(n39646), .C1(
        n31182), .C2(n39640), .ZN(n34545) );
  AOI221_X1 U29143 ( .B1(n39412), .B2(n31064), .C1(n39406), .C2(n31128), .A(
        n35819), .ZN(n35818) );
  OAI222_X1 U29144 ( .A1(n31246), .A2(n39400), .B1(n31310), .B2(n39394), .C1(
        n31182), .C2(n39388), .ZN(n35819) );
  AOI221_X1 U29145 ( .B1(n39664), .B2(n31063), .C1(n39658), .C2(n31127), .A(
        n34564), .ZN(n34563) );
  OAI222_X1 U29146 ( .A1(n31245), .A2(n39652), .B1(n31309), .B2(n39646), .C1(
        n31181), .C2(n39640), .ZN(n34564) );
  AOI221_X1 U29147 ( .B1(n39412), .B2(n31063), .C1(n39406), .C2(n31127), .A(
        n35838), .ZN(n35837) );
  OAI222_X1 U29148 ( .A1(n31245), .A2(n39400), .B1(n31309), .B2(n39394), .C1(
        n31181), .C2(n39388), .ZN(n35838) );
  AOI221_X1 U29149 ( .B1(n39664), .B2(n31062), .C1(n39658), .C2(n31126), .A(
        n34583), .ZN(n34582) );
  OAI222_X1 U29150 ( .A1(n31244), .A2(n39652), .B1(n31308), .B2(n39646), .C1(
        n31180), .C2(n39640), .ZN(n34583) );
  AOI221_X1 U29151 ( .B1(n39412), .B2(n31062), .C1(n39406), .C2(n31126), .A(
        n35857), .ZN(n35856) );
  OAI222_X1 U29152 ( .A1(n31244), .A2(n39400), .B1(n31308), .B2(n39394), .C1(
        n31180), .C2(n39388), .ZN(n35857) );
  AOI221_X1 U29153 ( .B1(n39664), .B2(n31061), .C1(n39658), .C2(n31125), .A(
        n34602), .ZN(n34601) );
  OAI222_X1 U29154 ( .A1(n31243), .A2(n39652), .B1(n31307), .B2(n39646), .C1(
        n31179), .C2(n39640), .ZN(n34602) );
  AOI221_X1 U29155 ( .B1(n39412), .B2(n31061), .C1(n39406), .C2(n31125), .A(
        n35876), .ZN(n35875) );
  OAI222_X1 U29156 ( .A1(n31243), .A2(n39400), .B1(n31307), .B2(n39394), .C1(
        n31179), .C2(n39388), .ZN(n35876) );
  AOI221_X1 U29157 ( .B1(n39664), .B2(n31060), .C1(n39658), .C2(n31124), .A(
        n34621), .ZN(n34620) );
  OAI222_X1 U29158 ( .A1(n31242), .A2(n39652), .B1(n31306), .B2(n39646), .C1(
        n31178), .C2(n39640), .ZN(n34621) );
  AOI221_X1 U29159 ( .B1(n39412), .B2(n31060), .C1(n39406), .C2(n31124), .A(
        n35895), .ZN(n35894) );
  OAI222_X1 U29160 ( .A1(n31242), .A2(n39400), .B1(n31306), .B2(n39394), .C1(
        n31178), .C2(n39388), .ZN(n35895) );
  AOI221_X1 U29161 ( .B1(n39664), .B2(n31059), .C1(n39658), .C2(n31123), .A(
        n34640), .ZN(n34639) );
  OAI222_X1 U29162 ( .A1(n31241), .A2(n39652), .B1(n31305), .B2(n39646), .C1(
        n31177), .C2(n39640), .ZN(n34640) );
  AOI221_X1 U29163 ( .B1(n39412), .B2(n31059), .C1(n39406), .C2(n31123), .A(
        n35914), .ZN(n35913) );
  OAI222_X1 U29164 ( .A1(n31241), .A2(n39400), .B1(n31305), .B2(n39394), .C1(
        n31177), .C2(n39388), .ZN(n35914) );
  AOI221_X1 U29165 ( .B1(n39664), .B2(n31058), .C1(n39658), .C2(n31122), .A(
        n34659), .ZN(n34658) );
  OAI222_X1 U29166 ( .A1(n31240), .A2(n39652), .B1(n31304), .B2(n39646), .C1(
        n31176), .C2(n39640), .ZN(n34659) );
  AOI221_X1 U29167 ( .B1(n39412), .B2(n31058), .C1(n39406), .C2(n31122), .A(
        n35933), .ZN(n35932) );
  OAI222_X1 U29168 ( .A1(n31240), .A2(n39400), .B1(n31304), .B2(n39394), .C1(
        n31176), .C2(n39388), .ZN(n35933) );
  AOI221_X1 U29169 ( .B1(n39664), .B2(n31057), .C1(n39658), .C2(n31121), .A(
        n34689), .ZN(n34688) );
  OAI222_X1 U29170 ( .A1(n31239), .A2(n39652), .B1(n31303), .B2(n39646), .C1(
        n31175), .C2(n39640), .ZN(n34689) );
  AOI221_X1 U29171 ( .B1(n39412), .B2(n31057), .C1(n39406), .C2(n31121), .A(
        n35963), .ZN(n35962) );
  OAI222_X1 U29172 ( .A1(n31239), .A2(n39400), .B1(n31303), .B2(n39394), .C1(
        n31175), .C2(n39388), .ZN(n35963) );
  AOI221_X1 U29173 ( .B1(n39132), .B2(n32815), .C1(n39126), .C2(n32767), .A(
        n37025), .ZN(n37022) );
  OAI222_X1 U29174 ( .A1(n30981), .A2(n39120), .B1(n31045), .B2(n39114), .C1(
        n30917), .C2(n39108), .ZN(n37025) );
  AOI221_X1 U29175 ( .B1(n39133), .B2(n32814), .C1(n39127), .C2(n32766), .A(
        n37006), .ZN(n37003) );
  OAI222_X1 U29176 ( .A1(n30980), .A2(n39121), .B1(n31044), .B2(n39115), .C1(
        n30916), .C2(n39109), .ZN(n37006) );
  AOI221_X1 U29177 ( .B1(n39133), .B2(n32813), .C1(n39127), .C2(n32765), .A(
        n36987), .ZN(n36984) );
  OAI222_X1 U29178 ( .A1(n30979), .A2(n39121), .B1(n31043), .B2(n39115), .C1(
        n30915), .C2(n39109), .ZN(n36987) );
  AOI221_X1 U29179 ( .B1(n39133), .B2(n32812), .C1(n39127), .C2(n32764), .A(
        n36968), .ZN(n36965) );
  OAI222_X1 U29180 ( .A1(n30978), .A2(n39121), .B1(n31042), .B2(n39115), .C1(
        n30914), .C2(n39109), .ZN(n36968) );
  AOI221_X1 U29181 ( .B1(n39133), .B2(n32811), .C1(n39127), .C2(n32763), .A(
        n36949), .ZN(n36946) );
  OAI222_X1 U29182 ( .A1(n30977), .A2(n39121), .B1(n31041), .B2(n39115), .C1(
        n30913), .C2(n39109), .ZN(n36949) );
  AOI221_X1 U29183 ( .B1(n39133), .B2(n32810), .C1(n39127), .C2(n32762), .A(
        n36930), .ZN(n36927) );
  OAI222_X1 U29184 ( .A1(n30976), .A2(n39121), .B1(n31040), .B2(n39115), .C1(
        n30912), .C2(n39109), .ZN(n36930) );
  AOI221_X1 U29185 ( .B1(n39133), .B2(n32809), .C1(n39127), .C2(n32761), .A(
        n36911), .ZN(n36908) );
  OAI222_X1 U29186 ( .A1(n30975), .A2(n39121), .B1(n31039), .B2(n39115), .C1(
        n30911), .C2(n39109), .ZN(n36911) );
  AOI221_X1 U29187 ( .B1(n39133), .B2(n32808), .C1(n39127), .C2(n32760), .A(
        n36892), .ZN(n36889) );
  OAI222_X1 U29188 ( .A1(n30974), .A2(n39121), .B1(n31038), .B2(n39115), .C1(
        n30910), .C2(n39109), .ZN(n36892) );
  AOI221_X1 U29189 ( .B1(n39133), .B2(n32807), .C1(n39127), .C2(n32759), .A(
        n36873), .ZN(n36870) );
  OAI222_X1 U29190 ( .A1(n30973), .A2(n39121), .B1(n31037), .B2(n39115), .C1(
        n30909), .C2(n39109), .ZN(n36873) );
  AOI221_X1 U29191 ( .B1(n39133), .B2(n32806), .C1(n39127), .C2(n32758), .A(
        n36854), .ZN(n36851) );
  OAI222_X1 U29192 ( .A1(n30972), .A2(n39121), .B1(n31036), .B2(n39115), .C1(
        n30908), .C2(n39109), .ZN(n36854) );
  AOI221_X1 U29193 ( .B1(n39133), .B2(n32805), .C1(n39127), .C2(n32757), .A(
        n36835), .ZN(n36832) );
  OAI222_X1 U29194 ( .A1(n30971), .A2(n39121), .B1(n31035), .B2(n39115), .C1(
        n30907), .C2(n39109), .ZN(n36835) );
  AOI221_X1 U29195 ( .B1(n39133), .B2(n32804), .C1(n39127), .C2(n32756), .A(
        n36816), .ZN(n36813) );
  OAI222_X1 U29196 ( .A1(n30970), .A2(n39121), .B1(n31034), .B2(n39115), .C1(
        n30906), .C2(n39109), .ZN(n36816) );
  AOI221_X1 U29197 ( .B1(n39133), .B2(n32803), .C1(n39127), .C2(n32755), .A(
        n36797), .ZN(n36794) );
  OAI222_X1 U29198 ( .A1(n30969), .A2(n39121), .B1(n31033), .B2(n39115), .C1(
        n30905), .C2(n39109), .ZN(n36797) );
  AOI221_X1 U29199 ( .B1(n39134), .B2(n32802), .C1(n39128), .C2(n32754), .A(
        n36778), .ZN(n36775) );
  OAI222_X1 U29200 ( .A1(n30968), .A2(n39122), .B1(n31032), .B2(n39116), .C1(
        n30904), .C2(n39110), .ZN(n36778) );
  AOI221_X1 U29201 ( .B1(n39134), .B2(n32801), .C1(n39128), .C2(n32753), .A(
        n36759), .ZN(n36756) );
  OAI222_X1 U29202 ( .A1(n30967), .A2(n39122), .B1(n31031), .B2(n39116), .C1(
        n30903), .C2(n39110), .ZN(n36759) );
  AOI221_X1 U29203 ( .B1(n39134), .B2(n32800), .C1(n39128), .C2(n32752), .A(
        n36740), .ZN(n36737) );
  OAI222_X1 U29204 ( .A1(n30966), .A2(n39122), .B1(n31030), .B2(n39116), .C1(
        n30902), .C2(n39110), .ZN(n36740) );
  AOI221_X1 U29205 ( .B1(n39134), .B2(n32799), .C1(n39128), .C2(n32751), .A(
        n36721), .ZN(n36718) );
  OAI222_X1 U29206 ( .A1(n30965), .A2(n39122), .B1(n31029), .B2(n39116), .C1(
        n30901), .C2(n39110), .ZN(n36721) );
  AOI221_X1 U29207 ( .B1(n39134), .B2(n32798), .C1(n39128), .C2(n32750), .A(
        n36702), .ZN(n36699) );
  OAI222_X1 U29208 ( .A1(n30964), .A2(n39122), .B1(n31028), .B2(n39116), .C1(
        n30900), .C2(n39110), .ZN(n36702) );
  AOI221_X1 U29209 ( .B1(n39134), .B2(n32797), .C1(n39128), .C2(n32749), .A(
        n36683), .ZN(n36680) );
  OAI222_X1 U29210 ( .A1(n30963), .A2(n39122), .B1(n31027), .B2(n39116), .C1(
        n30899), .C2(n39110), .ZN(n36683) );
  AOI221_X1 U29211 ( .B1(n39134), .B2(n32796), .C1(n39128), .C2(n32748), .A(
        n36664), .ZN(n36661) );
  OAI222_X1 U29212 ( .A1(n30962), .A2(n39122), .B1(n31026), .B2(n39116), .C1(
        n30898), .C2(n39110), .ZN(n36664) );
  AOI221_X1 U29213 ( .B1(n39134), .B2(n32795), .C1(n39128), .C2(n32747), .A(
        n36645), .ZN(n36642) );
  OAI222_X1 U29214 ( .A1(n30961), .A2(n39122), .B1(n31025), .B2(n39116), .C1(
        n30897), .C2(n39110), .ZN(n36645) );
  AOI221_X1 U29215 ( .B1(n39134), .B2(n32794), .C1(n39128), .C2(n32746), .A(
        n36626), .ZN(n36623) );
  OAI222_X1 U29216 ( .A1(n30960), .A2(n39122), .B1(n31024), .B2(n39116), .C1(
        n30896), .C2(n39110), .ZN(n36626) );
  AOI221_X1 U29217 ( .B1(n39134), .B2(n32793), .C1(n39128), .C2(n32745), .A(
        n36607), .ZN(n36604) );
  OAI222_X1 U29218 ( .A1(n30959), .A2(n39122), .B1(n31023), .B2(n39116), .C1(
        n30895), .C2(n39110), .ZN(n36607) );
  AOI221_X1 U29219 ( .B1(n39134), .B2(n32792), .C1(n39128), .C2(n32744), .A(
        n36588), .ZN(n36585) );
  OAI222_X1 U29220 ( .A1(n30958), .A2(n39122), .B1(n31022), .B2(n39116), .C1(
        n30894), .C2(n39110), .ZN(n36588) );
  AOI221_X1 U29221 ( .B1(n39134), .B2(n32791), .C1(n39128), .C2(n32743), .A(
        n36569), .ZN(n36566) );
  OAI222_X1 U29222 ( .A1(n30957), .A2(n39122), .B1(n31021), .B2(n39116), .C1(
        n30893), .C2(n39110), .ZN(n36569) );
  AOI221_X1 U29223 ( .B1(n39135), .B2(n32790), .C1(n39129), .C2(n32742), .A(
        n36550), .ZN(n36547) );
  OAI222_X1 U29224 ( .A1(n30956), .A2(n39123), .B1(n31020), .B2(n39117), .C1(
        n30892), .C2(n39111), .ZN(n36550) );
  AOI221_X1 U29225 ( .B1(n39135), .B2(n32789), .C1(n39129), .C2(n32741), .A(
        n36531), .ZN(n36528) );
  OAI222_X1 U29226 ( .A1(n30955), .A2(n39123), .B1(n31019), .B2(n39117), .C1(
        n30891), .C2(n39111), .ZN(n36531) );
  AOI221_X1 U29227 ( .B1(n39135), .B2(n32788), .C1(n39129), .C2(n32740), .A(
        n36512), .ZN(n36509) );
  OAI222_X1 U29228 ( .A1(n30954), .A2(n39123), .B1(n31018), .B2(n39117), .C1(
        n30890), .C2(n39111), .ZN(n36512) );
  AOI221_X1 U29229 ( .B1(n39135), .B2(n32787), .C1(n39129), .C2(n32739), .A(
        n36493), .ZN(n36490) );
  OAI222_X1 U29230 ( .A1(n30953), .A2(n39123), .B1(n31017), .B2(n39117), .C1(
        n30889), .C2(n39111), .ZN(n36493) );
  AOI221_X1 U29231 ( .B1(n39135), .B2(n32786), .C1(n39129), .C2(n32738), .A(
        n36474), .ZN(n36471) );
  OAI222_X1 U29232 ( .A1(n30952), .A2(n39123), .B1(n31016), .B2(n39117), .C1(
        n30888), .C2(n39111), .ZN(n36474) );
  AOI221_X1 U29233 ( .B1(n39135), .B2(n32785), .C1(n39129), .C2(n32737), .A(
        n36455), .ZN(n36452) );
  OAI222_X1 U29234 ( .A1(n30951), .A2(n39123), .B1(n31015), .B2(n39117), .C1(
        n30887), .C2(n39111), .ZN(n36455) );
  AOI221_X1 U29235 ( .B1(n39135), .B2(n32784), .C1(n39129), .C2(n32736), .A(
        n36436), .ZN(n36433) );
  OAI222_X1 U29236 ( .A1(n30950), .A2(n39123), .B1(n31014), .B2(n39117), .C1(
        n30886), .C2(n39111), .ZN(n36436) );
  AOI221_X1 U29237 ( .B1(n39135), .B2(n32783), .C1(n39129), .C2(n32735), .A(
        n36417), .ZN(n36414) );
  OAI222_X1 U29238 ( .A1(n30949), .A2(n39123), .B1(n31013), .B2(n39117), .C1(
        n30885), .C2(n39111), .ZN(n36417) );
  AOI221_X1 U29239 ( .B1(n39135), .B2(n32782), .C1(n39129), .C2(n32734), .A(
        n36398), .ZN(n36395) );
  OAI222_X1 U29240 ( .A1(n30948), .A2(n39123), .B1(n31012), .B2(n39117), .C1(
        n30884), .C2(n39111), .ZN(n36398) );
  AOI221_X1 U29241 ( .B1(n39135), .B2(n32781), .C1(n39129), .C2(n32733), .A(
        n36379), .ZN(n36376) );
  OAI222_X1 U29242 ( .A1(n30947), .A2(n39123), .B1(n31011), .B2(n39117), .C1(
        n30883), .C2(n39111), .ZN(n36379) );
  AOI221_X1 U29243 ( .B1(n39135), .B2(n32780), .C1(n39129), .C2(n32732), .A(
        n36360), .ZN(n36357) );
  OAI222_X1 U29244 ( .A1(n30946), .A2(n39123), .B1(n31010), .B2(n39117), .C1(
        n30882), .C2(n39111), .ZN(n36360) );
  AOI221_X1 U29245 ( .B1(n39135), .B2(n32779), .C1(n39129), .C2(n32731), .A(
        n36341), .ZN(n36338) );
  OAI222_X1 U29246 ( .A1(n30945), .A2(n39123), .B1(n31009), .B2(n39117), .C1(
        n30881), .C2(n39111), .ZN(n36341) );
  AOI221_X1 U29247 ( .B1(n39136), .B2(n32778), .C1(n39130), .C2(n32730), .A(
        n36322), .ZN(n36319) );
  OAI222_X1 U29248 ( .A1(n30944), .A2(n39124), .B1(n31008), .B2(n39118), .C1(
        n30880), .C2(n39112), .ZN(n36322) );
  AOI221_X1 U29249 ( .B1(n39136), .B2(n32777), .C1(n39130), .C2(n32729), .A(
        n36303), .ZN(n36300) );
  OAI222_X1 U29250 ( .A1(n30943), .A2(n39124), .B1(n31007), .B2(n39118), .C1(
        n30879), .C2(n39112), .ZN(n36303) );
  AOI221_X1 U29251 ( .B1(n39136), .B2(n32776), .C1(n39130), .C2(n32728), .A(
        n36284), .ZN(n36281) );
  OAI222_X1 U29252 ( .A1(n30942), .A2(n39124), .B1(n31006), .B2(n39118), .C1(
        n30878), .C2(n39112), .ZN(n36284) );
  AOI221_X1 U29253 ( .B1(n39136), .B2(n32775), .C1(n39130), .C2(n32727), .A(
        n36265), .ZN(n36262) );
  OAI222_X1 U29254 ( .A1(n30941), .A2(n39124), .B1(n31005), .B2(n39118), .C1(
        n30877), .C2(n39112), .ZN(n36265) );
  AOI221_X1 U29255 ( .B1(n39136), .B2(n32846), .C1(n39130), .C2(n32834), .A(
        n36246), .ZN(n36243) );
  OAI222_X1 U29256 ( .A1(n30940), .A2(n39124), .B1(n31004), .B2(n39118), .C1(
        n30876), .C2(n39112), .ZN(n36246) );
  AOI221_X1 U29257 ( .B1(n39136), .B2(n32845), .C1(n39130), .C2(n32833), .A(
        n36227), .ZN(n36224) );
  OAI222_X1 U29258 ( .A1(n30939), .A2(n39124), .B1(n31003), .B2(n39118), .C1(
        n30875), .C2(n39112), .ZN(n36227) );
  AOI221_X1 U29259 ( .B1(n39132), .B2(n32474), .C1(n39126), .C2(n32470), .A(
        n37215), .ZN(n37212) );
  OAI222_X1 U29260 ( .A1(n30991), .A2(n39120), .B1(n31055), .B2(n39114), .C1(
        n30927), .C2(n39108), .ZN(n37215) );
  AOI221_X1 U29261 ( .B1(n39132), .B2(n32473), .C1(n39126), .C2(n32469), .A(
        n37196), .ZN(n37193) );
  OAI222_X1 U29262 ( .A1(n30990), .A2(n39120), .B1(n31054), .B2(n39114), .C1(
        n30926), .C2(n39108), .ZN(n37196) );
  AOI221_X1 U29263 ( .B1(n39132), .B2(n32472), .C1(n39126), .C2(n32468), .A(
        n37177), .ZN(n37174) );
  OAI222_X1 U29264 ( .A1(n30989), .A2(n39120), .B1(n31053), .B2(n39114), .C1(
        n30925), .C2(n39108), .ZN(n37177) );
  AOI221_X1 U29265 ( .B1(n39132), .B2(n32822), .C1(n39126), .C2(n32774), .A(
        n37158), .ZN(n37155) );
  OAI222_X1 U29266 ( .A1(n30988), .A2(n39120), .B1(n31052), .B2(n39114), .C1(
        n30924), .C2(n39108), .ZN(n37158) );
  AOI221_X1 U29267 ( .B1(n39132), .B2(n32821), .C1(n39126), .C2(n32773), .A(
        n37139), .ZN(n37136) );
  OAI222_X1 U29268 ( .A1(n30987), .A2(n39120), .B1(n31051), .B2(n39114), .C1(
        n30923), .C2(n39108), .ZN(n37139) );
  AOI221_X1 U29269 ( .B1(n39137), .B2(n32838), .C1(n39131), .C2(n32826), .A(
        n36094), .ZN(n36091) );
  OAI222_X1 U29270 ( .A1(n30932), .A2(n39125), .B1(n30996), .B2(n39119), .C1(
        n30868), .C2(n39113), .ZN(n36094) );
  AOI221_X1 U29271 ( .B1(n39137), .B2(n32837), .C1(n39131), .C2(n32825), .A(
        n36075), .ZN(n36072) );
  OAI222_X1 U29272 ( .A1(n30931), .A2(n39125), .B1(n30995), .B2(n39119), .C1(
        n30867), .C2(n39113), .ZN(n36075) );
  AOI221_X1 U29273 ( .B1(n39137), .B2(n32836), .C1(n39131), .C2(n32824), .A(
        n36056), .ZN(n36053) );
  OAI222_X1 U29274 ( .A1(n30930), .A2(n39125), .B1(n30994), .B2(n39119), .C1(
        n30866), .C2(n39113), .ZN(n36056) );
  AOI221_X1 U29275 ( .B1(n39137), .B2(n32835), .C1(n39131), .C2(n32823), .A(
        n36024), .ZN(n36014) );
  OAI222_X1 U29276 ( .A1(n30929), .A2(n39125), .B1(n30993), .B2(n39119), .C1(
        n30865), .C2(n39113), .ZN(n36024) );
  AOI221_X1 U29277 ( .B1(n39132), .B2(n32475), .C1(n39126), .C2(n32471), .A(
        n37247), .ZN(n37243) );
  OAI222_X1 U29278 ( .A1(n30992), .A2(n39120), .B1(n31056), .B2(n39114), .C1(
        n30928), .C2(n39108), .ZN(n37247) );
  AOI221_X1 U29279 ( .B1(n39132), .B2(n32820), .C1(n39126), .C2(n32772), .A(
        n37120), .ZN(n37117) );
  OAI222_X1 U29280 ( .A1(n30986), .A2(n39120), .B1(n31050), .B2(n39114), .C1(
        n30922), .C2(n39108), .ZN(n37120) );
  AOI221_X1 U29281 ( .B1(n39132), .B2(n32819), .C1(n39126), .C2(n32771), .A(
        n37101), .ZN(n37098) );
  OAI222_X1 U29282 ( .A1(n30985), .A2(n39120), .B1(n31049), .B2(n39114), .C1(
        n30921), .C2(n39108), .ZN(n37101) );
  AOI221_X1 U29283 ( .B1(n39132), .B2(n32818), .C1(n39126), .C2(n32770), .A(
        n37082), .ZN(n37079) );
  OAI222_X1 U29284 ( .A1(n30984), .A2(n39120), .B1(n31048), .B2(n39114), .C1(
        n30920), .C2(n39108), .ZN(n37082) );
  AOI221_X1 U29285 ( .B1(n39132), .B2(n32817), .C1(n39126), .C2(n32769), .A(
        n37063), .ZN(n37060) );
  OAI222_X1 U29286 ( .A1(n30983), .A2(n39120), .B1(n31047), .B2(n39114), .C1(
        n30919), .C2(n39108), .ZN(n37063) );
  AOI221_X1 U29287 ( .B1(n39132), .B2(n32816), .C1(n39126), .C2(n32768), .A(
        n37044), .ZN(n37041) );
  OAI222_X1 U29288 ( .A1(n30982), .A2(n39120), .B1(n31046), .B2(n39114), .C1(
        n30918), .C2(n39108), .ZN(n37044) );
  AOI221_X1 U29289 ( .B1(n39136), .B2(n32844), .C1(n39130), .C2(n32832), .A(
        n36208), .ZN(n36205) );
  OAI222_X1 U29290 ( .A1(n30938), .A2(n39124), .B1(n31002), .B2(n39118), .C1(
        n30874), .C2(n39112), .ZN(n36208) );
  AOI221_X1 U29291 ( .B1(n39136), .B2(n32843), .C1(n39130), .C2(n32831), .A(
        n36189), .ZN(n36186) );
  OAI222_X1 U29292 ( .A1(n30937), .A2(n39124), .B1(n31001), .B2(n39118), .C1(
        n30873), .C2(n39112), .ZN(n36189) );
  AOI221_X1 U29293 ( .B1(n39136), .B2(n32842), .C1(n39130), .C2(n32830), .A(
        n36170), .ZN(n36167) );
  OAI222_X1 U29294 ( .A1(n30936), .A2(n39124), .B1(n31000), .B2(n39118), .C1(
        n30872), .C2(n39112), .ZN(n36170) );
  AOI221_X1 U29295 ( .B1(n39136), .B2(n32841), .C1(n39130), .C2(n32829), .A(
        n36151), .ZN(n36148) );
  OAI222_X1 U29296 ( .A1(n30935), .A2(n39124), .B1(n30999), .B2(n39118), .C1(
        n30871), .C2(n39112), .ZN(n36151) );
  AOI221_X1 U29297 ( .B1(n39136), .B2(n32840), .C1(n39130), .C2(n32828), .A(
        n36132), .ZN(n36129) );
  OAI222_X1 U29298 ( .A1(n30934), .A2(n39124), .B1(n30998), .B2(n39118), .C1(
        n30870), .C2(n39112), .ZN(n36132) );
  AOI221_X1 U29299 ( .B1(n39136), .B2(n32839), .C1(n39130), .C2(n32827), .A(
        n36113), .ZN(n36110) );
  OAI222_X1 U29300 ( .A1(n30933), .A2(n39124), .B1(n30997), .B2(n39118), .C1(
        n30869), .C2(n39112), .ZN(n36113) );
  AOI221_X1 U29301 ( .B1(n39639), .B2(n32475), .C1(n39633), .C2(n32471), .A(
        n33469), .ZN(n33459) );
  OAI222_X1 U29302 ( .A1(n30992), .A2(n39627), .B1(n31056), .B2(n39621), .C1(
        n30928), .C2(n39615), .ZN(n33469) );
  AOI221_X1 U29303 ( .B1(n39387), .B2(n32475), .C1(n39381), .C2(n32471), .A(
        n34743), .ZN(n34733) );
  OAI222_X1 U29304 ( .A1(n30992), .A2(n39375), .B1(n31056), .B2(n39369), .C1(
        n30928), .C2(n39363), .ZN(n34743) );
  AOI221_X1 U29305 ( .B1(n39639), .B2(n32474), .C1(n39633), .C2(n32470), .A(
        n33501), .ZN(n33498) );
  OAI222_X1 U29306 ( .A1(n30991), .A2(n39627), .B1(n31055), .B2(n39621), .C1(
        n30927), .C2(n39615), .ZN(n33501) );
  AOI221_X1 U29307 ( .B1(n39387), .B2(n32474), .C1(n39381), .C2(n32470), .A(
        n34775), .ZN(n34772) );
  OAI222_X1 U29308 ( .A1(n30991), .A2(n39375), .B1(n31055), .B2(n39369), .C1(
        n30927), .C2(n39363), .ZN(n34775) );
  AOI221_X1 U29309 ( .B1(n39639), .B2(n32473), .C1(n39633), .C2(n32469), .A(
        n33520), .ZN(n33517) );
  OAI222_X1 U29310 ( .A1(n30990), .A2(n39627), .B1(n31054), .B2(n39621), .C1(
        n30926), .C2(n39615), .ZN(n33520) );
  AOI221_X1 U29311 ( .B1(n39387), .B2(n32473), .C1(n39381), .C2(n32469), .A(
        n34794), .ZN(n34791) );
  OAI222_X1 U29312 ( .A1(n30990), .A2(n39375), .B1(n31054), .B2(n39369), .C1(
        n30926), .C2(n39363), .ZN(n34794) );
  AOI221_X1 U29313 ( .B1(n39639), .B2(n32472), .C1(n39633), .C2(n32468), .A(
        n33539), .ZN(n33536) );
  OAI222_X1 U29314 ( .A1(n30989), .A2(n39627), .B1(n31053), .B2(n39621), .C1(
        n30925), .C2(n39615), .ZN(n33539) );
  AOI221_X1 U29315 ( .B1(n39387), .B2(n32472), .C1(n39381), .C2(n32468), .A(
        n34813), .ZN(n34810) );
  OAI222_X1 U29316 ( .A1(n30989), .A2(n39375), .B1(n31053), .B2(n39369), .C1(
        n30925), .C2(n39363), .ZN(n34813) );
  OAI222_X1 U29317 ( .A1(n40593), .A2(n40745), .B1(n40586), .B2(n41129), .C1(
        n40577), .C2(n32321), .ZN(n9866) );
  OAI222_X1 U29318 ( .A1(n40593), .A2(n40751), .B1(n40586), .B2(n41135), .C1(
        n40578), .C2(n32320), .ZN(n9865) );
  OAI222_X1 U29319 ( .A1(n40593), .A2(n40757), .B1(n40586), .B2(n41141), .C1(
        n40578), .C2(n32319), .ZN(n9864) );
  OAI222_X1 U29320 ( .A1(n40593), .A2(n40763), .B1(n40586), .B2(n41147), .C1(
        n40578), .C2(n32318), .ZN(n9863) );
  OAI222_X1 U29321 ( .A1(n40592), .A2(n40769), .B1(n40585), .B2(n41153), .C1(
        n40578), .C2(n32317), .ZN(n9862) );
  OAI222_X1 U29322 ( .A1(n40592), .A2(n40775), .B1(n40585), .B2(n41159), .C1(
        n40578), .C2(n32316), .ZN(n9861) );
  OAI222_X1 U29323 ( .A1(n40592), .A2(n40781), .B1(n40585), .B2(n41165), .C1(
        n40578), .C2(n32315), .ZN(n9860) );
  OAI222_X1 U29324 ( .A1(n40592), .A2(n40787), .B1(n40585), .B2(n41171), .C1(
        n40578), .C2(n32314), .ZN(n9859) );
  OAI222_X1 U29325 ( .A1(n40592), .A2(n40793), .B1(n40585), .B2(n41177), .C1(
        n40578), .C2(n32313), .ZN(n9858) );
  OAI222_X1 U29326 ( .A1(n40592), .A2(n40799), .B1(n40585), .B2(n41183), .C1(
        n40578), .C2(n32312), .ZN(n9857) );
  OAI222_X1 U29327 ( .A1(n40592), .A2(n40805), .B1(n40585), .B2(n41189), .C1(
        n40578), .C2(n32311), .ZN(n9856) );
  OAI222_X1 U29328 ( .A1(n40592), .A2(n40811), .B1(n40585), .B2(n41195), .C1(
        n40578), .C2(n32310), .ZN(n9855) );
  OAI222_X1 U29329 ( .A1(n40592), .A2(n40817), .B1(n40585), .B2(n41201), .C1(
        n40579), .C2(n32309), .ZN(n9854) );
  OAI222_X1 U29330 ( .A1(n40592), .A2(n40823), .B1(n40585), .B2(n41207), .C1(
        n40579), .C2(n32308), .ZN(n9853) );
  OAI222_X1 U29331 ( .A1(n40592), .A2(n40829), .B1(n40585), .B2(n41213), .C1(
        n40579), .C2(n32307), .ZN(n9852) );
  OAI222_X1 U29332 ( .A1(n40592), .A2(n40835), .B1(n40585), .B2(n41219), .C1(
        n40579), .C2(n32306), .ZN(n9851) );
  OAI222_X1 U29333 ( .A1(n40591), .A2(n40841), .B1(n40584), .B2(n41225), .C1(
        n40579), .C2(n32305), .ZN(n9850) );
  OAI222_X1 U29334 ( .A1(n40591), .A2(n40847), .B1(n40584), .B2(n41231), .C1(
        n40579), .C2(n32304), .ZN(n9849) );
  OAI222_X1 U29335 ( .A1(n40591), .A2(n40853), .B1(n40584), .B2(n41237), .C1(
        n40579), .C2(n32303), .ZN(n9848) );
  OAI222_X1 U29336 ( .A1(n40591), .A2(n40859), .B1(n40584), .B2(n41243), .C1(
        n40579), .C2(n32302), .ZN(n9847) );
  OAI222_X1 U29337 ( .A1(n40591), .A2(n40865), .B1(n40584), .B2(n41249), .C1(
        n40579), .C2(n32301), .ZN(n9846) );
  OAI222_X1 U29338 ( .A1(n40591), .A2(n40871), .B1(n40584), .B2(n41255), .C1(
        n40579), .C2(n32300), .ZN(n9845) );
  OAI222_X1 U29339 ( .A1(n40591), .A2(n40877), .B1(n40584), .B2(n41261), .C1(
        n40579), .C2(n32299), .ZN(n9844) );
  OAI222_X1 U29340 ( .A1(n40591), .A2(n40883), .B1(n40584), .B2(n41267), .C1(
        n40579), .C2(n32298), .ZN(n9843) );
  OAI222_X1 U29341 ( .A1(n40591), .A2(n40889), .B1(n40584), .B2(n41273), .C1(
        n40580), .C2(n32297), .ZN(n9842) );
  OAI222_X1 U29342 ( .A1(n40591), .A2(n40895), .B1(n40584), .B2(n41279), .C1(
        n40580), .C2(n32296), .ZN(n9841) );
  OAI222_X1 U29343 ( .A1(n40591), .A2(n40901), .B1(n40584), .B2(n41285), .C1(
        n40580), .C2(n32295), .ZN(n9840) );
  OAI222_X1 U29344 ( .A1(n40591), .A2(n40907), .B1(n40584), .B2(n41291), .C1(
        n40580), .C2(n32294), .ZN(n9839) );
  OAI222_X1 U29345 ( .A1(n40590), .A2(n40913), .B1(n40583), .B2(n41297), .C1(
        n40580), .C2(n32293), .ZN(n9838) );
  OAI222_X1 U29346 ( .A1(n40590), .A2(n40919), .B1(n40583), .B2(n41303), .C1(
        n40580), .C2(n32292), .ZN(n9837) );
  OAI222_X1 U29347 ( .A1(n40590), .A2(n40925), .B1(n40583), .B2(n41309), .C1(
        n40580), .C2(n32291), .ZN(n9836) );
  OAI222_X1 U29348 ( .A1(n40590), .A2(n40931), .B1(n40583), .B2(n41315), .C1(
        n40580), .C2(n32290), .ZN(n9835) );
  OAI222_X1 U29349 ( .A1(n40590), .A2(n40937), .B1(n40583), .B2(n41321), .C1(
        n40580), .C2(n32289), .ZN(n9834) );
  OAI222_X1 U29350 ( .A1(n40590), .A2(n40943), .B1(n40583), .B2(n41327), .C1(
        n40580), .C2(n32288), .ZN(n9833) );
  OAI222_X1 U29351 ( .A1(n40590), .A2(n40949), .B1(n40583), .B2(n41333), .C1(
        n40580), .C2(n32287), .ZN(n9832) );
  OAI222_X1 U29352 ( .A1(n40590), .A2(n40961), .B1(n40583), .B2(n41345), .C1(
        n40580), .C2(n32286), .ZN(n9830) );
  OAI222_X1 U29353 ( .A1(n40601), .A2(n40555), .B1(n40985), .B2(n40548), .C1(
        n40536), .C2(n32285), .ZN(n9762) );
  OAI222_X1 U29354 ( .A1(n40607), .A2(n40555), .B1(n40991), .B2(n40548), .C1(
        n40536), .C2(n32284), .ZN(n9761) );
  OAI222_X1 U29355 ( .A1(n40613), .A2(n40555), .B1(n40997), .B2(n40548), .C1(
        n40536), .C2(n32283), .ZN(n9760) );
  OAI222_X1 U29356 ( .A1(n40619), .A2(n40555), .B1(n41003), .B2(n40548), .C1(
        n40536), .C2(n32282), .ZN(n9759) );
  OAI222_X1 U29357 ( .A1(n40601), .A2(n40575), .B1(n40985), .B2(n40568), .C1(
        n40556), .C2(n32281), .ZN(n9826) );
  OAI222_X1 U29358 ( .A1(n40607), .A2(n40575), .B1(n40991), .B2(n40568), .C1(
        n40556), .C2(n32280), .ZN(n9825) );
  OAI222_X1 U29359 ( .A1(n40613), .A2(n40575), .B1(n40997), .B2(n40568), .C1(
        n40556), .C2(n32279), .ZN(n9824) );
  OAI222_X1 U29360 ( .A1(n40619), .A2(n40575), .B1(n41003), .B2(n40568), .C1(
        n40556), .C2(n32278), .ZN(n9823) );
  OAI222_X1 U29361 ( .A1(n40600), .A2(n40455), .B1(n40984), .B2(n40448), .C1(
        n40436), .C2(n32277), .ZN(n9442) );
  OAI222_X1 U29362 ( .A1(n40606), .A2(n40455), .B1(n40990), .B2(n40448), .C1(
        n40436), .C2(n32276), .ZN(n9441) );
  OAI222_X1 U29363 ( .A1(n40612), .A2(n40455), .B1(n40996), .B2(n40448), .C1(
        n40436), .C2(n32275), .ZN(n9440) );
  OAI222_X1 U29364 ( .A1(n40618), .A2(n40455), .B1(n41002), .B2(n40448), .C1(
        n40436), .C2(n32274), .ZN(n9439) );
  OAI222_X1 U29365 ( .A1(n40600), .A2(n40495), .B1(n40984), .B2(n40488), .C1(
        n40476), .C2(n32273), .ZN(n9570) );
  OAI222_X1 U29366 ( .A1(n40606), .A2(n40495), .B1(n40990), .B2(n40488), .C1(
        n40476), .C2(n32272), .ZN(n9569) );
  OAI222_X1 U29367 ( .A1(n40612), .A2(n40495), .B1(n40996), .B2(n40488), .C1(
        n40476), .C2(n32271), .ZN(n9568) );
  OAI222_X1 U29368 ( .A1(n40618), .A2(n40495), .B1(n41002), .B2(n40488), .C1(
        n40476), .C2(n32270), .ZN(n9567) );
  OAI222_X1 U29369 ( .A1(n40600), .A2(n40475), .B1(n40984), .B2(n40468), .C1(
        n40456), .C2(n32269), .ZN(n9506) );
  OAI222_X1 U29370 ( .A1(n40606), .A2(n40475), .B1(n40990), .B2(n40468), .C1(
        n40456), .C2(n32268), .ZN(n9505) );
  OAI222_X1 U29371 ( .A1(n40612), .A2(n40475), .B1(n40996), .B2(n40468), .C1(
        n40456), .C2(n32267), .ZN(n9504) );
  OAI222_X1 U29372 ( .A1(n40618), .A2(n40475), .B1(n41002), .B2(n40468), .C1(
        n40456), .C2(n32266), .ZN(n9503) );
  OAI222_X1 U29373 ( .A1(n40595), .A2(n40601), .B1(n40588), .B2(n40985), .C1(
        n40576), .C2(n32265), .ZN(n9890) );
  OAI222_X1 U29374 ( .A1(n40595), .A2(n40607), .B1(n40588), .B2(n40991), .C1(
        n40576), .C2(n32264), .ZN(n9889) );
  OAI222_X1 U29375 ( .A1(n40595), .A2(n40613), .B1(n40588), .B2(n40997), .C1(
        n40576), .C2(n32263), .ZN(n9888) );
  OAI222_X1 U29376 ( .A1(n40595), .A2(n40619), .B1(n40588), .B2(n41003), .C1(
        n40576), .C2(n32262), .ZN(n9887) );
  OAI222_X1 U29377 ( .A1(n40594), .A2(n40625), .B1(n40587), .B2(n41009), .C1(
        n40576), .C2(n32074), .ZN(n9886) );
  OAI222_X1 U29378 ( .A1(n40594), .A2(n40631), .B1(n40587), .B2(n41015), .C1(
        n40576), .C2(n32073), .ZN(n9885) );
  OAI222_X1 U29379 ( .A1(n40594), .A2(n40637), .B1(n40587), .B2(n41021), .C1(
        n40576), .C2(n32072), .ZN(n9884) );
  OAI222_X1 U29380 ( .A1(n40594), .A2(n40643), .B1(n40587), .B2(n41027), .C1(
        n40576), .C2(n32071), .ZN(n9883) );
  OAI222_X1 U29381 ( .A1(n40594), .A2(n40649), .B1(n40587), .B2(n41033), .C1(
        n40576), .C2(n32070), .ZN(n9882) );
  OAI222_X1 U29382 ( .A1(n40594), .A2(n40655), .B1(n40587), .B2(n41039), .C1(
        n40576), .C2(n32069), .ZN(n9881) );
  OAI222_X1 U29383 ( .A1(n40594), .A2(n40661), .B1(n40587), .B2(n41045), .C1(
        n40576), .C2(n32068), .ZN(n9880) );
  OAI222_X1 U29384 ( .A1(n40594), .A2(n40667), .B1(n40587), .B2(n41051), .C1(
        n40576), .C2(n32067), .ZN(n9879) );
  OAI222_X1 U29385 ( .A1(n40594), .A2(n40673), .B1(n40587), .B2(n41057), .C1(
        n40577), .C2(n32066), .ZN(n9878) );
  OAI222_X1 U29386 ( .A1(n40594), .A2(n40679), .B1(n40587), .B2(n41063), .C1(
        n40577), .C2(n32065), .ZN(n9877) );
  OAI222_X1 U29387 ( .A1(n40594), .A2(n40685), .B1(n40587), .B2(n41069), .C1(
        n40577), .C2(n32064), .ZN(n9876) );
  OAI222_X1 U29388 ( .A1(n40594), .A2(n40691), .B1(n40587), .B2(n41075), .C1(
        n40578), .C2(n32063), .ZN(n9875) );
  OAI222_X1 U29389 ( .A1(n40593), .A2(n40697), .B1(n40586), .B2(n41081), .C1(
        n40577), .C2(n32062), .ZN(n9874) );
  OAI222_X1 U29390 ( .A1(n40593), .A2(n40703), .B1(n40586), .B2(n41087), .C1(
        n40577), .C2(n32061), .ZN(n9873) );
  OAI222_X1 U29391 ( .A1(n40593), .A2(n40709), .B1(n40586), .B2(n41093), .C1(
        n40577), .C2(n32060), .ZN(n9872) );
  OAI222_X1 U29392 ( .A1(n40593), .A2(n40715), .B1(n40586), .B2(n41099), .C1(
        n40577), .C2(n32059), .ZN(n9871) );
  OAI222_X1 U29393 ( .A1(n40593), .A2(n40721), .B1(n40586), .B2(n41105), .C1(
        n40577), .C2(n32058), .ZN(n9870) );
  OAI222_X1 U29394 ( .A1(n40593), .A2(n40727), .B1(n40586), .B2(n41111), .C1(
        n40577), .C2(n32057), .ZN(n9869) );
  OAI222_X1 U29395 ( .A1(n40593), .A2(n40733), .B1(n40586), .B2(n41117), .C1(
        n40577), .C2(n32056), .ZN(n9868) );
  OAI222_X1 U29396 ( .A1(n40593), .A2(n40739), .B1(n40586), .B2(n41123), .C1(
        n40577), .C2(n32055), .ZN(n9867) );
  OAI222_X1 U29397 ( .A1(n40625), .A2(n40574), .B1(n41009), .B2(n40567), .C1(
        n40556), .C2(n32050), .ZN(n9822) );
  OAI222_X1 U29398 ( .A1(n40631), .A2(n40574), .B1(n41015), .B2(n40567), .C1(
        n40556), .C2(n32049), .ZN(n9821) );
  OAI222_X1 U29399 ( .A1(n40637), .A2(n40574), .B1(n41021), .B2(n40567), .C1(
        n40556), .C2(n32048), .ZN(n9820) );
  OAI222_X1 U29400 ( .A1(n40643), .A2(n40574), .B1(n41027), .B2(n40567), .C1(
        n40556), .C2(n32047), .ZN(n9819) );
  OAI222_X1 U29401 ( .A1(n40649), .A2(n40574), .B1(n41033), .B2(n40567), .C1(
        n40556), .C2(n32046), .ZN(n9818) );
  OAI222_X1 U29402 ( .A1(n40655), .A2(n40574), .B1(n41039), .B2(n40567), .C1(
        n40556), .C2(n32045), .ZN(n9817) );
  OAI222_X1 U29403 ( .A1(n40661), .A2(n40574), .B1(n41045), .B2(n40567), .C1(
        n40556), .C2(n32044), .ZN(n9816) );
  OAI222_X1 U29404 ( .A1(n40667), .A2(n40574), .B1(n41051), .B2(n40567), .C1(
        n40556), .C2(n32043), .ZN(n9815) );
  OAI222_X1 U29405 ( .A1(n40673), .A2(n40574), .B1(n41057), .B2(n40567), .C1(
        n40557), .C2(n32042), .ZN(n9814) );
  OAI222_X1 U29406 ( .A1(n40679), .A2(n40574), .B1(n41063), .B2(n40567), .C1(
        n40557), .C2(n32041), .ZN(n9813) );
  OAI222_X1 U29407 ( .A1(n40685), .A2(n40574), .B1(n41069), .B2(n40567), .C1(
        n40557), .C2(n32040), .ZN(n9812) );
  OAI222_X1 U29408 ( .A1(n40691), .A2(n40574), .B1(n41075), .B2(n40567), .C1(
        n40558), .C2(n32039), .ZN(n9811) );
  OAI222_X1 U29409 ( .A1(n40697), .A2(n40573), .B1(n41081), .B2(n40566), .C1(
        n40557), .C2(n32038), .ZN(n9810) );
  OAI222_X1 U29410 ( .A1(n40703), .A2(n40573), .B1(n41087), .B2(n40566), .C1(
        n40557), .C2(n32037), .ZN(n9809) );
  OAI222_X1 U29411 ( .A1(n40709), .A2(n40573), .B1(n41093), .B2(n40566), .C1(
        n40557), .C2(n32036), .ZN(n9808) );
  OAI222_X1 U29412 ( .A1(n40715), .A2(n40573), .B1(n41099), .B2(n40566), .C1(
        n40557), .C2(n32035), .ZN(n9807) );
  OAI222_X1 U29413 ( .A1(n40721), .A2(n40573), .B1(n41105), .B2(n40566), .C1(
        n40557), .C2(n32034), .ZN(n9806) );
  OAI222_X1 U29414 ( .A1(n40727), .A2(n40573), .B1(n41111), .B2(n40566), .C1(
        n40557), .C2(n32033), .ZN(n9805) );
  OAI222_X1 U29415 ( .A1(n40733), .A2(n40573), .B1(n41117), .B2(n40566), .C1(
        n40557), .C2(n32032), .ZN(n9804) );
  OAI222_X1 U29416 ( .A1(n40739), .A2(n40573), .B1(n41123), .B2(n40566), .C1(
        n40557), .C2(n32031), .ZN(n9803) );
  OAI222_X1 U29417 ( .A1(n40745), .A2(n40573), .B1(n41129), .B2(n40566), .C1(
        n40557), .C2(n32030), .ZN(n9802) );
  OAI222_X1 U29418 ( .A1(n40751), .A2(n40573), .B1(n41135), .B2(n40566), .C1(
        n40558), .C2(n32029), .ZN(n9801) );
  OAI222_X1 U29419 ( .A1(n40757), .A2(n40573), .B1(n41141), .B2(n40566), .C1(
        n40558), .C2(n32028), .ZN(n9800) );
  OAI222_X1 U29420 ( .A1(n40763), .A2(n40573), .B1(n41147), .B2(n40566), .C1(
        n40558), .C2(n32027), .ZN(n9799) );
  OAI222_X1 U29421 ( .A1(n40769), .A2(n40572), .B1(n41153), .B2(n40565), .C1(
        n40558), .C2(n32026), .ZN(n9798) );
  OAI222_X1 U29422 ( .A1(n40775), .A2(n40572), .B1(n41159), .B2(n40565), .C1(
        n40558), .C2(n32025), .ZN(n9797) );
  OAI222_X1 U29423 ( .A1(n40781), .A2(n40572), .B1(n41165), .B2(n40565), .C1(
        n40558), .C2(n32024), .ZN(n9796) );
  OAI222_X1 U29424 ( .A1(n40787), .A2(n40572), .B1(n41171), .B2(n40565), .C1(
        n40558), .C2(n32023), .ZN(n9795) );
  OAI222_X1 U29425 ( .A1(n40793), .A2(n40572), .B1(n41177), .B2(n40565), .C1(
        n40558), .C2(n32022), .ZN(n9794) );
  OAI222_X1 U29426 ( .A1(n40799), .A2(n40572), .B1(n41183), .B2(n40565), .C1(
        n40558), .C2(n32021), .ZN(n9793) );
  OAI222_X1 U29427 ( .A1(n40805), .A2(n40572), .B1(n41189), .B2(n40565), .C1(
        n40558), .C2(n32020), .ZN(n9792) );
  OAI222_X1 U29428 ( .A1(n40811), .A2(n40572), .B1(n41195), .B2(n40565), .C1(
        n40558), .C2(n32019), .ZN(n9791) );
  OAI222_X1 U29429 ( .A1(n40817), .A2(n40572), .B1(n41201), .B2(n40565), .C1(
        n40559), .C2(n32018), .ZN(n9790) );
  OAI222_X1 U29430 ( .A1(n40823), .A2(n40572), .B1(n41207), .B2(n40565), .C1(
        n40559), .C2(n32017), .ZN(n9789) );
  OAI222_X1 U29431 ( .A1(n40829), .A2(n40572), .B1(n41213), .B2(n40565), .C1(
        n40559), .C2(n32016), .ZN(n9788) );
  OAI222_X1 U29432 ( .A1(n40835), .A2(n40572), .B1(n41219), .B2(n40565), .C1(
        n40559), .C2(n32015), .ZN(n9787) );
  OAI222_X1 U29433 ( .A1(n40841), .A2(n40571), .B1(n41225), .B2(n40564), .C1(
        n40559), .C2(n32014), .ZN(n9786) );
  OAI222_X1 U29434 ( .A1(n40847), .A2(n40571), .B1(n41231), .B2(n40564), .C1(
        n40559), .C2(n32013), .ZN(n9785) );
  OAI222_X1 U29435 ( .A1(n40853), .A2(n40571), .B1(n41237), .B2(n40564), .C1(
        n40559), .C2(n32012), .ZN(n9784) );
  OAI222_X1 U29436 ( .A1(n40859), .A2(n40571), .B1(n41243), .B2(n40564), .C1(
        n40559), .C2(n32011), .ZN(n9783) );
  OAI222_X1 U29437 ( .A1(n40865), .A2(n40571), .B1(n41249), .B2(n40564), .C1(
        n40559), .C2(n32010), .ZN(n9782) );
  OAI222_X1 U29438 ( .A1(n40871), .A2(n40571), .B1(n41255), .B2(n40564), .C1(
        n40559), .C2(n32009), .ZN(n9781) );
  OAI222_X1 U29439 ( .A1(n40877), .A2(n40571), .B1(n41261), .B2(n40564), .C1(
        n40559), .C2(n32008), .ZN(n9780) );
  OAI222_X1 U29440 ( .A1(n40883), .A2(n40571), .B1(n41267), .B2(n40564), .C1(
        n40559), .C2(n32007), .ZN(n9779) );
  OAI222_X1 U29441 ( .A1(n40889), .A2(n40571), .B1(n41273), .B2(n40564), .C1(
        n40560), .C2(n32006), .ZN(n9778) );
  OAI222_X1 U29442 ( .A1(n40895), .A2(n40571), .B1(n41279), .B2(n40564), .C1(
        n40560), .C2(n32005), .ZN(n9777) );
  OAI222_X1 U29443 ( .A1(n40901), .A2(n40571), .B1(n41285), .B2(n40564), .C1(
        n40560), .C2(n32004), .ZN(n9776) );
  OAI222_X1 U29444 ( .A1(n40907), .A2(n40571), .B1(n41291), .B2(n40564), .C1(
        n40560), .C2(n32003), .ZN(n9775) );
  OAI222_X1 U29445 ( .A1(n40913), .A2(n40570), .B1(n41297), .B2(n40563), .C1(
        n40560), .C2(n32002), .ZN(n9774) );
  OAI222_X1 U29446 ( .A1(n40919), .A2(n40570), .B1(n41303), .B2(n40563), .C1(
        n40560), .C2(n32001), .ZN(n9773) );
  OAI222_X1 U29447 ( .A1(n40925), .A2(n40570), .B1(n41309), .B2(n40563), .C1(
        n40560), .C2(n32000), .ZN(n9772) );
  OAI222_X1 U29448 ( .A1(n40931), .A2(n40570), .B1(n41315), .B2(n40563), .C1(
        n40560), .C2(n31999), .ZN(n9771) );
  OAI222_X1 U29449 ( .A1(n40937), .A2(n40570), .B1(n41321), .B2(n40563), .C1(
        n40560), .C2(n31998), .ZN(n9770) );
  OAI222_X1 U29450 ( .A1(n40943), .A2(n40570), .B1(n41327), .B2(n40563), .C1(
        n40560), .C2(n31997), .ZN(n9769) );
  OAI222_X1 U29451 ( .A1(n40949), .A2(n40570), .B1(n41333), .B2(n40563), .C1(
        n40560), .C2(n31996), .ZN(n9768) );
  OAI222_X1 U29452 ( .A1(n40961), .A2(n40570), .B1(n41345), .B2(n40563), .C1(
        n40560), .C2(n31994), .ZN(n9766) );
  OAI222_X1 U29453 ( .A1(n40625), .A2(n40554), .B1(n41009), .B2(n40547), .C1(
        n40536), .C2(n31990), .ZN(n9758) );
  OAI222_X1 U29454 ( .A1(n40631), .A2(n40554), .B1(n41015), .B2(n40547), .C1(
        n40536), .C2(n31989), .ZN(n9757) );
  OAI222_X1 U29455 ( .A1(n40637), .A2(n40554), .B1(n41021), .B2(n40547), .C1(
        n40536), .C2(n31988), .ZN(n9756) );
  OAI222_X1 U29456 ( .A1(n40643), .A2(n40554), .B1(n41027), .B2(n40547), .C1(
        n40536), .C2(n31987), .ZN(n9755) );
  OAI222_X1 U29457 ( .A1(n40649), .A2(n40554), .B1(n41033), .B2(n40547), .C1(
        n40536), .C2(n31986), .ZN(n9754) );
  OAI222_X1 U29458 ( .A1(n40655), .A2(n40554), .B1(n41039), .B2(n40547), .C1(
        n40536), .C2(n31985), .ZN(n9753) );
  OAI222_X1 U29459 ( .A1(n40661), .A2(n40554), .B1(n41045), .B2(n40547), .C1(
        n40536), .C2(n31984), .ZN(n9752) );
  OAI222_X1 U29460 ( .A1(n40667), .A2(n40554), .B1(n41051), .B2(n40547), .C1(
        n40536), .C2(n31983), .ZN(n9751) );
  OAI222_X1 U29461 ( .A1(n40673), .A2(n40554), .B1(n41057), .B2(n40547), .C1(
        n40537), .C2(n31982), .ZN(n9750) );
  OAI222_X1 U29462 ( .A1(n40679), .A2(n40554), .B1(n41063), .B2(n40547), .C1(
        n40537), .C2(n31981), .ZN(n9749) );
  OAI222_X1 U29463 ( .A1(n40685), .A2(n40554), .B1(n41069), .B2(n40547), .C1(
        n40537), .C2(n31980), .ZN(n9748) );
  OAI222_X1 U29464 ( .A1(n40691), .A2(n40554), .B1(n41075), .B2(n40547), .C1(
        n40538), .C2(n31979), .ZN(n9747) );
  OAI222_X1 U29465 ( .A1(n40697), .A2(n40553), .B1(n41081), .B2(n40546), .C1(
        n40537), .C2(n31978), .ZN(n9746) );
  OAI222_X1 U29466 ( .A1(n40703), .A2(n40553), .B1(n41087), .B2(n40546), .C1(
        n40537), .C2(n31977), .ZN(n9745) );
  OAI222_X1 U29467 ( .A1(n40709), .A2(n40553), .B1(n41093), .B2(n40546), .C1(
        n40537), .C2(n31976), .ZN(n9744) );
  OAI222_X1 U29468 ( .A1(n40715), .A2(n40553), .B1(n41099), .B2(n40546), .C1(
        n40537), .C2(n31975), .ZN(n9743) );
  OAI222_X1 U29469 ( .A1(n40721), .A2(n40553), .B1(n41105), .B2(n40546), .C1(
        n40537), .C2(n31974), .ZN(n9742) );
  OAI222_X1 U29470 ( .A1(n40727), .A2(n40553), .B1(n41111), .B2(n40546), .C1(
        n40537), .C2(n31973), .ZN(n9741) );
  OAI222_X1 U29471 ( .A1(n40733), .A2(n40553), .B1(n41117), .B2(n40546), .C1(
        n40537), .C2(n31972), .ZN(n9740) );
  OAI222_X1 U29472 ( .A1(n40739), .A2(n40553), .B1(n41123), .B2(n40546), .C1(
        n40537), .C2(n31971), .ZN(n9739) );
  OAI222_X1 U29473 ( .A1(n40745), .A2(n40553), .B1(n41129), .B2(n40546), .C1(
        n40537), .C2(n31970), .ZN(n9738) );
  OAI222_X1 U29474 ( .A1(n40751), .A2(n40553), .B1(n41135), .B2(n40546), .C1(
        n40538), .C2(n31969), .ZN(n9737) );
  OAI222_X1 U29475 ( .A1(n40757), .A2(n40553), .B1(n41141), .B2(n40546), .C1(
        n40538), .C2(n31968), .ZN(n9736) );
  OAI222_X1 U29476 ( .A1(n40763), .A2(n40553), .B1(n41147), .B2(n40546), .C1(
        n40538), .C2(n31967), .ZN(n9735) );
  OAI222_X1 U29477 ( .A1(n40769), .A2(n40552), .B1(n41153), .B2(n40545), .C1(
        n40538), .C2(n31966), .ZN(n9734) );
  OAI222_X1 U29478 ( .A1(n40775), .A2(n40552), .B1(n41159), .B2(n40545), .C1(
        n40538), .C2(n31965), .ZN(n9733) );
  OAI222_X1 U29479 ( .A1(n40781), .A2(n40552), .B1(n41165), .B2(n40545), .C1(
        n40538), .C2(n31964), .ZN(n9732) );
  OAI222_X1 U29480 ( .A1(n40787), .A2(n40552), .B1(n41171), .B2(n40545), .C1(
        n40538), .C2(n31963), .ZN(n9731) );
  OAI222_X1 U29481 ( .A1(n40793), .A2(n40552), .B1(n41177), .B2(n40545), .C1(
        n40538), .C2(n31962), .ZN(n9730) );
  OAI222_X1 U29482 ( .A1(n40799), .A2(n40552), .B1(n41183), .B2(n40545), .C1(
        n40538), .C2(n31961), .ZN(n9729) );
  OAI222_X1 U29483 ( .A1(n40805), .A2(n40552), .B1(n41189), .B2(n40545), .C1(
        n40538), .C2(n31960), .ZN(n9728) );
  OAI222_X1 U29484 ( .A1(n40811), .A2(n40552), .B1(n41195), .B2(n40545), .C1(
        n40538), .C2(n31959), .ZN(n9727) );
  OAI222_X1 U29485 ( .A1(n40817), .A2(n40552), .B1(n41201), .B2(n40545), .C1(
        n40539), .C2(n31958), .ZN(n9726) );
  OAI222_X1 U29486 ( .A1(n40823), .A2(n40552), .B1(n41207), .B2(n40545), .C1(
        n40539), .C2(n31957), .ZN(n9725) );
  OAI222_X1 U29487 ( .A1(n40829), .A2(n40552), .B1(n41213), .B2(n40545), .C1(
        n40539), .C2(n31956), .ZN(n9724) );
  OAI222_X1 U29488 ( .A1(n40835), .A2(n40552), .B1(n41219), .B2(n40545), .C1(
        n40539), .C2(n31955), .ZN(n9723) );
  OAI222_X1 U29489 ( .A1(n40841), .A2(n40551), .B1(n41225), .B2(n40544), .C1(
        n40539), .C2(n31954), .ZN(n9722) );
  OAI222_X1 U29490 ( .A1(n40847), .A2(n40551), .B1(n41231), .B2(n40544), .C1(
        n40539), .C2(n31953), .ZN(n9721) );
  OAI222_X1 U29491 ( .A1(n40853), .A2(n40551), .B1(n41237), .B2(n40544), .C1(
        n40539), .C2(n31952), .ZN(n9720) );
  OAI222_X1 U29492 ( .A1(n40859), .A2(n40551), .B1(n41243), .B2(n40544), .C1(
        n40539), .C2(n31951), .ZN(n9719) );
  OAI222_X1 U29493 ( .A1(n40865), .A2(n40551), .B1(n41249), .B2(n40544), .C1(
        n40539), .C2(n31950), .ZN(n9718) );
  OAI222_X1 U29494 ( .A1(n40871), .A2(n40551), .B1(n41255), .B2(n40544), .C1(
        n40539), .C2(n31949), .ZN(n9717) );
  OAI222_X1 U29495 ( .A1(n40877), .A2(n40551), .B1(n41261), .B2(n40544), .C1(
        n40539), .C2(n31948), .ZN(n9716) );
  OAI222_X1 U29496 ( .A1(n40883), .A2(n40551), .B1(n41267), .B2(n40544), .C1(
        n40539), .C2(n31947), .ZN(n9715) );
  OAI222_X1 U29497 ( .A1(n40889), .A2(n40551), .B1(n41273), .B2(n40544), .C1(
        n40540), .C2(n31946), .ZN(n9714) );
  OAI222_X1 U29498 ( .A1(n40895), .A2(n40551), .B1(n41279), .B2(n40544), .C1(
        n40540), .C2(n31945), .ZN(n9713) );
  OAI222_X1 U29499 ( .A1(n40901), .A2(n40551), .B1(n41285), .B2(n40544), .C1(
        n40540), .C2(n31944), .ZN(n9712) );
  OAI222_X1 U29500 ( .A1(n40907), .A2(n40551), .B1(n41291), .B2(n40544), .C1(
        n40540), .C2(n31943), .ZN(n9711) );
  OAI222_X1 U29501 ( .A1(n40913), .A2(n40550), .B1(n41297), .B2(n40543), .C1(
        n40540), .C2(n31942), .ZN(n9710) );
  OAI222_X1 U29502 ( .A1(n40919), .A2(n40550), .B1(n41303), .B2(n40543), .C1(
        n40540), .C2(n31941), .ZN(n9709) );
  OAI222_X1 U29503 ( .A1(n40925), .A2(n40550), .B1(n41309), .B2(n40543), .C1(
        n40540), .C2(n31940), .ZN(n9708) );
  OAI222_X1 U29504 ( .A1(n40931), .A2(n40550), .B1(n41315), .B2(n40543), .C1(
        n40540), .C2(n31939), .ZN(n9707) );
  OAI222_X1 U29505 ( .A1(n40937), .A2(n40550), .B1(n41321), .B2(n40543), .C1(
        n40540), .C2(n31938), .ZN(n9706) );
  OAI222_X1 U29506 ( .A1(n40943), .A2(n40550), .B1(n41327), .B2(n40543), .C1(
        n40540), .C2(n31937), .ZN(n9705) );
  OAI222_X1 U29507 ( .A1(n40949), .A2(n40550), .B1(n41333), .B2(n40543), .C1(
        n40540), .C2(n31936), .ZN(n9704) );
  OAI222_X1 U29508 ( .A1(n40961), .A2(n40550), .B1(n41345), .B2(n40543), .C1(
        n40540), .C2(n31934), .ZN(n9702) );
  OAI222_X1 U29509 ( .A1(n40624), .A2(n40494), .B1(n41008), .B2(n40487), .C1(
        n40476), .C2(n31930), .ZN(n9566) );
  OAI222_X1 U29510 ( .A1(n40630), .A2(n40494), .B1(n41014), .B2(n40487), .C1(
        n40476), .C2(n31929), .ZN(n9565) );
  OAI222_X1 U29511 ( .A1(n40636), .A2(n40494), .B1(n41020), .B2(n40487), .C1(
        n40476), .C2(n31928), .ZN(n9564) );
  OAI222_X1 U29512 ( .A1(n40642), .A2(n40494), .B1(n41026), .B2(n40487), .C1(
        n40476), .C2(n31927), .ZN(n9563) );
  OAI222_X1 U29513 ( .A1(n40648), .A2(n40494), .B1(n41032), .B2(n40487), .C1(
        n40476), .C2(n31926), .ZN(n9562) );
  OAI222_X1 U29514 ( .A1(n40654), .A2(n40494), .B1(n41038), .B2(n40487), .C1(
        n40476), .C2(n31925), .ZN(n9561) );
  OAI222_X1 U29515 ( .A1(n40660), .A2(n40494), .B1(n41044), .B2(n40487), .C1(
        n40476), .C2(n31924), .ZN(n9560) );
  OAI222_X1 U29516 ( .A1(n40666), .A2(n40494), .B1(n41050), .B2(n40487), .C1(
        n40476), .C2(n31923), .ZN(n9559) );
  OAI222_X1 U29517 ( .A1(n40672), .A2(n40494), .B1(n41056), .B2(n40487), .C1(
        n40477), .C2(n31922), .ZN(n9558) );
  OAI222_X1 U29518 ( .A1(n40678), .A2(n40494), .B1(n41062), .B2(n40487), .C1(
        n40477), .C2(n31921), .ZN(n9557) );
  OAI222_X1 U29519 ( .A1(n40684), .A2(n40494), .B1(n41068), .B2(n40487), .C1(
        n40477), .C2(n31920), .ZN(n9556) );
  OAI222_X1 U29520 ( .A1(n40690), .A2(n40494), .B1(n41074), .B2(n40487), .C1(
        n40478), .C2(n31919), .ZN(n9555) );
  OAI222_X1 U29521 ( .A1(n40696), .A2(n40493), .B1(n41080), .B2(n40486), .C1(
        n40477), .C2(n31918), .ZN(n9554) );
  OAI222_X1 U29522 ( .A1(n40702), .A2(n40493), .B1(n41086), .B2(n40486), .C1(
        n40477), .C2(n31917), .ZN(n9553) );
  OAI222_X1 U29523 ( .A1(n40708), .A2(n40493), .B1(n41092), .B2(n40486), .C1(
        n40477), .C2(n31916), .ZN(n9552) );
  OAI222_X1 U29524 ( .A1(n40714), .A2(n40493), .B1(n41098), .B2(n40486), .C1(
        n40477), .C2(n31915), .ZN(n9551) );
  OAI222_X1 U29525 ( .A1(n40720), .A2(n40493), .B1(n41104), .B2(n40486), .C1(
        n40477), .C2(n31914), .ZN(n9550) );
  OAI222_X1 U29526 ( .A1(n40726), .A2(n40493), .B1(n41110), .B2(n40486), .C1(
        n40477), .C2(n31913), .ZN(n9549) );
  OAI222_X1 U29527 ( .A1(n40732), .A2(n40493), .B1(n41116), .B2(n40486), .C1(
        n40477), .C2(n31912), .ZN(n9548) );
  OAI222_X1 U29528 ( .A1(n40738), .A2(n40493), .B1(n41122), .B2(n40486), .C1(
        n40477), .C2(n31911), .ZN(n9547) );
  OAI222_X1 U29529 ( .A1(n40744), .A2(n40493), .B1(n41128), .B2(n40486), .C1(
        n40477), .C2(n31910), .ZN(n9546) );
  OAI222_X1 U29530 ( .A1(n40750), .A2(n40493), .B1(n41134), .B2(n40486), .C1(
        n40478), .C2(n31909), .ZN(n9545) );
  OAI222_X1 U29531 ( .A1(n40756), .A2(n40493), .B1(n41140), .B2(n40486), .C1(
        n40478), .C2(n31908), .ZN(n9544) );
  OAI222_X1 U29532 ( .A1(n40762), .A2(n40493), .B1(n41146), .B2(n40486), .C1(
        n40478), .C2(n31907), .ZN(n9543) );
  OAI222_X1 U29533 ( .A1(n40768), .A2(n40492), .B1(n41152), .B2(n40485), .C1(
        n40478), .C2(n31906), .ZN(n9542) );
  OAI222_X1 U29534 ( .A1(n40774), .A2(n40492), .B1(n41158), .B2(n40485), .C1(
        n40478), .C2(n31905), .ZN(n9541) );
  OAI222_X1 U29535 ( .A1(n40780), .A2(n40492), .B1(n41164), .B2(n40485), .C1(
        n40478), .C2(n31904), .ZN(n9540) );
  OAI222_X1 U29536 ( .A1(n40786), .A2(n40492), .B1(n41170), .B2(n40485), .C1(
        n40478), .C2(n31903), .ZN(n9539) );
  OAI222_X1 U29537 ( .A1(n40792), .A2(n40492), .B1(n41176), .B2(n40485), .C1(
        n40478), .C2(n31902), .ZN(n9538) );
  OAI222_X1 U29538 ( .A1(n40798), .A2(n40492), .B1(n41182), .B2(n40485), .C1(
        n40478), .C2(n31901), .ZN(n9537) );
  OAI222_X1 U29539 ( .A1(n40804), .A2(n40492), .B1(n41188), .B2(n40485), .C1(
        n40478), .C2(n31900), .ZN(n9536) );
  OAI222_X1 U29540 ( .A1(n40810), .A2(n40492), .B1(n41194), .B2(n40485), .C1(
        n40478), .C2(n31899), .ZN(n9535) );
  OAI222_X1 U29541 ( .A1(n40816), .A2(n40492), .B1(n41200), .B2(n40485), .C1(
        n40479), .C2(n31898), .ZN(n9534) );
  OAI222_X1 U29542 ( .A1(n40822), .A2(n40492), .B1(n41206), .B2(n40485), .C1(
        n40479), .C2(n31897), .ZN(n9533) );
  OAI222_X1 U29543 ( .A1(n40828), .A2(n40492), .B1(n41212), .B2(n40485), .C1(
        n40479), .C2(n31896), .ZN(n9532) );
  OAI222_X1 U29544 ( .A1(n40834), .A2(n40492), .B1(n41218), .B2(n40485), .C1(
        n40479), .C2(n31895), .ZN(n9531) );
  OAI222_X1 U29545 ( .A1(n40840), .A2(n40491), .B1(n41224), .B2(n40484), .C1(
        n40479), .C2(n31894), .ZN(n9530) );
  OAI222_X1 U29546 ( .A1(n40846), .A2(n40491), .B1(n41230), .B2(n40484), .C1(
        n40479), .C2(n31893), .ZN(n9529) );
  OAI222_X1 U29547 ( .A1(n40852), .A2(n40491), .B1(n41236), .B2(n40484), .C1(
        n40479), .C2(n31892), .ZN(n9528) );
  OAI222_X1 U29548 ( .A1(n40858), .A2(n40491), .B1(n41242), .B2(n40484), .C1(
        n40479), .C2(n31891), .ZN(n9527) );
  OAI222_X1 U29549 ( .A1(n40864), .A2(n40491), .B1(n41248), .B2(n40484), .C1(
        n40479), .C2(n31890), .ZN(n9526) );
  OAI222_X1 U29550 ( .A1(n40870), .A2(n40491), .B1(n41254), .B2(n40484), .C1(
        n40479), .C2(n31889), .ZN(n9525) );
  OAI222_X1 U29551 ( .A1(n40876), .A2(n40491), .B1(n41260), .B2(n40484), .C1(
        n40479), .C2(n31888), .ZN(n9524) );
  OAI222_X1 U29552 ( .A1(n40882), .A2(n40491), .B1(n41266), .B2(n40484), .C1(
        n40479), .C2(n31887), .ZN(n9523) );
  OAI222_X1 U29553 ( .A1(n40888), .A2(n40491), .B1(n41272), .B2(n40484), .C1(
        n40480), .C2(n31886), .ZN(n9522) );
  OAI222_X1 U29554 ( .A1(n40894), .A2(n40491), .B1(n41278), .B2(n40484), .C1(
        n40480), .C2(n31885), .ZN(n9521) );
  OAI222_X1 U29555 ( .A1(n40900), .A2(n40491), .B1(n41284), .B2(n40484), .C1(
        n40480), .C2(n31884), .ZN(n9520) );
  OAI222_X1 U29556 ( .A1(n40906), .A2(n40491), .B1(n41290), .B2(n40484), .C1(
        n40480), .C2(n31883), .ZN(n9519) );
  OAI222_X1 U29557 ( .A1(n40912), .A2(n40490), .B1(n41296), .B2(n40483), .C1(
        n40480), .C2(n31882), .ZN(n9518) );
  OAI222_X1 U29558 ( .A1(n40918), .A2(n40490), .B1(n41302), .B2(n40483), .C1(
        n40480), .C2(n31881), .ZN(n9517) );
  OAI222_X1 U29559 ( .A1(n40924), .A2(n40490), .B1(n41308), .B2(n40483), .C1(
        n40480), .C2(n31880), .ZN(n9516) );
  OAI222_X1 U29560 ( .A1(n40930), .A2(n40490), .B1(n41314), .B2(n40483), .C1(
        n40480), .C2(n31879), .ZN(n9515) );
  OAI222_X1 U29561 ( .A1(n40936), .A2(n40490), .B1(n41320), .B2(n40483), .C1(
        n40480), .C2(n31878), .ZN(n9514) );
  OAI222_X1 U29562 ( .A1(n40942), .A2(n40490), .B1(n41326), .B2(n40483), .C1(
        n40480), .C2(n31877), .ZN(n9513) );
  OAI222_X1 U29563 ( .A1(n40948), .A2(n40490), .B1(n41332), .B2(n40483), .C1(
        n40480), .C2(n31876), .ZN(n9512) );
  OAI222_X1 U29564 ( .A1(n40960), .A2(n40490), .B1(n41344), .B2(n40483), .C1(
        n40480), .C2(n31874), .ZN(n9510) );
  OAI222_X1 U29565 ( .A1(n40624), .A2(n40474), .B1(n41008), .B2(n40467), .C1(
        n40456), .C2(n31870), .ZN(n9502) );
  OAI222_X1 U29566 ( .A1(n40630), .A2(n40474), .B1(n41014), .B2(n40467), .C1(
        n40456), .C2(n31869), .ZN(n9501) );
  OAI222_X1 U29567 ( .A1(n40636), .A2(n40474), .B1(n41020), .B2(n40467), .C1(
        n40456), .C2(n31868), .ZN(n9500) );
  OAI222_X1 U29568 ( .A1(n40642), .A2(n40474), .B1(n41026), .B2(n40467), .C1(
        n40456), .C2(n31867), .ZN(n9499) );
  OAI222_X1 U29569 ( .A1(n40648), .A2(n40474), .B1(n41032), .B2(n40467), .C1(
        n40456), .C2(n31866), .ZN(n9498) );
  OAI222_X1 U29570 ( .A1(n40654), .A2(n40474), .B1(n41038), .B2(n40467), .C1(
        n40456), .C2(n31865), .ZN(n9497) );
  OAI222_X1 U29571 ( .A1(n40660), .A2(n40474), .B1(n41044), .B2(n40467), .C1(
        n40456), .C2(n31864), .ZN(n9496) );
  OAI222_X1 U29572 ( .A1(n40666), .A2(n40474), .B1(n41050), .B2(n40467), .C1(
        n40456), .C2(n31863), .ZN(n9495) );
  OAI222_X1 U29573 ( .A1(n40672), .A2(n40474), .B1(n41056), .B2(n40467), .C1(
        n40457), .C2(n31862), .ZN(n9494) );
  OAI222_X1 U29574 ( .A1(n40678), .A2(n40474), .B1(n41062), .B2(n40467), .C1(
        n40457), .C2(n31861), .ZN(n9493) );
  OAI222_X1 U29575 ( .A1(n40684), .A2(n40474), .B1(n41068), .B2(n40467), .C1(
        n40457), .C2(n31860), .ZN(n9492) );
  OAI222_X1 U29576 ( .A1(n40690), .A2(n40474), .B1(n41074), .B2(n40467), .C1(
        n40458), .C2(n31859), .ZN(n9491) );
  OAI222_X1 U29577 ( .A1(n40696), .A2(n40473), .B1(n41080), .B2(n40466), .C1(
        n40457), .C2(n31858), .ZN(n9490) );
  OAI222_X1 U29578 ( .A1(n40702), .A2(n40473), .B1(n41086), .B2(n40466), .C1(
        n40457), .C2(n31857), .ZN(n9489) );
  OAI222_X1 U29579 ( .A1(n40708), .A2(n40473), .B1(n41092), .B2(n40466), .C1(
        n40457), .C2(n31856), .ZN(n9488) );
  OAI222_X1 U29580 ( .A1(n40714), .A2(n40473), .B1(n41098), .B2(n40466), .C1(
        n40457), .C2(n31855), .ZN(n9487) );
  OAI222_X1 U29581 ( .A1(n40720), .A2(n40473), .B1(n41104), .B2(n40466), .C1(
        n40457), .C2(n31854), .ZN(n9486) );
  OAI222_X1 U29582 ( .A1(n40726), .A2(n40473), .B1(n41110), .B2(n40466), .C1(
        n40457), .C2(n31853), .ZN(n9485) );
  OAI222_X1 U29583 ( .A1(n40732), .A2(n40473), .B1(n41116), .B2(n40466), .C1(
        n40457), .C2(n31852), .ZN(n9484) );
  OAI222_X1 U29584 ( .A1(n40738), .A2(n40473), .B1(n41122), .B2(n40466), .C1(
        n40457), .C2(n31851), .ZN(n9483) );
  OAI222_X1 U29585 ( .A1(n40744), .A2(n40473), .B1(n41128), .B2(n40466), .C1(
        n40457), .C2(n31850), .ZN(n9482) );
  OAI222_X1 U29586 ( .A1(n40750), .A2(n40473), .B1(n41134), .B2(n40466), .C1(
        n40458), .C2(n31849), .ZN(n9481) );
  OAI222_X1 U29587 ( .A1(n40756), .A2(n40473), .B1(n41140), .B2(n40466), .C1(
        n40458), .C2(n31848), .ZN(n9480) );
  OAI222_X1 U29588 ( .A1(n40762), .A2(n40473), .B1(n41146), .B2(n40466), .C1(
        n40458), .C2(n31847), .ZN(n9479) );
  OAI222_X1 U29589 ( .A1(n40768), .A2(n40472), .B1(n41152), .B2(n40465), .C1(
        n40458), .C2(n31846), .ZN(n9478) );
  OAI222_X1 U29590 ( .A1(n40774), .A2(n40472), .B1(n41158), .B2(n40465), .C1(
        n40458), .C2(n31845), .ZN(n9477) );
  OAI222_X1 U29591 ( .A1(n40780), .A2(n40472), .B1(n41164), .B2(n40465), .C1(
        n40458), .C2(n31844), .ZN(n9476) );
  OAI222_X1 U29592 ( .A1(n40786), .A2(n40472), .B1(n41170), .B2(n40465), .C1(
        n40458), .C2(n31843), .ZN(n9475) );
  OAI222_X1 U29593 ( .A1(n40792), .A2(n40472), .B1(n41176), .B2(n40465), .C1(
        n40458), .C2(n31842), .ZN(n9474) );
  OAI222_X1 U29594 ( .A1(n40798), .A2(n40472), .B1(n41182), .B2(n40465), .C1(
        n40458), .C2(n31841), .ZN(n9473) );
  OAI222_X1 U29595 ( .A1(n40804), .A2(n40472), .B1(n41188), .B2(n40465), .C1(
        n40458), .C2(n31840), .ZN(n9472) );
  OAI222_X1 U29596 ( .A1(n40810), .A2(n40472), .B1(n41194), .B2(n40465), .C1(
        n40458), .C2(n31839), .ZN(n9471) );
  OAI222_X1 U29597 ( .A1(n40816), .A2(n40472), .B1(n41200), .B2(n40465), .C1(
        n40459), .C2(n31838), .ZN(n9470) );
  OAI222_X1 U29598 ( .A1(n40822), .A2(n40472), .B1(n41206), .B2(n40465), .C1(
        n40459), .C2(n31837), .ZN(n9469) );
  OAI222_X1 U29599 ( .A1(n40828), .A2(n40472), .B1(n41212), .B2(n40465), .C1(
        n40459), .C2(n31836), .ZN(n9468) );
  OAI222_X1 U29600 ( .A1(n40834), .A2(n40472), .B1(n41218), .B2(n40465), .C1(
        n40459), .C2(n31835), .ZN(n9467) );
  OAI222_X1 U29601 ( .A1(n40840), .A2(n40471), .B1(n41224), .B2(n40464), .C1(
        n40459), .C2(n31834), .ZN(n9466) );
  OAI222_X1 U29602 ( .A1(n40846), .A2(n40471), .B1(n41230), .B2(n40464), .C1(
        n40459), .C2(n31833), .ZN(n9465) );
  OAI222_X1 U29603 ( .A1(n40852), .A2(n40471), .B1(n41236), .B2(n40464), .C1(
        n40459), .C2(n31832), .ZN(n9464) );
  OAI222_X1 U29604 ( .A1(n40858), .A2(n40471), .B1(n41242), .B2(n40464), .C1(
        n40459), .C2(n31831), .ZN(n9463) );
  OAI222_X1 U29605 ( .A1(n40864), .A2(n40471), .B1(n41248), .B2(n40464), .C1(
        n40459), .C2(n31830), .ZN(n9462) );
  OAI222_X1 U29606 ( .A1(n40870), .A2(n40471), .B1(n41254), .B2(n40464), .C1(
        n40459), .C2(n31829), .ZN(n9461) );
  OAI222_X1 U29607 ( .A1(n40876), .A2(n40471), .B1(n41260), .B2(n40464), .C1(
        n40459), .C2(n31828), .ZN(n9460) );
  OAI222_X1 U29608 ( .A1(n40882), .A2(n40471), .B1(n41266), .B2(n40464), .C1(
        n40459), .C2(n31827), .ZN(n9459) );
  OAI222_X1 U29609 ( .A1(n40888), .A2(n40471), .B1(n41272), .B2(n40464), .C1(
        n40460), .C2(n31826), .ZN(n9458) );
  OAI222_X1 U29610 ( .A1(n40894), .A2(n40471), .B1(n41278), .B2(n40464), .C1(
        n40460), .C2(n31825), .ZN(n9457) );
  OAI222_X1 U29611 ( .A1(n40900), .A2(n40471), .B1(n41284), .B2(n40464), .C1(
        n40460), .C2(n31824), .ZN(n9456) );
  OAI222_X1 U29612 ( .A1(n40906), .A2(n40471), .B1(n41290), .B2(n40464), .C1(
        n40460), .C2(n31823), .ZN(n9455) );
  OAI222_X1 U29613 ( .A1(n40912), .A2(n40470), .B1(n41296), .B2(n40463), .C1(
        n40460), .C2(n31822), .ZN(n9454) );
  OAI222_X1 U29614 ( .A1(n40918), .A2(n40470), .B1(n41302), .B2(n40463), .C1(
        n40460), .C2(n31821), .ZN(n9453) );
  OAI222_X1 U29615 ( .A1(n40924), .A2(n40470), .B1(n41308), .B2(n40463), .C1(
        n40460), .C2(n31820), .ZN(n9452) );
  OAI222_X1 U29616 ( .A1(n40930), .A2(n40470), .B1(n41314), .B2(n40463), .C1(
        n40460), .C2(n31819), .ZN(n9451) );
  OAI222_X1 U29617 ( .A1(n40936), .A2(n40470), .B1(n41320), .B2(n40463), .C1(
        n40460), .C2(n31818), .ZN(n9450) );
  OAI222_X1 U29618 ( .A1(n40942), .A2(n40470), .B1(n41326), .B2(n40463), .C1(
        n40460), .C2(n31817), .ZN(n9449) );
  OAI222_X1 U29619 ( .A1(n40948), .A2(n40470), .B1(n41332), .B2(n40463), .C1(
        n40460), .C2(n31816), .ZN(n9448) );
  OAI222_X1 U29620 ( .A1(n40960), .A2(n40470), .B1(n41344), .B2(n40463), .C1(
        n40460), .C2(n31814), .ZN(n9446) );
  OAI222_X1 U29621 ( .A1(n40624), .A2(n40454), .B1(n41008), .B2(n40447), .C1(
        n40436), .C2(n31810), .ZN(n9438) );
  OAI222_X1 U29622 ( .A1(n40630), .A2(n40454), .B1(n41014), .B2(n40447), .C1(
        n40436), .C2(n31809), .ZN(n9437) );
  OAI222_X1 U29623 ( .A1(n40636), .A2(n40454), .B1(n41020), .B2(n40447), .C1(
        n40436), .C2(n31808), .ZN(n9436) );
  OAI222_X1 U29624 ( .A1(n40642), .A2(n40454), .B1(n41026), .B2(n40447), .C1(
        n40436), .C2(n31807), .ZN(n9435) );
  OAI222_X1 U29625 ( .A1(n40648), .A2(n40454), .B1(n41032), .B2(n40447), .C1(
        n40436), .C2(n31806), .ZN(n9434) );
  OAI222_X1 U29626 ( .A1(n40654), .A2(n40454), .B1(n41038), .B2(n40447), .C1(
        n40436), .C2(n31805), .ZN(n9433) );
  OAI222_X1 U29627 ( .A1(n40660), .A2(n40454), .B1(n41044), .B2(n40447), .C1(
        n40436), .C2(n31804), .ZN(n9432) );
  OAI222_X1 U29628 ( .A1(n40666), .A2(n40454), .B1(n41050), .B2(n40447), .C1(
        n40436), .C2(n31803), .ZN(n9431) );
  OAI222_X1 U29629 ( .A1(n40672), .A2(n40454), .B1(n41056), .B2(n40447), .C1(
        n40437), .C2(n31802), .ZN(n9430) );
  OAI222_X1 U29630 ( .A1(n40678), .A2(n40454), .B1(n41062), .B2(n40447), .C1(
        n40437), .C2(n31801), .ZN(n9429) );
  OAI222_X1 U29631 ( .A1(n40684), .A2(n40454), .B1(n41068), .B2(n40447), .C1(
        n40437), .C2(n31800), .ZN(n9428) );
  OAI222_X1 U29632 ( .A1(n40690), .A2(n40454), .B1(n41074), .B2(n40447), .C1(
        n40438), .C2(n31799), .ZN(n9427) );
  OAI222_X1 U29633 ( .A1(n40696), .A2(n40453), .B1(n41080), .B2(n40446), .C1(
        n40437), .C2(n31798), .ZN(n9426) );
  OAI222_X1 U29634 ( .A1(n40702), .A2(n40453), .B1(n41086), .B2(n40446), .C1(
        n40437), .C2(n31797), .ZN(n9425) );
  OAI222_X1 U29635 ( .A1(n40708), .A2(n40453), .B1(n41092), .B2(n40446), .C1(
        n40437), .C2(n31796), .ZN(n9424) );
  OAI222_X1 U29636 ( .A1(n40714), .A2(n40453), .B1(n41098), .B2(n40446), .C1(
        n40437), .C2(n31795), .ZN(n9423) );
  OAI222_X1 U29637 ( .A1(n40720), .A2(n40453), .B1(n41104), .B2(n40446), .C1(
        n40437), .C2(n31794), .ZN(n9422) );
  OAI222_X1 U29638 ( .A1(n40726), .A2(n40453), .B1(n41110), .B2(n40446), .C1(
        n40437), .C2(n31793), .ZN(n9421) );
  OAI222_X1 U29639 ( .A1(n40732), .A2(n40453), .B1(n41116), .B2(n40446), .C1(
        n40437), .C2(n31792), .ZN(n9420) );
  OAI222_X1 U29640 ( .A1(n40738), .A2(n40453), .B1(n41122), .B2(n40446), .C1(
        n40437), .C2(n31791), .ZN(n9419) );
  OAI222_X1 U29641 ( .A1(n40744), .A2(n40453), .B1(n41128), .B2(n40446), .C1(
        n40437), .C2(n31790), .ZN(n9418) );
  OAI222_X1 U29642 ( .A1(n40750), .A2(n40453), .B1(n41134), .B2(n40446), .C1(
        n40438), .C2(n31789), .ZN(n9417) );
  OAI222_X1 U29643 ( .A1(n40756), .A2(n40453), .B1(n41140), .B2(n40446), .C1(
        n40438), .C2(n31788), .ZN(n9416) );
  OAI222_X1 U29644 ( .A1(n40762), .A2(n40453), .B1(n41146), .B2(n40446), .C1(
        n40438), .C2(n31787), .ZN(n9415) );
  OAI222_X1 U29645 ( .A1(n40768), .A2(n40452), .B1(n41152), .B2(n40445), .C1(
        n40438), .C2(n31786), .ZN(n9414) );
  OAI222_X1 U29646 ( .A1(n40774), .A2(n40452), .B1(n41158), .B2(n40445), .C1(
        n40438), .C2(n31785), .ZN(n9413) );
  OAI222_X1 U29647 ( .A1(n40780), .A2(n40452), .B1(n41164), .B2(n40445), .C1(
        n40438), .C2(n31784), .ZN(n9412) );
  OAI222_X1 U29648 ( .A1(n40786), .A2(n40452), .B1(n41170), .B2(n40445), .C1(
        n40438), .C2(n31783), .ZN(n9411) );
  OAI222_X1 U29649 ( .A1(n40792), .A2(n40452), .B1(n41176), .B2(n40445), .C1(
        n40438), .C2(n31782), .ZN(n9410) );
  OAI222_X1 U29650 ( .A1(n40798), .A2(n40452), .B1(n41182), .B2(n40445), .C1(
        n40438), .C2(n31781), .ZN(n9409) );
  OAI222_X1 U29651 ( .A1(n40804), .A2(n40452), .B1(n41188), .B2(n40445), .C1(
        n40438), .C2(n31780), .ZN(n9408) );
  OAI222_X1 U29652 ( .A1(n40810), .A2(n40452), .B1(n41194), .B2(n40445), .C1(
        n40438), .C2(n31779), .ZN(n9407) );
  OAI222_X1 U29653 ( .A1(n40816), .A2(n40452), .B1(n41200), .B2(n40445), .C1(
        n40439), .C2(n31778), .ZN(n9406) );
  OAI222_X1 U29654 ( .A1(n40822), .A2(n40452), .B1(n41206), .B2(n40445), .C1(
        n40439), .C2(n31777), .ZN(n9405) );
  OAI222_X1 U29655 ( .A1(n40828), .A2(n40452), .B1(n41212), .B2(n40445), .C1(
        n40439), .C2(n31776), .ZN(n9404) );
  OAI222_X1 U29656 ( .A1(n40834), .A2(n40452), .B1(n41218), .B2(n40445), .C1(
        n40439), .C2(n31775), .ZN(n9403) );
  OAI222_X1 U29657 ( .A1(n40840), .A2(n40451), .B1(n41224), .B2(n40444), .C1(
        n40439), .C2(n31774), .ZN(n9402) );
  OAI222_X1 U29658 ( .A1(n40846), .A2(n40451), .B1(n41230), .B2(n40444), .C1(
        n40439), .C2(n31773), .ZN(n9401) );
  OAI222_X1 U29659 ( .A1(n40852), .A2(n40451), .B1(n41236), .B2(n40444), .C1(
        n40439), .C2(n31772), .ZN(n9400) );
  OAI222_X1 U29660 ( .A1(n40858), .A2(n40451), .B1(n41242), .B2(n40444), .C1(
        n40439), .C2(n31771), .ZN(n9399) );
  OAI222_X1 U29661 ( .A1(n40864), .A2(n40451), .B1(n41248), .B2(n40444), .C1(
        n40439), .C2(n31770), .ZN(n9398) );
  OAI222_X1 U29662 ( .A1(n40870), .A2(n40451), .B1(n41254), .B2(n40444), .C1(
        n40439), .C2(n31769), .ZN(n9397) );
  OAI222_X1 U29663 ( .A1(n40876), .A2(n40451), .B1(n41260), .B2(n40444), .C1(
        n40439), .C2(n31768), .ZN(n9396) );
  OAI222_X1 U29664 ( .A1(n40882), .A2(n40451), .B1(n41266), .B2(n40444), .C1(
        n40439), .C2(n31767), .ZN(n9395) );
  OAI222_X1 U29665 ( .A1(n40888), .A2(n40451), .B1(n41272), .B2(n40444), .C1(
        n40440), .C2(n31766), .ZN(n9394) );
  OAI222_X1 U29666 ( .A1(n40894), .A2(n40451), .B1(n41278), .B2(n40444), .C1(
        n40440), .C2(n31765), .ZN(n9393) );
  OAI222_X1 U29667 ( .A1(n40900), .A2(n40451), .B1(n41284), .B2(n40444), .C1(
        n40440), .C2(n31764), .ZN(n9392) );
  OAI222_X1 U29668 ( .A1(n40906), .A2(n40451), .B1(n41290), .B2(n40444), .C1(
        n40440), .C2(n31763), .ZN(n9391) );
  OAI222_X1 U29669 ( .A1(n40912), .A2(n40450), .B1(n41296), .B2(n40443), .C1(
        n40440), .C2(n31762), .ZN(n9390) );
  OAI222_X1 U29670 ( .A1(n40918), .A2(n40450), .B1(n41302), .B2(n40443), .C1(
        n40440), .C2(n31761), .ZN(n9389) );
  OAI222_X1 U29671 ( .A1(n40924), .A2(n40450), .B1(n41308), .B2(n40443), .C1(
        n40440), .C2(n31760), .ZN(n9388) );
  OAI222_X1 U29672 ( .A1(n40930), .A2(n40450), .B1(n41314), .B2(n40443), .C1(
        n40440), .C2(n31759), .ZN(n9387) );
  OAI222_X1 U29673 ( .A1(n40936), .A2(n40450), .B1(n41320), .B2(n40443), .C1(
        n40440), .C2(n31758), .ZN(n9386) );
  OAI222_X1 U29674 ( .A1(n40942), .A2(n40450), .B1(n41326), .B2(n40443), .C1(
        n40440), .C2(n31757), .ZN(n9385) );
  OAI222_X1 U29675 ( .A1(n40948), .A2(n40450), .B1(n41332), .B2(n40443), .C1(
        n40440), .C2(n31756), .ZN(n9384) );
  OAI222_X1 U29676 ( .A1(n40960), .A2(n40450), .B1(n41344), .B2(n40443), .C1(
        n40440), .C2(n31754), .ZN(n9382) );
  OAI222_X1 U29677 ( .A1(n40600), .A2(n40395), .B1(n40984), .B2(n40388), .C1(
        n40376), .C2(n31750), .ZN(n9250) );
  OAI222_X1 U29678 ( .A1(n40606), .A2(n40395), .B1(n40990), .B2(n40388), .C1(
        n40376), .C2(n31749), .ZN(n9249) );
  OAI222_X1 U29679 ( .A1(n40612), .A2(n40395), .B1(n40996), .B2(n40388), .C1(
        n40376), .C2(n31748), .ZN(n9248) );
  OAI222_X1 U29680 ( .A1(n40618), .A2(n40395), .B1(n41002), .B2(n40388), .C1(
        n40376), .C2(n31747), .ZN(n9247) );
  OAI222_X1 U29681 ( .A1(n40624), .A2(n40394), .B1(n41008), .B2(n40387), .C1(
        n40376), .C2(n31746), .ZN(n9246) );
  OAI222_X1 U29682 ( .A1(n40630), .A2(n40394), .B1(n41014), .B2(n40387), .C1(
        n40376), .C2(n31745), .ZN(n9245) );
  OAI222_X1 U29683 ( .A1(n40636), .A2(n40394), .B1(n41020), .B2(n40387), .C1(
        n40376), .C2(n31744), .ZN(n9244) );
  OAI222_X1 U29684 ( .A1(n40642), .A2(n40394), .B1(n41026), .B2(n40387), .C1(
        n40376), .C2(n31743), .ZN(n9243) );
  OAI222_X1 U29685 ( .A1(n40648), .A2(n40394), .B1(n41032), .B2(n40387), .C1(
        n40376), .C2(n31742), .ZN(n9242) );
  OAI222_X1 U29686 ( .A1(n40654), .A2(n40394), .B1(n41038), .B2(n40387), .C1(
        n40376), .C2(n31741), .ZN(n9241) );
  OAI222_X1 U29687 ( .A1(n40660), .A2(n40394), .B1(n41044), .B2(n40387), .C1(
        n40376), .C2(n31740), .ZN(n9240) );
  OAI222_X1 U29688 ( .A1(n40666), .A2(n40394), .B1(n41050), .B2(n40387), .C1(
        n40376), .C2(n31739), .ZN(n9239) );
  OAI222_X1 U29689 ( .A1(n40672), .A2(n40394), .B1(n41056), .B2(n40387), .C1(
        n40377), .C2(n31738), .ZN(n9238) );
  OAI222_X1 U29690 ( .A1(n40678), .A2(n40394), .B1(n41062), .B2(n40387), .C1(
        n40377), .C2(n31737), .ZN(n9237) );
  OAI222_X1 U29691 ( .A1(n40684), .A2(n40394), .B1(n41068), .B2(n40387), .C1(
        n40377), .C2(n31736), .ZN(n9236) );
  OAI222_X1 U29692 ( .A1(n40690), .A2(n40394), .B1(n41074), .B2(n40387), .C1(
        n40378), .C2(n31735), .ZN(n9235) );
  OAI222_X1 U29693 ( .A1(n40696), .A2(n40393), .B1(n41080), .B2(n40386), .C1(
        n40377), .C2(n31734), .ZN(n9234) );
  OAI222_X1 U29694 ( .A1(n40702), .A2(n40393), .B1(n41086), .B2(n40386), .C1(
        n40377), .C2(n31733), .ZN(n9233) );
  OAI222_X1 U29695 ( .A1(n40708), .A2(n40393), .B1(n41092), .B2(n40386), .C1(
        n40377), .C2(n31732), .ZN(n9232) );
  OAI222_X1 U29696 ( .A1(n40714), .A2(n40393), .B1(n41098), .B2(n40386), .C1(
        n40377), .C2(n31731), .ZN(n9231) );
  OAI222_X1 U29697 ( .A1(n40720), .A2(n40393), .B1(n41104), .B2(n40386), .C1(
        n40377), .C2(n31730), .ZN(n9230) );
  OAI222_X1 U29698 ( .A1(n40726), .A2(n40393), .B1(n41110), .B2(n40386), .C1(
        n40377), .C2(n31729), .ZN(n9229) );
  OAI222_X1 U29699 ( .A1(n40732), .A2(n40393), .B1(n41116), .B2(n40386), .C1(
        n40377), .C2(n31728), .ZN(n9228) );
  OAI222_X1 U29700 ( .A1(n40738), .A2(n40393), .B1(n41122), .B2(n40386), .C1(
        n40377), .C2(n31727), .ZN(n9227) );
  OAI222_X1 U29701 ( .A1(n40744), .A2(n40393), .B1(n41128), .B2(n40386), .C1(
        n40377), .C2(n31726), .ZN(n9226) );
  OAI222_X1 U29702 ( .A1(n40750), .A2(n40393), .B1(n41134), .B2(n40386), .C1(
        n40378), .C2(n31725), .ZN(n9225) );
  OAI222_X1 U29703 ( .A1(n40756), .A2(n40393), .B1(n41140), .B2(n40386), .C1(
        n40378), .C2(n31724), .ZN(n9224) );
  OAI222_X1 U29704 ( .A1(n40762), .A2(n40393), .B1(n41146), .B2(n40386), .C1(
        n40378), .C2(n31723), .ZN(n9223) );
  OAI222_X1 U29705 ( .A1(n40768), .A2(n40392), .B1(n41152), .B2(n40385), .C1(
        n40378), .C2(n31722), .ZN(n9222) );
  OAI222_X1 U29706 ( .A1(n40774), .A2(n40392), .B1(n41158), .B2(n40385), .C1(
        n40378), .C2(n31721), .ZN(n9221) );
  OAI222_X1 U29707 ( .A1(n40780), .A2(n40392), .B1(n41164), .B2(n40385), .C1(
        n40378), .C2(n31720), .ZN(n9220) );
  OAI222_X1 U29708 ( .A1(n40786), .A2(n40392), .B1(n41170), .B2(n40385), .C1(
        n40378), .C2(n31719), .ZN(n9219) );
  OAI222_X1 U29709 ( .A1(n40792), .A2(n40392), .B1(n41176), .B2(n40385), .C1(
        n40378), .C2(n31718), .ZN(n9218) );
  OAI222_X1 U29710 ( .A1(n40798), .A2(n40392), .B1(n41182), .B2(n40385), .C1(
        n40378), .C2(n31717), .ZN(n9217) );
  OAI222_X1 U29711 ( .A1(n40804), .A2(n40392), .B1(n41188), .B2(n40385), .C1(
        n40378), .C2(n31716), .ZN(n9216) );
  OAI222_X1 U29712 ( .A1(n40810), .A2(n40392), .B1(n41194), .B2(n40385), .C1(
        n40378), .C2(n31715), .ZN(n9215) );
  OAI222_X1 U29713 ( .A1(n40816), .A2(n40392), .B1(n41200), .B2(n40385), .C1(
        n40379), .C2(n31714), .ZN(n9214) );
  OAI222_X1 U29714 ( .A1(n40822), .A2(n40392), .B1(n41206), .B2(n40385), .C1(
        n40379), .C2(n31713), .ZN(n9213) );
  OAI222_X1 U29715 ( .A1(n40828), .A2(n40392), .B1(n41212), .B2(n40385), .C1(
        n40379), .C2(n31712), .ZN(n9212) );
  OAI222_X1 U29716 ( .A1(n40834), .A2(n40392), .B1(n41218), .B2(n40385), .C1(
        n40379), .C2(n31711), .ZN(n9211) );
  OAI222_X1 U29717 ( .A1(n40840), .A2(n40391), .B1(n41224), .B2(n40384), .C1(
        n40379), .C2(n31710), .ZN(n9210) );
  OAI222_X1 U29718 ( .A1(n40846), .A2(n40391), .B1(n41230), .B2(n40384), .C1(
        n40379), .C2(n31709), .ZN(n9209) );
  OAI222_X1 U29719 ( .A1(n40852), .A2(n40391), .B1(n41236), .B2(n40384), .C1(
        n40379), .C2(n31708), .ZN(n9208) );
  OAI222_X1 U29720 ( .A1(n40858), .A2(n40391), .B1(n41242), .B2(n40384), .C1(
        n40379), .C2(n31707), .ZN(n9207) );
  OAI222_X1 U29721 ( .A1(n40864), .A2(n40391), .B1(n41248), .B2(n40384), .C1(
        n40379), .C2(n31706), .ZN(n9206) );
  OAI222_X1 U29722 ( .A1(n40870), .A2(n40391), .B1(n41254), .B2(n40384), .C1(
        n40379), .C2(n31705), .ZN(n9205) );
  OAI222_X1 U29723 ( .A1(n40876), .A2(n40391), .B1(n41260), .B2(n40384), .C1(
        n40379), .C2(n31704), .ZN(n9204) );
  OAI222_X1 U29724 ( .A1(n40882), .A2(n40391), .B1(n41266), .B2(n40384), .C1(
        n40379), .C2(n31703), .ZN(n9203) );
  OAI222_X1 U29725 ( .A1(n40888), .A2(n40391), .B1(n41272), .B2(n40384), .C1(
        n40380), .C2(n31702), .ZN(n9202) );
  OAI222_X1 U29726 ( .A1(n40894), .A2(n40391), .B1(n41278), .B2(n40384), .C1(
        n40380), .C2(n31701), .ZN(n9201) );
  OAI222_X1 U29727 ( .A1(n40900), .A2(n40391), .B1(n41284), .B2(n40384), .C1(
        n40380), .C2(n31700), .ZN(n9200) );
  OAI222_X1 U29728 ( .A1(n40906), .A2(n40391), .B1(n41290), .B2(n40384), .C1(
        n40380), .C2(n31699), .ZN(n9199) );
  OAI222_X1 U29729 ( .A1(n40912), .A2(n40390), .B1(n41296), .B2(n40383), .C1(
        n40380), .C2(n31698), .ZN(n9198) );
  OAI222_X1 U29730 ( .A1(n40918), .A2(n40390), .B1(n41302), .B2(n40383), .C1(
        n40380), .C2(n31697), .ZN(n9197) );
  OAI222_X1 U29731 ( .A1(n40924), .A2(n40390), .B1(n41308), .B2(n40383), .C1(
        n40380), .C2(n31696), .ZN(n9196) );
  OAI222_X1 U29732 ( .A1(n40930), .A2(n40390), .B1(n41314), .B2(n40383), .C1(
        n40380), .C2(n31695), .ZN(n9195) );
  OAI222_X1 U29733 ( .A1(n40936), .A2(n40390), .B1(n41320), .B2(n40383), .C1(
        n40380), .C2(n31694), .ZN(n9194) );
  OAI222_X1 U29734 ( .A1(n40942), .A2(n40390), .B1(n41326), .B2(n40383), .C1(
        n40380), .C2(n31693), .ZN(n9193) );
  OAI222_X1 U29735 ( .A1(n40948), .A2(n40390), .B1(n41332), .B2(n40383), .C1(
        n40380), .C2(n31692), .ZN(n9192) );
  OAI222_X1 U29736 ( .A1(n40960), .A2(n40390), .B1(n41344), .B2(n40383), .C1(
        n40380), .C2(n31690), .ZN(n9190) );
  OAI222_X1 U29737 ( .A1(n40600), .A2(n40375), .B1(n40984), .B2(n40368), .C1(
        n40356), .C2(n31686), .ZN(n9186) );
  OAI222_X1 U29738 ( .A1(n40606), .A2(n40375), .B1(n40990), .B2(n40368), .C1(
        n40356), .C2(n31685), .ZN(n9185) );
  OAI222_X1 U29739 ( .A1(n40612), .A2(n40375), .B1(n40996), .B2(n40368), .C1(
        n40356), .C2(n31684), .ZN(n9184) );
  OAI222_X1 U29740 ( .A1(n40618), .A2(n40375), .B1(n41002), .B2(n40368), .C1(
        n40356), .C2(n31683), .ZN(n9183) );
  OAI222_X1 U29741 ( .A1(n40624), .A2(n40374), .B1(n41008), .B2(n40367), .C1(
        n40356), .C2(n31682), .ZN(n9182) );
  OAI222_X1 U29742 ( .A1(n40630), .A2(n40374), .B1(n41014), .B2(n40367), .C1(
        n40356), .C2(n31681), .ZN(n9181) );
  OAI222_X1 U29743 ( .A1(n40636), .A2(n40374), .B1(n41020), .B2(n40367), .C1(
        n40356), .C2(n31680), .ZN(n9180) );
  OAI222_X1 U29744 ( .A1(n40642), .A2(n40374), .B1(n41026), .B2(n40367), .C1(
        n40356), .C2(n31679), .ZN(n9179) );
  OAI222_X1 U29745 ( .A1(n40648), .A2(n40374), .B1(n41032), .B2(n40367), .C1(
        n40356), .C2(n31678), .ZN(n9178) );
  OAI222_X1 U29746 ( .A1(n40654), .A2(n40374), .B1(n41038), .B2(n40367), .C1(
        n40356), .C2(n31677), .ZN(n9177) );
  OAI222_X1 U29747 ( .A1(n40660), .A2(n40374), .B1(n41044), .B2(n40367), .C1(
        n40356), .C2(n31676), .ZN(n9176) );
  OAI222_X1 U29748 ( .A1(n40666), .A2(n40374), .B1(n41050), .B2(n40367), .C1(
        n40356), .C2(n31675), .ZN(n9175) );
  OAI222_X1 U29749 ( .A1(n40672), .A2(n40374), .B1(n41056), .B2(n40367), .C1(
        n40357), .C2(n31674), .ZN(n9174) );
  OAI222_X1 U29750 ( .A1(n40678), .A2(n40374), .B1(n41062), .B2(n40367), .C1(
        n40357), .C2(n31673), .ZN(n9173) );
  OAI222_X1 U29751 ( .A1(n40684), .A2(n40374), .B1(n41068), .B2(n40367), .C1(
        n40357), .C2(n31672), .ZN(n9172) );
  OAI222_X1 U29752 ( .A1(n40690), .A2(n40374), .B1(n41074), .B2(n40367), .C1(
        n40358), .C2(n31671), .ZN(n9171) );
  OAI222_X1 U29753 ( .A1(n40696), .A2(n40373), .B1(n41080), .B2(n40366), .C1(
        n40357), .C2(n31670), .ZN(n9170) );
  OAI222_X1 U29754 ( .A1(n40702), .A2(n40373), .B1(n41086), .B2(n40366), .C1(
        n40357), .C2(n31669), .ZN(n9169) );
  OAI222_X1 U29755 ( .A1(n40708), .A2(n40373), .B1(n41092), .B2(n40366), .C1(
        n40357), .C2(n31668), .ZN(n9168) );
  OAI222_X1 U29756 ( .A1(n40714), .A2(n40373), .B1(n41098), .B2(n40366), .C1(
        n40357), .C2(n31667), .ZN(n9167) );
  OAI222_X1 U29757 ( .A1(n40720), .A2(n40373), .B1(n41104), .B2(n40366), .C1(
        n40357), .C2(n31666), .ZN(n9166) );
  OAI222_X1 U29758 ( .A1(n40726), .A2(n40373), .B1(n41110), .B2(n40366), .C1(
        n40357), .C2(n31665), .ZN(n9165) );
  OAI222_X1 U29759 ( .A1(n40732), .A2(n40373), .B1(n41116), .B2(n40366), .C1(
        n40357), .C2(n31664), .ZN(n9164) );
  OAI222_X1 U29760 ( .A1(n40738), .A2(n40373), .B1(n41122), .B2(n40366), .C1(
        n40357), .C2(n31663), .ZN(n9163) );
  OAI222_X1 U29761 ( .A1(n40744), .A2(n40373), .B1(n41128), .B2(n40366), .C1(
        n40357), .C2(n31662), .ZN(n9162) );
  OAI222_X1 U29762 ( .A1(n40750), .A2(n40373), .B1(n41134), .B2(n40366), .C1(
        n40358), .C2(n31661), .ZN(n9161) );
  OAI222_X1 U29763 ( .A1(n40756), .A2(n40373), .B1(n41140), .B2(n40366), .C1(
        n40358), .C2(n31660), .ZN(n9160) );
  OAI222_X1 U29764 ( .A1(n40762), .A2(n40373), .B1(n41146), .B2(n40366), .C1(
        n40358), .C2(n31659), .ZN(n9159) );
  OAI222_X1 U29765 ( .A1(n40768), .A2(n40372), .B1(n41152), .B2(n40365), .C1(
        n40358), .C2(n31658), .ZN(n9158) );
  OAI222_X1 U29766 ( .A1(n40774), .A2(n40372), .B1(n41158), .B2(n40365), .C1(
        n40358), .C2(n31657), .ZN(n9157) );
  OAI222_X1 U29767 ( .A1(n40780), .A2(n40372), .B1(n41164), .B2(n40365), .C1(
        n40358), .C2(n31656), .ZN(n9156) );
  OAI222_X1 U29768 ( .A1(n40786), .A2(n40372), .B1(n41170), .B2(n40365), .C1(
        n40358), .C2(n31655), .ZN(n9155) );
  OAI222_X1 U29769 ( .A1(n40792), .A2(n40372), .B1(n41176), .B2(n40365), .C1(
        n40358), .C2(n31654), .ZN(n9154) );
  OAI222_X1 U29770 ( .A1(n40798), .A2(n40372), .B1(n41182), .B2(n40365), .C1(
        n40358), .C2(n31653), .ZN(n9153) );
  OAI222_X1 U29771 ( .A1(n40804), .A2(n40372), .B1(n41188), .B2(n40365), .C1(
        n40358), .C2(n31652), .ZN(n9152) );
  OAI222_X1 U29772 ( .A1(n40810), .A2(n40372), .B1(n41194), .B2(n40365), .C1(
        n40358), .C2(n31651), .ZN(n9151) );
  OAI222_X1 U29773 ( .A1(n40816), .A2(n40372), .B1(n41200), .B2(n40365), .C1(
        n40359), .C2(n31650), .ZN(n9150) );
  OAI222_X1 U29774 ( .A1(n40822), .A2(n40372), .B1(n41206), .B2(n40365), .C1(
        n40359), .C2(n31649), .ZN(n9149) );
  OAI222_X1 U29775 ( .A1(n40828), .A2(n40372), .B1(n41212), .B2(n40365), .C1(
        n40359), .C2(n31648), .ZN(n9148) );
  OAI222_X1 U29776 ( .A1(n40834), .A2(n40372), .B1(n41218), .B2(n40365), .C1(
        n40359), .C2(n31647), .ZN(n9147) );
  OAI222_X1 U29777 ( .A1(n40840), .A2(n40371), .B1(n41224), .B2(n40364), .C1(
        n40359), .C2(n31646), .ZN(n9146) );
  OAI222_X1 U29778 ( .A1(n40846), .A2(n40371), .B1(n41230), .B2(n40364), .C1(
        n40359), .C2(n31645), .ZN(n9145) );
  OAI222_X1 U29779 ( .A1(n40852), .A2(n40371), .B1(n41236), .B2(n40364), .C1(
        n40359), .C2(n31644), .ZN(n9144) );
  OAI222_X1 U29780 ( .A1(n40858), .A2(n40371), .B1(n41242), .B2(n40364), .C1(
        n40359), .C2(n31643), .ZN(n9143) );
  OAI222_X1 U29781 ( .A1(n40864), .A2(n40371), .B1(n41248), .B2(n40364), .C1(
        n40359), .C2(n31642), .ZN(n9142) );
  OAI222_X1 U29782 ( .A1(n40870), .A2(n40371), .B1(n41254), .B2(n40364), .C1(
        n40359), .C2(n31641), .ZN(n9141) );
  OAI222_X1 U29783 ( .A1(n40876), .A2(n40371), .B1(n41260), .B2(n40364), .C1(
        n40359), .C2(n31640), .ZN(n9140) );
  OAI222_X1 U29784 ( .A1(n40882), .A2(n40371), .B1(n41266), .B2(n40364), .C1(
        n40359), .C2(n31639), .ZN(n9139) );
  OAI222_X1 U29785 ( .A1(n40888), .A2(n40371), .B1(n41272), .B2(n40364), .C1(
        n40360), .C2(n31638), .ZN(n9138) );
  OAI222_X1 U29786 ( .A1(n40894), .A2(n40371), .B1(n41278), .B2(n40364), .C1(
        n40360), .C2(n31637), .ZN(n9137) );
  OAI222_X1 U29787 ( .A1(n40900), .A2(n40371), .B1(n41284), .B2(n40364), .C1(
        n40360), .C2(n31636), .ZN(n9136) );
  OAI222_X1 U29788 ( .A1(n40906), .A2(n40371), .B1(n41290), .B2(n40364), .C1(
        n40360), .C2(n31635), .ZN(n9135) );
  OAI222_X1 U29789 ( .A1(n40912), .A2(n40370), .B1(n41296), .B2(n40363), .C1(
        n40360), .C2(n31634), .ZN(n9134) );
  OAI222_X1 U29790 ( .A1(n40918), .A2(n40370), .B1(n41302), .B2(n40363), .C1(
        n40360), .C2(n31633), .ZN(n9133) );
  OAI222_X1 U29791 ( .A1(n40924), .A2(n40370), .B1(n41308), .B2(n40363), .C1(
        n40360), .C2(n31632), .ZN(n9132) );
  OAI222_X1 U29792 ( .A1(n40930), .A2(n40370), .B1(n41314), .B2(n40363), .C1(
        n40360), .C2(n31631), .ZN(n9131) );
  OAI222_X1 U29793 ( .A1(n40936), .A2(n40370), .B1(n41320), .B2(n40363), .C1(
        n40360), .C2(n31630), .ZN(n9130) );
  OAI222_X1 U29794 ( .A1(n40942), .A2(n40370), .B1(n41326), .B2(n40363), .C1(
        n40360), .C2(n31629), .ZN(n9129) );
  OAI222_X1 U29795 ( .A1(n40948), .A2(n40370), .B1(n41332), .B2(n40363), .C1(
        n40360), .C2(n31628), .ZN(n9128) );
  OAI222_X1 U29796 ( .A1(n40960), .A2(n40370), .B1(n41344), .B2(n40363), .C1(
        n40360), .C2(n31626), .ZN(n9126) );
  OAI222_X1 U29797 ( .A1(n40600), .A2(n40355), .B1(n40984), .B2(n40348), .C1(
        n40336), .C2(n31622), .ZN(n9122) );
  OAI222_X1 U29798 ( .A1(n40606), .A2(n40355), .B1(n40990), .B2(n40348), .C1(
        n40336), .C2(n31621), .ZN(n9121) );
  OAI222_X1 U29799 ( .A1(n40612), .A2(n40355), .B1(n40996), .B2(n40348), .C1(
        n40336), .C2(n31620), .ZN(n9120) );
  OAI222_X1 U29800 ( .A1(n40618), .A2(n40355), .B1(n41002), .B2(n40348), .C1(
        n40336), .C2(n31619), .ZN(n9119) );
  OAI222_X1 U29801 ( .A1(n40624), .A2(n40354), .B1(n41008), .B2(n40347), .C1(
        n40336), .C2(n31618), .ZN(n9118) );
  OAI222_X1 U29802 ( .A1(n40630), .A2(n40354), .B1(n41014), .B2(n40347), .C1(
        n40336), .C2(n31617), .ZN(n9117) );
  OAI222_X1 U29803 ( .A1(n40636), .A2(n40354), .B1(n41020), .B2(n40347), .C1(
        n40336), .C2(n31616), .ZN(n9116) );
  OAI222_X1 U29804 ( .A1(n40642), .A2(n40354), .B1(n41026), .B2(n40347), .C1(
        n40336), .C2(n31615), .ZN(n9115) );
  OAI222_X1 U29805 ( .A1(n40648), .A2(n40354), .B1(n41032), .B2(n40347), .C1(
        n40336), .C2(n31614), .ZN(n9114) );
  OAI222_X1 U29806 ( .A1(n40654), .A2(n40354), .B1(n41038), .B2(n40347), .C1(
        n40336), .C2(n31613), .ZN(n9113) );
  OAI222_X1 U29807 ( .A1(n40660), .A2(n40354), .B1(n41044), .B2(n40347), .C1(
        n40336), .C2(n31612), .ZN(n9112) );
  OAI222_X1 U29808 ( .A1(n40666), .A2(n40354), .B1(n41050), .B2(n40347), .C1(
        n40336), .C2(n31611), .ZN(n9111) );
  OAI222_X1 U29809 ( .A1(n40672), .A2(n40354), .B1(n41056), .B2(n40347), .C1(
        n40337), .C2(n31610), .ZN(n9110) );
  OAI222_X1 U29810 ( .A1(n40678), .A2(n40354), .B1(n41062), .B2(n40347), .C1(
        n40337), .C2(n31609), .ZN(n9109) );
  OAI222_X1 U29811 ( .A1(n40684), .A2(n40354), .B1(n41068), .B2(n40347), .C1(
        n40337), .C2(n31608), .ZN(n9108) );
  OAI222_X1 U29812 ( .A1(n40690), .A2(n40354), .B1(n41074), .B2(n40347), .C1(
        n40338), .C2(n31607), .ZN(n9107) );
  OAI222_X1 U29813 ( .A1(n40696), .A2(n40353), .B1(n41080), .B2(n40346), .C1(
        n40337), .C2(n31606), .ZN(n9106) );
  OAI222_X1 U29814 ( .A1(n40702), .A2(n40353), .B1(n41086), .B2(n40346), .C1(
        n40337), .C2(n31605), .ZN(n9105) );
  OAI222_X1 U29815 ( .A1(n40708), .A2(n40353), .B1(n41092), .B2(n40346), .C1(
        n40337), .C2(n31604), .ZN(n9104) );
  OAI222_X1 U29816 ( .A1(n40714), .A2(n40353), .B1(n41098), .B2(n40346), .C1(
        n40337), .C2(n31603), .ZN(n9103) );
  OAI222_X1 U29817 ( .A1(n40720), .A2(n40353), .B1(n41104), .B2(n40346), .C1(
        n40337), .C2(n31602), .ZN(n9102) );
  OAI222_X1 U29818 ( .A1(n40726), .A2(n40353), .B1(n41110), .B2(n40346), .C1(
        n40337), .C2(n31601), .ZN(n9101) );
  OAI222_X1 U29819 ( .A1(n40732), .A2(n40353), .B1(n41116), .B2(n40346), .C1(
        n40337), .C2(n31600), .ZN(n9100) );
  OAI222_X1 U29820 ( .A1(n40738), .A2(n40353), .B1(n41122), .B2(n40346), .C1(
        n40337), .C2(n31599), .ZN(n9099) );
  OAI222_X1 U29821 ( .A1(n40744), .A2(n40353), .B1(n41128), .B2(n40346), .C1(
        n40337), .C2(n31598), .ZN(n9098) );
  OAI222_X1 U29822 ( .A1(n40750), .A2(n40353), .B1(n41134), .B2(n40346), .C1(
        n40338), .C2(n31597), .ZN(n9097) );
  OAI222_X1 U29823 ( .A1(n40756), .A2(n40353), .B1(n41140), .B2(n40346), .C1(
        n40338), .C2(n31596), .ZN(n9096) );
  OAI222_X1 U29824 ( .A1(n40762), .A2(n40353), .B1(n41146), .B2(n40346), .C1(
        n40338), .C2(n31595), .ZN(n9095) );
  OAI222_X1 U29825 ( .A1(n40768), .A2(n40352), .B1(n41152), .B2(n40345), .C1(
        n40338), .C2(n31594), .ZN(n9094) );
  OAI222_X1 U29826 ( .A1(n40774), .A2(n40352), .B1(n41158), .B2(n40345), .C1(
        n40338), .C2(n31593), .ZN(n9093) );
  OAI222_X1 U29827 ( .A1(n40780), .A2(n40352), .B1(n41164), .B2(n40345), .C1(
        n40338), .C2(n31592), .ZN(n9092) );
  OAI222_X1 U29828 ( .A1(n40786), .A2(n40352), .B1(n41170), .B2(n40345), .C1(
        n40338), .C2(n31591), .ZN(n9091) );
  OAI222_X1 U29829 ( .A1(n40792), .A2(n40352), .B1(n41176), .B2(n40345), .C1(
        n40338), .C2(n31590), .ZN(n9090) );
  OAI222_X1 U29830 ( .A1(n40798), .A2(n40352), .B1(n41182), .B2(n40345), .C1(
        n40338), .C2(n31589), .ZN(n9089) );
  OAI222_X1 U29831 ( .A1(n40804), .A2(n40352), .B1(n41188), .B2(n40345), .C1(
        n40338), .C2(n31588), .ZN(n9088) );
  OAI222_X1 U29832 ( .A1(n40810), .A2(n40352), .B1(n41194), .B2(n40345), .C1(
        n40338), .C2(n31587), .ZN(n9087) );
  OAI222_X1 U29833 ( .A1(n40816), .A2(n40352), .B1(n41200), .B2(n40345), .C1(
        n40339), .C2(n31586), .ZN(n9086) );
  OAI222_X1 U29834 ( .A1(n40822), .A2(n40352), .B1(n41206), .B2(n40345), .C1(
        n40339), .C2(n31585), .ZN(n9085) );
  OAI222_X1 U29835 ( .A1(n40828), .A2(n40352), .B1(n41212), .B2(n40345), .C1(
        n40339), .C2(n31584), .ZN(n9084) );
  OAI222_X1 U29836 ( .A1(n40834), .A2(n40352), .B1(n41218), .B2(n40345), .C1(
        n40339), .C2(n31583), .ZN(n9083) );
  OAI222_X1 U29837 ( .A1(n40840), .A2(n40351), .B1(n41224), .B2(n40344), .C1(
        n40339), .C2(n31582), .ZN(n9082) );
  OAI222_X1 U29838 ( .A1(n40846), .A2(n40351), .B1(n41230), .B2(n40344), .C1(
        n40339), .C2(n31581), .ZN(n9081) );
  OAI222_X1 U29839 ( .A1(n40852), .A2(n40351), .B1(n41236), .B2(n40344), .C1(
        n40339), .C2(n31580), .ZN(n9080) );
  OAI222_X1 U29840 ( .A1(n40858), .A2(n40351), .B1(n41242), .B2(n40344), .C1(
        n40339), .C2(n31579), .ZN(n9079) );
  OAI222_X1 U29841 ( .A1(n40864), .A2(n40351), .B1(n41248), .B2(n40344), .C1(
        n40339), .C2(n31578), .ZN(n9078) );
  OAI222_X1 U29842 ( .A1(n40870), .A2(n40351), .B1(n41254), .B2(n40344), .C1(
        n40339), .C2(n31577), .ZN(n9077) );
  OAI222_X1 U29843 ( .A1(n40876), .A2(n40351), .B1(n41260), .B2(n40344), .C1(
        n40339), .C2(n31576), .ZN(n9076) );
  OAI222_X1 U29844 ( .A1(n40882), .A2(n40351), .B1(n41266), .B2(n40344), .C1(
        n40339), .C2(n31575), .ZN(n9075) );
  OAI222_X1 U29845 ( .A1(n40888), .A2(n40351), .B1(n41272), .B2(n40344), .C1(
        n40340), .C2(n31574), .ZN(n9074) );
  OAI222_X1 U29846 ( .A1(n40894), .A2(n40351), .B1(n41278), .B2(n40344), .C1(
        n40340), .C2(n31573), .ZN(n9073) );
  OAI222_X1 U29847 ( .A1(n40900), .A2(n40351), .B1(n41284), .B2(n40344), .C1(
        n40340), .C2(n31572), .ZN(n9072) );
  OAI222_X1 U29848 ( .A1(n40906), .A2(n40351), .B1(n41290), .B2(n40344), .C1(
        n40340), .C2(n31571), .ZN(n9071) );
  OAI222_X1 U29849 ( .A1(n40912), .A2(n40350), .B1(n41296), .B2(n40343), .C1(
        n40340), .C2(n31570), .ZN(n9070) );
  OAI222_X1 U29850 ( .A1(n40918), .A2(n40350), .B1(n41302), .B2(n40343), .C1(
        n40340), .C2(n31569), .ZN(n9069) );
  OAI222_X1 U29851 ( .A1(n40924), .A2(n40350), .B1(n41308), .B2(n40343), .C1(
        n40340), .C2(n31568), .ZN(n9068) );
  OAI222_X1 U29852 ( .A1(n40930), .A2(n40350), .B1(n41314), .B2(n40343), .C1(
        n40340), .C2(n31567), .ZN(n9067) );
  OAI222_X1 U29853 ( .A1(n40936), .A2(n40350), .B1(n41320), .B2(n40343), .C1(
        n40340), .C2(n31566), .ZN(n9066) );
  OAI222_X1 U29854 ( .A1(n40942), .A2(n40350), .B1(n41326), .B2(n40343), .C1(
        n40340), .C2(n31565), .ZN(n9065) );
  OAI222_X1 U29855 ( .A1(n40948), .A2(n40350), .B1(n41332), .B2(n40343), .C1(
        n40340), .C2(n31564), .ZN(n9064) );
  OAI222_X1 U29856 ( .A1(n40960), .A2(n40350), .B1(n41344), .B2(n40343), .C1(
        n40340), .C2(n31562), .ZN(n9062) );
  OAI222_X1 U29857 ( .A1(n40600), .A2(n40295), .B1(n40984), .B2(n40288), .C1(
        n40276), .C2(n31558), .ZN(n8930) );
  OAI222_X1 U29858 ( .A1(n40606), .A2(n40295), .B1(n40990), .B2(n40288), .C1(
        n40276), .C2(n31557), .ZN(n8929) );
  OAI222_X1 U29859 ( .A1(n40612), .A2(n40295), .B1(n40996), .B2(n40288), .C1(
        n40276), .C2(n31556), .ZN(n8928) );
  OAI222_X1 U29860 ( .A1(n40618), .A2(n40295), .B1(n41002), .B2(n40288), .C1(
        n40276), .C2(n31555), .ZN(n8927) );
  OAI222_X1 U29861 ( .A1(n40624), .A2(n40294), .B1(n41008), .B2(n40287), .C1(
        n40276), .C2(n31554), .ZN(n8926) );
  OAI222_X1 U29862 ( .A1(n40630), .A2(n40294), .B1(n41014), .B2(n40287), .C1(
        n40276), .C2(n31553), .ZN(n8925) );
  OAI222_X1 U29863 ( .A1(n40636), .A2(n40294), .B1(n41020), .B2(n40287), .C1(
        n40276), .C2(n31552), .ZN(n8924) );
  OAI222_X1 U29864 ( .A1(n40642), .A2(n40294), .B1(n41026), .B2(n40287), .C1(
        n40276), .C2(n31551), .ZN(n8923) );
  OAI222_X1 U29865 ( .A1(n40648), .A2(n40294), .B1(n41032), .B2(n40287), .C1(
        n40276), .C2(n31550), .ZN(n8922) );
  OAI222_X1 U29866 ( .A1(n40654), .A2(n40294), .B1(n41038), .B2(n40287), .C1(
        n40276), .C2(n31549), .ZN(n8921) );
  OAI222_X1 U29867 ( .A1(n40660), .A2(n40294), .B1(n41044), .B2(n40287), .C1(
        n40276), .C2(n31548), .ZN(n8920) );
  OAI222_X1 U29868 ( .A1(n40666), .A2(n40294), .B1(n41050), .B2(n40287), .C1(
        n40276), .C2(n31547), .ZN(n8919) );
  OAI222_X1 U29869 ( .A1(n40672), .A2(n40294), .B1(n41056), .B2(n40287), .C1(
        n40277), .C2(n31546), .ZN(n8918) );
  OAI222_X1 U29870 ( .A1(n40678), .A2(n40294), .B1(n41062), .B2(n40287), .C1(
        n40277), .C2(n31545), .ZN(n8917) );
  OAI222_X1 U29871 ( .A1(n40684), .A2(n40294), .B1(n41068), .B2(n40287), .C1(
        n40277), .C2(n31544), .ZN(n8916) );
  OAI222_X1 U29872 ( .A1(n40690), .A2(n40294), .B1(n41074), .B2(n40287), .C1(
        n40278), .C2(n31543), .ZN(n8915) );
  OAI222_X1 U29873 ( .A1(n40696), .A2(n40293), .B1(n41080), .B2(n40286), .C1(
        n40277), .C2(n31542), .ZN(n8914) );
  OAI222_X1 U29874 ( .A1(n40702), .A2(n40293), .B1(n41086), .B2(n40286), .C1(
        n40277), .C2(n31541), .ZN(n8913) );
  OAI222_X1 U29875 ( .A1(n40708), .A2(n40293), .B1(n41092), .B2(n40286), .C1(
        n40277), .C2(n31540), .ZN(n8912) );
  OAI222_X1 U29876 ( .A1(n40714), .A2(n40293), .B1(n41098), .B2(n40286), .C1(
        n40277), .C2(n31539), .ZN(n8911) );
  OAI222_X1 U29877 ( .A1(n40720), .A2(n40293), .B1(n41104), .B2(n40286), .C1(
        n40277), .C2(n31538), .ZN(n8910) );
  OAI222_X1 U29878 ( .A1(n40726), .A2(n40293), .B1(n41110), .B2(n40286), .C1(
        n40277), .C2(n31537), .ZN(n8909) );
  OAI222_X1 U29879 ( .A1(n40732), .A2(n40293), .B1(n41116), .B2(n40286), .C1(
        n40277), .C2(n31536), .ZN(n8908) );
  OAI222_X1 U29880 ( .A1(n40738), .A2(n40293), .B1(n41122), .B2(n40286), .C1(
        n40277), .C2(n31535), .ZN(n8907) );
  OAI222_X1 U29881 ( .A1(n40744), .A2(n40293), .B1(n41128), .B2(n40286), .C1(
        n40277), .C2(n31534), .ZN(n8906) );
  OAI222_X1 U29882 ( .A1(n40750), .A2(n40293), .B1(n41134), .B2(n40286), .C1(
        n40278), .C2(n31533), .ZN(n8905) );
  OAI222_X1 U29883 ( .A1(n40756), .A2(n40293), .B1(n41140), .B2(n40286), .C1(
        n40278), .C2(n31532), .ZN(n8904) );
  OAI222_X1 U29884 ( .A1(n40762), .A2(n40293), .B1(n41146), .B2(n40286), .C1(
        n40278), .C2(n31531), .ZN(n8903) );
  OAI222_X1 U29885 ( .A1(n40768), .A2(n40292), .B1(n41152), .B2(n40285), .C1(
        n40278), .C2(n31530), .ZN(n8902) );
  OAI222_X1 U29886 ( .A1(n40774), .A2(n40292), .B1(n41158), .B2(n40285), .C1(
        n40278), .C2(n31529), .ZN(n8901) );
  OAI222_X1 U29887 ( .A1(n40780), .A2(n40292), .B1(n41164), .B2(n40285), .C1(
        n40278), .C2(n31528), .ZN(n8900) );
  OAI222_X1 U29888 ( .A1(n40786), .A2(n40292), .B1(n41170), .B2(n40285), .C1(
        n40278), .C2(n31527), .ZN(n8899) );
  OAI222_X1 U29889 ( .A1(n40792), .A2(n40292), .B1(n41176), .B2(n40285), .C1(
        n40278), .C2(n31526), .ZN(n8898) );
  OAI222_X1 U29890 ( .A1(n40798), .A2(n40292), .B1(n41182), .B2(n40285), .C1(
        n40278), .C2(n31525), .ZN(n8897) );
  OAI222_X1 U29891 ( .A1(n40804), .A2(n40292), .B1(n41188), .B2(n40285), .C1(
        n40278), .C2(n31524), .ZN(n8896) );
  OAI222_X1 U29892 ( .A1(n40810), .A2(n40292), .B1(n41194), .B2(n40285), .C1(
        n40278), .C2(n31523), .ZN(n8895) );
  OAI222_X1 U29893 ( .A1(n40816), .A2(n40292), .B1(n41200), .B2(n40285), .C1(
        n40279), .C2(n31522), .ZN(n8894) );
  OAI222_X1 U29894 ( .A1(n40822), .A2(n40292), .B1(n41206), .B2(n40285), .C1(
        n40279), .C2(n31521), .ZN(n8893) );
  OAI222_X1 U29895 ( .A1(n40828), .A2(n40292), .B1(n41212), .B2(n40285), .C1(
        n40279), .C2(n31520), .ZN(n8892) );
  OAI222_X1 U29896 ( .A1(n40834), .A2(n40292), .B1(n41218), .B2(n40285), .C1(
        n40279), .C2(n31519), .ZN(n8891) );
  OAI222_X1 U29897 ( .A1(n40840), .A2(n40291), .B1(n41224), .B2(n40284), .C1(
        n40279), .C2(n31518), .ZN(n8890) );
  OAI222_X1 U29898 ( .A1(n40846), .A2(n40291), .B1(n41230), .B2(n40284), .C1(
        n40279), .C2(n31517), .ZN(n8889) );
  OAI222_X1 U29899 ( .A1(n40852), .A2(n40291), .B1(n41236), .B2(n40284), .C1(
        n40279), .C2(n31516), .ZN(n8888) );
  OAI222_X1 U29900 ( .A1(n40858), .A2(n40291), .B1(n41242), .B2(n40284), .C1(
        n40279), .C2(n31515), .ZN(n8887) );
  OAI222_X1 U29901 ( .A1(n40864), .A2(n40291), .B1(n41248), .B2(n40284), .C1(
        n40279), .C2(n31514), .ZN(n8886) );
  OAI222_X1 U29902 ( .A1(n40870), .A2(n40291), .B1(n41254), .B2(n40284), .C1(
        n40279), .C2(n31513), .ZN(n8885) );
  OAI222_X1 U29903 ( .A1(n40876), .A2(n40291), .B1(n41260), .B2(n40284), .C1(
        n40279), .C2(n31512), .ZN(n8884) );
  OAI222_X1 U29904 ( .A1(n40882), .A2(n40291), .B1(n41266), .B2(n40284), .C1(
        n40279), .C2(n31511), .ZN(n8883) );
  OAI222_X1 U29905 ( .A1(n40888), .A2(n40291), .B1(n41272), .B2(n40284), .C1(
        n40280), .C2(n31510), .ZN(n8882) );
  OAI222_X1 U29906 ( .A1(n40894), .A2(n40291), .B1(n41278), .B2(n40284), .C1(
        n40280), .C2(n31509), .ZN(n8881) );
  OAI222_X1 U29907 ( .A1(n40900), .A2(n40291), .B1(n41284), .B2(n40284), .C1(
        n40280), .C2(n31508), .ZN(n8880) );
  OAI222_X1 U29908 ( .A1(n40906), .A2(n40291), .B1(n41290), .B2(n40284), .C1(
        n40280), .C2(n31507), .ZN(n8879) );
  OAI222_X1 U29909 ( .A1(n40912), .A2(n40290), .B1(n41296), .B2(n40283), .C1(
        n40280), .C2(n31506), .ZN(n8878) );
  OAI222_X1 U29910 ( .A1(n40918), .A2(n40290), .B1(n41302), .B2(n40283), .C1(
        n40280), .C2(n31505), .ZN(n8877) );
  OAI222_X1 U29911 ( .A1(n40924), .A2(n40290), .B1(n41308), .B2(n40283), .C1(
        n40280), .C2(n31504), .ZN(n8876) );
  OAI222_X1 U29912 ( .A1(n40930), .A2(n40290), .B1(n41314), .B2(n40283), .C1(
        n40280), .C2(n31503), .ZN(n8875) );
  OAI222_X1 U29913 ( .A1(n40936), .A2(n40290), .B1(n41320), .B2(n40283), .C1(
        n40280), .C2(n31502), .ZN(n8874) );
  OAI222_X1 U29914 ( .A1(n40942), .A2(n40290), .B1(n41326), .B2(n40283), .C1(
        n40280), .C2(n31501), .ZN(n8873) );
  OAI222_X1 U29915 ( .A1(n40948), .A2(n40290), .B1(n41332), .B2(n40283), .C1(
        n40280), .C2(n31500), .ZN(n8872) );
  OAI222_X1 U29916 ( .A1(n40960), .A2(n40290), .B1(n41344), .B2(n40283), .C1(
        n40280), .C2(n31498), .ZN(n8870) );
  OAI222_X1 U29917 ( .A1(n40599), .A2(n40275), .B1(n40983), .B2(n40268), .C1(
        n40256), .C2(n31494), .ZN(n8866) );
  OAI222_X1 U29918 ( .A1(n40605), .A2(n40275), .B1(n40989), .B2(n40268), .C1(
        n40256), .C2(n31493), .ZN(n8865) );
  OAI222_X1 U29919 ( .A1(n40611), .A2(n40275), .B1(n40995), .B2(n40268), .C1(
        n40256), .C2(n31492), .ZN(n8864) );
  OAI222_X1 U29920 ( .A1(n40617), .A2(n40275), .B1(n41001), .B2(n40268), .C1(
        n40256), .C2(n31491), .ZN(n8863) );
  OAI222_X1 U29921 ( .A1(n40623), .A2(n40274), .B1(n41007), .B2(n40267), .C1(
        n40256), .C2(n31490), .ZN(n8862) );
  OAI222_X1 U29922 ( .A1(n40629), .A2(n40274), .B1(n41013), .B2(n40267), .C1(
        n40256), .C2(n31489), .ZN(n8861) );
  OAI222_X1 U29923 ( .A1(n40635), .A2(n40274), .B1(n41019), .B2(n40267), .C1(
        n40256), .C2(n31488), .ZN(n8860) );
  OAI222_X1 U29924 ( .A1(n40641), .A2(n40274), .B1(n41025), .B2(n40267), .C1(
        n40256), .C2(n31487), .ZN(n8859) );
  OAI222_X1 U29925 ( .A1(n40647), .A2(n40274), .B1(n41031), .B2(n40267), .C1(
        n40256), .C2(n31486), .ZN(n8858) );
  OAI222_X1 U29926 ( .A1(n40653), .A2(n40274), .B1(n41037), .B2(n40267), .C1(
        n40256), .C2(n31485), .ZN(n8857) );
  OAI222_X1 U29927 ( .A1(n40659), .A2(n40274), .B1(n41043), .B2(n40267), .C1(
        n40256), .C2(n31484), .ZN(n8856) );
  OAI222_X1 U29928 ( .A1(n40665), .A2(n40274), .B1(n41049), .B2(n40267), .C1(
        n40256), .C2(n31483), .ZN(n8855) );
  OAI222_X1 U29929 ( .A1(n40671), .A2(n40274), .B1(n41055), .B2(n40267), .C1(
        n40257), .C2(n31482), .ZN(n8854) );
  OAI222_X1 U29930 ( .A1(n40677), .A2(n40274), .B1(n41061), .B2(n40267), .C1(
        n40257), .C2(n31481), .ZN(n8853) );
  OAI222_X1 U29931 ( .A1(n40683), .A2(n40274), .B1(n41067), .B2(n40267), .C1(
        n40257), .C2(n31480), .ZN(n8852) );
  OAI222_X1 U29932 ( .A1(n40689), .A2(n40274), .B1(n41073), .B2(n40267), .C1(
        n40258), .C2(n31479), .ZN(n8851) );
  OAI222_X1 U29933 ( .A1(n40695), .A2(n40273), .B1(n41079), .B2(n40266), .C1(
        n40257), .C2(n31478), .ZN(n8850) );
  OAI222_X1 U29934 ( .A1(n40701), .A2(n40273), .B1(n41085), .B2(n40266), .C1(
        n40257), .C2(n31477), .ZN(n8849) );
  OAI222_X1 U29935 ( .A1(n40707), .A2(n40273), .B1(n41091), .B2(n40266), .C1(
        n40257), .C2(n31476), .ZN(n8848) );
  OAI222_X1 U29936 ( .A1(n40713), .A2(n40273), .B1(n41097), .B2(n40266), .C1(
        n40257), .C2(n31475), .ZN(n8847) );
  OAI222_X1 U29937 ( .A1(n40719), .A2(n40273), .B1(n41103), .B2(n40266), .C1(
        n40257), .C2(n31474), .ZN(n8846) );
  OAI222_X1 U29938 ( .A1(n40725), .A2(n40273), .B1(n41109), .B2(n40266), .C1(
        n40257), .C2(n31473), .ZN(n8845) );
  OAI222_X1 U29939 ( .A1(n40731), .A2(n40273), .B1(n41115), .B2(n40266), .C1(
        n40257), .C2(n31472), .ZN(n8844) );
  OAI222_X1 U29940 ( .A1(n40737), .A2(n40273), .B1(n41121), .B2(n40266), .C1(
        n40257), .C2(n31471), .ZN(n8843) );
  OAI222_X1 U29941 ( .A1(n40743), .A2(n40273), .B1(n41127), .B2(n40266), .C1(
        n40257), .C2(n31470), .ZN(n8842) );
  OAI222_X1 U29942 ( .A1(n40749), .A2(n40273), .B1(n41133), .B2(n40266), .C1(
        n40258), .C2(n31469), .ZN(n8841) );
  OAI222_X1 U29943 ( .A1(n40755), .A2(n40273), .B1(n41139), .B2(n40266), .C1(
        n40258), .C2(n31468), .ZN(n8840) );
  OAI222_X1 U29944 ( .A1(n40761), .A2(n40273), .B1(n41145), .B2(n40266), .C1(
        n40258), .C2(n31467), .ZN(n8839) );
  OAI222_X1 U29945 ( .A1(n40767), .A2(n40272), .B1(n41151), .B2(n40265), .C1(
        n40258), .C2(n31466), .ZN(n8838) );
  OAI222_X1 U29946 ( .A1(n40773), .A2(n40272), .B1(n41157), .B2(n40265), .C1(
        n40258), .C2(n31465), .ZN(n8837) );
  OAI222_X1 U29947 ( .A1(n40779), .A2(n40272), .B1(n41163), .B2(n40265), .C1(
        n40258), .C2(n31464), .ZN(n8836) );
  OAI222_X1 U29948 ( .A1(n40785), .A2(n40272), .B1(n41169), .B2(n40265), .C1(
        n40258), .C2(n31463), .ZN(n8835) );
  OAI222_X1 U29949 ( .A1(n40791), .A2(n40272), .B1(n41175), .B2(n40265), .C1(
        n40258), .C2(n31462), .ZN(n8834) );
  OAI222_X1 U29950 ( .A1(n40797), .A2(n40272), .B1(n41181), .B2(n40265), .C1(
        n40258), .C2(n31461), .ZN(n8833) );
  OAI222_X1 U29951 ( .A1(n40803), .A2(n40272), .B1(n41187), .B2(n40265), .C1(
        n40258), .C2(n31460), .ZN(n8832) );
  OAI222_X1 U29952 ( .A1(n40809), .A2(n40272), .B1(n41193), .B2(n40265), .C1(
        n40258), .C2(n31459), .ZN(n8831) );
  OAI222_X1 U29953 ( .A1(n40815), .A2(n40272), .B1(n41199), .B2(n40265), .C1(
        n40259), .C2(n31458), .ZN(n8830) );
  OAI222_X1 U29954 ( .A1(n40821), .A2(n40272), .B1(n41205), .B2(n40265), .C1(
        n40259), .C2(n31457), .ZN(n8829) );
  OAI222_X1 U29955 ( .A1(n40827), .A2(n40272), .B1(n41211), .B2(n40265), .C1(
        n40259), .C2(n31456), .ZN(n8828) );
  OAI222_X1 U29956 ( .A1(n40833), .A2(n40272), .B1(n41217), .B2(n40265), .C1(
        n40259), .C2(n31455), .ZN(n8827) );
  OAI222_X1 U29957 ( .A1(n40839), .A2(n40271), .B1(n41223), .B2(n40264), .C1(
        n40259), .C2(n31454), .ZN(n8826) );
  OAI222_X1 U29958 ( .A1(n40845), .A2(n40271), .B1(n41229), .B2(n40264), .C1(
        n40259), .C2(n31453), .ZN(n8825) );
  OAI222_X1 U29959 ( .A1(n40851), .A2(n40271), .B1(n41235), .B2(n40264), .C1(
        n40259), .C2(n31452), .ZN(n8824) );
  OAI222_X1 U29960 ( .A1(n40857), .A2(n40271), .B1(n41241), .B2(n40264), .C1(
        n40259), .C2(n31451), .ZN(n8823) );
  OAI222_X1 U29961 ( .A1(n40863), .A2(n40271), .B1(n41247), .B2(n40264), .C1(
        n40259), .C2(n31450), .ZN(n8822) );
  OAI222_X1 U29962 ( .A1(n40869), .A2(n40271), .B1(n41253), .B2(n40264), .C1(
        n40259), .C2(n31449), .ZN(n8821) );
  OAI222_X1 U29963 ( .A1(n40875), .A2(n40271), .B1(n41259), .B2(n40264), .C1(
        n40259), .C2(n31448), .ZN(n8820) );
  OAI222_X1 U29964 ( .A1(n40881), .A2(n40271), .B1(n41265), .B2(n40264), .C1(
        n40259), .C2(n31447), .ZN(n8819) );
  OAI222_X1 U29965 ( .A1(n40887), .A2(n40271), .B1(n41271), .B2(n40264), .C1(
        n40260), .C2(n31446), .ZN(n8818) );
  OAI222_X1 U29966 ( .A1(n40893), .A2(n40271), .B1(n41277), .B2(n40264), .C1(
        n40260), .C2(n31445), .ZN(n8817) );
  OAI222_X1 U29967 ( .A1(n40899), .A2(n40271), .B1(n41283), .B2(n40264), .C1(
        n40260), .C2(n31444), .ZN(n8816) );
  OAI222_X1 U29968 ( .A1(n40905), .A2(n40271), .B1(n41289), .B2(n40264), .C1(
        n40260), .C2(n31443), .ZN(n8815) );
  OAI222_X1 U29969 ( .A1(n40911), .A2(n40270), .B1(n41295), .B2(n40263), .C1(
        n40260), .C2(n31442), .ZN(n8814) );
  OAI222_X1 U29970 ( .A1(n40917), .A2(n40270), .B1(n41301), .B2(n40263), .C1(
        n40260), .C2(n31441), .ZN(n8813) );
  OAI222_X1 U29971 ( .A1(n40923), .A2(n40270), .B1(n41307), .B2(n40263), .C1(
        n40260), .C2(n31440), .ZN(n8812) );
  OAI222_X1 U29972 ( .A1(n40929), .A2(n40270), .B1(n41313), .B2(n40263), .C1(
        n40260), .C2(n31439), .ZN(n8811) );
  OAI222_X1 U29973 ( .A1(n40935), .A2(n40270), .B1(n41319), .B2(n40263), .C1(
        n40260), .C2(n31438), .ZN(n8810) );
  OAI222_X1 U29974 ( .A1(n40941), .A2(n40270), .B1(n41325), .B2(n40263), .C1(
        n40260), .C2(n31437), .ZN(n8809) );
  OAI222_X1 U29975 ( .A1(n40947), .A2(n40270), .B1(n41331), .B2(n40263), .C1(
        n40260), .C2(n31436), .ZN(n8808) );
  OAI222_X1 U29976 ( .A1(n40959), .A2(n40270), .B1(n41343), .B2(n40263), .C1(
        n40260), .C2(n31434), .ZN(n8806) );
  OAI222_X1 U29977 ( .A1(n40599), .A2(n40255), .B1(n40983), .B2(n40248), .C1(
        n40236), .C2(n31430), .ZN(n8802) );
  OAI222_X1 U29978 ( .A1(n40605), .A2(n40255), .B1(n40989), .B2(n40248), .C1(
        n40236), .C2(n31429), .ZN(n8801) );
  OAI222_X1 U29979 ( .A1(n40611), .A2(n40255), .B1(n40995), .B2(n40248), .C1(
        n40236), .C2(n31428), .ZN(n8800) );
  OAI222_X1 U29980 ( .A1(n40617), .A2(n40255), .B1(n41001), .B2(n40248), .C1(
        n40236), .C2(n31427), .ZN(n8799) );
  OAI222_X1 U29981 ( .A1(n40623), .A2(n40254), .B1(n41007), .B2(n40247), .C1(
        n40236), .C2(n31426), .ZN(n8798) );
  OAI222_X1 U29982 ( .A1(n40629), .A2(n40254), .B1(n41013), .B2(n40247), .C1(
        n40236), .C2(n31425), .ZN(n8797) );
  OAI222_X1 U29983 ( .A1(n40635), .A2(n40254), .B1(n41019), .B2(n40247), .C1(
        n40236), .C2(n31424), .ZN(n8796) );
  OAI222_X1 U29984 ( .A1(n40641), .A2(n40254), .B1(n41025), .B2(n40247), .C1(
        n40236), .C2(n31423), .ZN(n8795) );
  OAI222_X1 U29985 ( .A1(n40647), .A2(n40254), .B1(n41031), .B2(n40247), .C1(
        n40236), .C2(n31422), .ZN(n8794) );
  OAI222_X1 U29986 ( .A1(n40653), .A2(n40254), .B1(n41037), .B2(n40247), .C1(
        n40236), .C2(n31421), .ZN(n8793) );
  OAI222_X1 U29987 ( .A1(n40659), .A2(n40254), .B1(n41043), .B2(n40247), .C1(
        n40236), .C2(n31420), .ZN(n8792) );
  OAI222_X1 U29988 ( .A1(n40665), .A2(n40254), .B1(n41049), .B2(n40247), .C1(
        n40236), .C2(n31419), .ZN(n8791) );
  OAI222_X1 U29989 ( .A1(n40671), .A2(n40254), .B1(n41055), .B2(n40247), .C1(
        n40237), .C2(n31418), .ZN(n8790) );
  OAI222_X1 U29990 ( .A1(n40677), .A2(n40254), .B1(n41061), .B2(n40247), .C1(
        n40237), .C2(n31417), .ZN(n8789) );
  OAI222_X1 U29991 ( .A1(n40683), .A2(n40254), .B1(n41067), .B2(n40247), .C1(
        n40237), .C2(n31416), .ZN(n8788) );
  OAI222_X1 U29992 ( .A1(n40689), .A2(n40254), .B1(n41073), .B2(n40247), .C1(
        n40238), .C2(n31415), .ZN(n8787) );
  OAI222_X1 U29993 ( .A1(n40695), .A2(n40253), .B1(n41079), .B2(n40246), .C1(
        n40237), .C2(n31414), .ZN(n8786) );
  OAI222_X1 U29994 ( .A1(n40701), .A2(n40253), .B1(n41085), .B2(n40246), .C1(
        n40237), .C2(n31413), .ZN(n8785) );
  OAI222_X1 U29995 ( .A1(n40707), .A2(n40253), .B1(n41091), .B2(n40246), .C1(
        n40237), .C2(n31412), .ZN(n8784) );
  OAI222_X1 U29996 ( .A1(n40713), .A2(n40253), .B1(n41097), .B2(n40246), .C1(
        n40237), .C2(n31411), .ZN(n8783) );
  OAI222_X1 U29997 ( .A1(n40719), .A2(n40253), .B1(n41103), .B2(n40246), .C1(
        n40237), .C2(n31410), .ZN(n8782) );
  OAI222_X1 U29998 ( .A1(n40725), .A2(n40253), .B1(n41109), .B2(n40246), .C1(
        n40237), .C2(n31409), .ZN(n8781) );
  OAI222_X1 U29999 ( .A1(n40731), .A2(n40253), .B1(n41115), .B2(n40246), .C1(
        n40237), .C2(n31408), .ZN(n8780) );
  OAI222_X1 U30000 ( .A1(n40737), .A2(n40253), .B1(n41121), .B2(n40246), .C1(
        n40237), .C2(n31407), .ZN(n8779) );
  OAI222_X1 U30001 ( .A1(n40743), .A2(n40253), .B1(n41127), .B2(n40246), .C1(
        n40237), .C2(n31406), .ZN(n8778) );
  OAI222_X1 U30002 ( .A1(n40749), .A2(n40253), .B1(n41133), .B2(n40246), .C1(
        n40238), .C2(n31405), .ZN(n8777) );
  OAI222_X1 U30003 ( .A1(n40755), .A2(n40253), .B1(n41139), .B2(n40246), .C1(
        n40238), .C2(n31404), .ZN(n8776) );
  OAI222_X1 U30004 ( .A1(n40761), .A2(n40253), .B1(n41145), .B2(n40246), .C1(
        n40238), .C2(n31403), .ZN(n8775) );
  OAI222_X1 U30005 ( .A1(n40767), .A2(n40252), .B1(n41151), .B2(n40245), .C1(
        n40238), .C2(n31402), .ZN(n8774) );
  OAI222_X1 U30006 ( .A1(n40773), .A2(n40252), .B1(n41157), .B2(n40245), .C1(
        n40238), .C2(n31401), .ZN(n8773) );
  OAI222_X1 U30007 ( .A1(n40779), .A2(n40252), .B1(n41163), .B2(n40245), .C1(
        n40238), .C2(n31400), .ZN(n8772) );
  OAI222_X1 U30008 ( .A1(n40785), .A2(n40252), .B1(n41169), .B2(n40245), .C1(
        n40238), .C2(n31399), .ZN(n8771) );
  OAI222_X1 U30009 ( .A1(n40791), .A2(n40252), .B1(n41175), .B2(n40245), .C1(
        n40238), .C2(n31398), .ZN(n8770) );
  OAI222_X1 U30010 ( .A1(n40797), .A2(n40252), .B1(n41181), .B2(n40245), .C1(
        n40238), .C2(n31397), .ZN(n8769) );
  OAI222_X1 U30011 ( .A1(n40803), .A2(n40252), .B1(n41187), .B2(n40245), .C1(
        n40238), .C2(n31396), .ZN(n8768) );
  OAI222_X1 U30012 ( .A1(n40809), .A2(n40252), .B1(n41193), .B2(n40245), .C1(
        n40238), .C2(n31395), .ZN(n8767) );
  OAI222_X1 U30013 ( .A1(n40815), .A2(n40252), .B1(n41199), .B2(n40245), .C1(
        n40239), .C2(n31394), .ZN(n8766) );
  OAI222_X1 U30014 ( .A1(n40821), .A2(n40252), .B1(n41205), .B2(n40245), .C1(
        n40239), .C2(n31393), .ZN(n8765) );
  OAI222_X1 U30015 ( .A1(n40827), .A2(n40252), .B1(n41211), .B2(n40245), .C1(
        n40239), .C2(n31392), .ZN(n8764) );
  OAI222_X1 U30016 ( .A1(n40833), .A2(n40252), .B1(n41217), .B2(n40245), .C1(
        n40239), .C2(n31391), .ZN(n8763) );
  OAI222_X1 U30017 ( .A1(n40839), .A2(n40251), .B1(n41223), .B2(n40244), .C1(
        n40239), .C2(n31390), .ZN(n8762) );
  OAI222_X1 U30018 ( .A1(n40845), .A2(n40251), .B1(n41229), .B2(n40244), .C1(
        n40239), .C2(n31389), .ZN(n8761) );
  OAI222_X1 U30019 ( .A1(n40851), .A2(n40251), .B1(n41235), .B2(n40244), .C1(
        n40239), .C2(n31388), .ZN(n8760) );
  OAI222_X1 U30020 ( .A1(n40857), .A2(n40251), .B1(n41241), .B2(n40244), .C1(
        n40239), .C2(n31387), .ZN(n8759) );
  OAI222_X1 U30021 ( .A1(n40863), .A2(n40251), .B1(n41247), .B2(n40244), .C1(
        n40239), .C2(n31386), .ZN(n8758) );
  OAI222_X1 U30022 ( .A1(n40869), .A2(n40251), .B1(n41253), .B2(n40244), .C1(
        n40239), .C2(n31385), .ZN(n8757) );
  OAI222_X1 U30023 ( .A1(n40875), .A2(n40251), .B1(n41259), .B2(n40244), .C1(
        n40239), .C2(n31384), .ZN(n8756) );
  OAI222_X1 U30024 ( .A1(n40881), .A2(n40251), .B1(n41265), .B2(n40244), .C1(
        n40239), .C2(n31383), .ZN(n8755) );
  OAI222_X1 U30025 ( .A1(n40887), .A2(n40251), .B1(n41271), .B2(n40244), .C1(
        n40240), .C2(n31382), .ZN(n8754) );
  OAI222_X1 U30026 ( .A1(n40893), .A2(n40251), .B1(n41277), .B2(n40244), .C1(
        n40240), .C2(n31381), .ZN(n8753) );
  OAI222_X1 U30027 ( .A1(n40899), .A2(n40251), .B1(n41283), .B2(n40244), .C1(
        n40240), .C2(n31380), .ZN(n8752) );
  OAI222_X1 U30028 ( .A1(n40905), .A2(n40251), .B1(n41289), .B2(n40244), .C1(
        n40240), .C2(n31379), .ZN(n8751) );
  OAI222_X1 U30029 ( .A1(n40911), .A2(n40250), .B1(n41295), .B2(n40243), .C1(
        n40240), .C2(n31378), .ZN(n8750) );
  OAI222_X1 U30030 ( .A1(n40917), .A2(n40250), .B1(n41301), .B2(n40243), .C1(
        n40240), .C2(n31377), .ZN(n8749) );
  OAI222_X1 U30031 ( .A1(n40923), .A2(n40250), .B1(n41307), .B2(n40243), .C1(
        n40240), .C2(n31376), .ZN(n8748) );
  OAI222_X1 U30032 ( .A1(n40929), .A2(n40250), .B1(n41313), .B2(n40243), .C1(
        n40240), .C2(n31375), .ZN(n8747) );
  OAI222_X1 U30033 ( .A1(n40935), .A2(n40250), .B1(n41319), .B2(n40243), .C1(
        n40240), .C2(n31374), .ZN(n8746) );
  OAI222_X1 U30034 ( .A1(n40941), .A2(n40250), .B1(n41325), .B2(n40243), .C1(
        n40240), .C2(n31373), .ZN(n8745) );
  OAI222_X1 U30035 ( .A1(n40947), .A2(n40250), .B1(n41331), .B2(n40243), .C1(
        n40240), .C2(n31372), .ZN(n8744) );
  OAI222_X1 U30036 ( .A1(n40959), .A2(n40250), .B1(n41343), .B2(n40243), .C1(
        n40240), .C2(n31370), .ZN(n8742) );
  OAI222_X1 U30037 ( .A1(n40599), .A2(n40195), .B1(n40983), .B2(n40188), .C1(
        n40176), .C2(n31366), .ZN(n8610) );
  OAI222_X1 U30038 ( .A1(n40605), .A2(n40195), .B1(n40989), .B2(n40188), .C1(
        n40176), .C2(n31365), .ZN(n8609) );
  OAI222_X1 U30039 ( .A1(n40611), .A2(n40195), .B1(n40995), .B2(n40188), .C1(
        n40176), .C2(n31364), .ZN(n8608) );
  OAI222_X1 U30040 ( .A1(n40617), .A2(n40195), .B1(n41001), .B2(n40188), .C1(
        n40176), .C2(n31363), .ZN(n8607) );
  OAI222_X1 U30041 ( .A1(n40623), .A2(n40194), .B1(n41007), .B2(n40187), .C1(
        n40176), .C2(n31362), .ZN(n8606) );
  OAI222_X1 U30042 ( .A1(n40629), .A2(n40194), .B1(n41013), .B2(n40187), .C1(
        n40176), .C2(n31361), .ZN(n8605) );
  OAI222_X1 U30043 ( .A1(n40635), .A2(n40194), .B1(n41019), .B2(n40187), .C1(
        n40176), .C2(n31360), .ZN(n8604) );
  OAI222_X1 U30044 ( .A1(n40641), .A2(n40194), .B1(n41025), .B2(n40187), .C1(
        n40176), .C2(n31359), .ZN(n8603) );
  OAI222_X1 U30045 ( .A1(n40647), .A2(n40194), .B1(n41031), .B2(n40187), .C1(
        n40176), .C2(n31358), .ZN(n8602) );
  OAI222_X1 U30046 ( .A1(n40653), .A2(n40194), .B1(n41037), .B2(n40187), .C1(
        n40176), .C2(n31357), .ZN(n8601) );
  OAI222_X1 U30047 ( .A1(n40659), .A2(n40194), .B1(n41043), .B2(n40187), .C1(
        n40176), .C2(n31356), .ZN(n8600) );
  OAI222_X1 U30048 ( .A1(n40665), .A2(n40194), .B1(n41049), .B2(n40187), .C1(
        n40176), .C2(n31355), .ZN(n8599) );
  OAI222_X1 U30049 ( .A1(n40671), .A2(n40194), .B1(n41055), .B2(n40187), .C1(
        n40177), .C2(n31354), .ZN(n8598) );
  OAI222_X1 U30050 ( .A1(n40677), .A2(n40194), .B1(n41061), .B2(n40187), .C1(
        n40177), .C2(n31353), .ZN(n8597) );
  OAI222_X1 U30051 ( .A1(n40683), .A2(n40194), .B1(n41067), .B2(n40187), .C1(
        n40177), .C2(n31352), .ZN(n8596) );
  OAI222_X1 U30052 ( .A1(n40689), .A2(n40194), .B1(n41073), .B2(n40187), .C1(
        n40178), .C2(n31351), .ZN(n8595) );
  OAI222_X1 U30053 ( .A1(n40695), .A2(n40193), .B1(n41079), .B2(n40186), .C1(
        n40177), .C2(n31350), .ZN(n8594) );
  OAI222_X1 U30054 ( .A1(n40701), .A2(n40193), .B1(n41085), .B2(n40186), .C1(
        n40177), .C2(n31349), .ZN(n8593) );
  OAI222_X1 U30055 ( .A1(n40707), .A2(n40193), .B1(n41091), .B2(n40186), .C1(
        n40177), .C2(n31348), .ZN(n8592) );
  OAI222_X1 U30056 ( .A1(n40713), .A2(n40193), .B1(n41097), .B2(n40186), .C1(
        n40177), .C2(n31347), .ZN(n8591) );
  OAI222_X1 U30057 ( .A1(n40719), .A2(n40193), .B1(n41103), .B2(n40186), .C1(
        n40177), .C2(n31346), .ZN(n8590) );
  OAI222_X1 U30058 ( .A1(n40725), .A2(n40193), .B1(n41109), .B2(n40186), .C1(
        n40177), .C2(n31345), .ZN(n8589) );
  OAI222_X1 U30059 ( .A1(n40731), .A2(n40193), .B1(n41115), .B2(n40186), .C1(
        n40177), .C2(n31344), .ZN(n8588) );
  OAI222_X1 U30060 ( .A1(n40737), .A2(n40193), .B1(n41121), .B2(n40186), .C1(
        n40177), .C2(n31343), .ZN(n8587) );
  OAI222_X1 U30061 ( .A1(n40743), .A2(n40193), .B1(n41127), .B2(n40186), .C1(
        n40177), .C2(n31342), .ZN(n8586) );
  OAI222_X1 U30062 ( .A1(n40749), .A2(n40193), .B1(n41133), .B2(n40186), .C1(
        n40178), .C2(n31341), .ZN(n8585) );
  OAI222_X1 U30063 ( .A1(n40755), .A2(n40193), .B1(n41139), .B2(n40186), .C1(
        n40178), .C2(n31340), .ZN(n8584) );
  OAI222_X1 U30064 ( .A1(n40761), .A2(n40193), .B1(n41145), .B2(n40186), .C1(
        n40178), .C2(n31339), .ZN(n8583) );
  OAI222_X1 U30065 ( .A1(n40767), .A2(n40192), .B1(n41151), .B2(n40185), .C1(
        n40178), .C2(n31338), .ZN(n8582) );
  OAI222_X1 U30066 ( .A1(n40773), .A2(n40192), .B1(n41157), .B2(n40185), .C1(
        n40178), .C2(n31337), .ZN(n8581) );
  OAI222_X1 U30067 ( .A1(n40779), .A2(n40192), .B1(n41163), .B2(n40185), .C1(
        n40178), .C2(n31336), .ZN(n8580) );
  OAI222_X1 U30068 ( .A1(n40785), .A2(n40192), .B1(n41169), .B2(n40185), .C1(
        n40178), .C2(n31335), .ZN(n8579) );
  OAI222_X1 U30069 ( .A1(n40791), .A2(n40192), .B1(n41175), .B2(n40185), .C1(
        n40178), .C2(n31334), .ZN(n8578) );
  OAI222_X1 U30070 ( .A1(n40797), .A2(n40192), .B1(n41181), .B2(n40185), .C1(
        n40178), .C2(n31333), .ZN(n8577) );
  OAI222_X1 U30071 ( .A1(n40803), .A2(n40192), .B1(n41187), .B2(n40185), .C1(
        n40178), .C2(n31332), .ZN(n8576) );
  OAI222_X1 U30072 ( .A1(n40809), .A2(n40192), .B1(n41193), .B2(n40185), .C1(
        n40178), .C2(n31331), .ZN(n8575) );
  OAI222_X1 U30073 ( .A1(n40815), .A2(n40192), .B1(n41199), .B2(n40185), .C1(
        n40179), .C2(n31330), .ZN(n8574) );
  OAI222_X1 U30074 ( .A1(n40821), .A2(n40192), .B1(n41205), .B2(n40185), .C1(
        n40179), .C2(n31329), .ZN(n8573) );
  OAI222_X1 U30075 ( .A1(n40827), .A2(n40192), .B1(n41211), .B2(n40185), .C1(
        n40179), .C2(n31328), .ZN(n8572) );
  OAI222_X1 U30076 ( .A1(n40833), .A2(n40192), .B1(n41217), .B2(n40185), .C1(
        n40179), .C2(n31327), .ZN(n8571) );
  OAI222_X1 U30077 ( .A1(n40839), .A2(n40191), .B1(n41223), .B2(n40184), .C1(
        n40179), .C2(n31326), .ZN(n8570) );
  OAI222_X1 U30078 ( .A1(n40845), .A2(n40191), .B1(n41229), .B2(n40184), .C1(
        n40179), .C2(n31325), .ZN(n8569) );
  OAI222_X1 U30079 ( .A1(n40851), .A2(n40191), .B1(n41235), .B2(n40184), .C1(
        n40179), .C2(n31324), .ZN(n8568) );
  OAI222_X1 U30080 ( .A1(n40857), .A2(n40191), .B1(n41241), .B2(n40184), .C1(
        n40179), .C2(n31323), .ZN(n8567) );
  OAI222_X1 U30081 ( .A1(n40863), .A2(n40191), .B1(n41247), .B2(n40184), .C1(
        n40179), .C2(n31322), .ZN(n8566) );
  OAI222_X1 U30082 ( .A1(n40869), .A2(n40191), .B1(n41253), .B2(n40184), .C1(
        n40179), .C2(n31321), .ZN(n8565) );
  OAI222_X1 U30083 ( .A1(n40875), .A2(n40191), .B1(n41259), .B2(n40184), .C1(
        n40179), .C2(n31320), .ZN(n8564) );
  OAI222_X1 U30084 ( .A1(n40881), .A2(n40191), .B1(n41265), .B2(n40184), .C1(
        n40179), .C2(n31319), .ZN(n8563) );
  OAI222_X1 U30085 ( .A1(n40887), .A2(n40191), .B1(n41271), .B2(n40184), .C1(
        n40180), .C2(n31318), .ZN(n8562) );
  OAI222_X1 U30086 ( .A1(n40893), .A2(n40191), .B1(n41277), .B2(n40184), .C1(
        n40180), .C2(n31317), .ZN(n8561) );
  OAI222_X1 U30087 ( .A1(n40899), .A2(n40191), .B1(n41283), .B2(n40184), .C1(
        n40180), .C2(n31316), .ZN(n8560) );
  OAI222_X1 U30088 ( .A1(n40905), .A2(n40191), .B1(n41289), .B2(n40184), .C1(
        n40180), .C2(n31315), .ZN(n8559) );
  OAI222_X1 U30089 ( .A1(n40911), .A2(n40190), .B1(n41295), .B2(n40183), .C1(
        n40180), .C2(n31314), .ZN(n8558) );
  OAI222_X1 U30090 ( .A1(n40917), .A2(n40190), .B1(n41301), .B2(n40183), .C1(
        n40180), .C2(n31313), .ZN(n8557) );
  OAI222_X1 U30091 ( .A1(n40923), .A2(n40190), .B1(n41307), .B2(n40183), .C1(
        n40180), .C2(n31312), .ZN(n8556) );
  OAI222_X1 U30092 ( .A1(n40929), .A2(n40190), .B1(n41313), .B2(n40183), .C1(
        n40180), .C2(n31311), .ZN(n8555) );
  OAI222_X1 U30093 ( .A1(n40935), .A2(n40190), .B1(n41319), .B2(n40183), .C1(
        n40180), .C2(n31310), .ZN(n8554) );
  OAI222_X1 U30094 ( .A1(n40941), .A2(n40190), .B1(n41325), .B2(n40183), .C1(
        n40180), .C2(n31309), .ZN(n8553) );
  OAI222_X1 U30095 ( .A1(n40947), .A2(n40190), .B1(n41331), .B2(n40183), .C1(
        n40180), .C2(n31308), .ZN(n8552) );
  OAI222_X1 U30096 ( .A1(n40959), .A2(n40190), .B1(n41343), .B2(n40183), .C1(
        n40180), .C2(n31306), .ZN(n8550) );
  OAI222_X1 U30097 ( .A1(n40599), .A2(n40175), .B1(n40983), .B2(n40168), .C1(
        n40156), .C2(n31302), .ZN(n8546) );
  OAI222_X1 U30098 ( .A1(n40605), .A2(n40175), .B1(n40989), .B2(n40168), .C1(
        n40156), .C2(n31301), .ZN(n8545) );
  OAI222_X1 U30099 ( .A1(n40611), .A2(n40175), .B1(n40995), .B2(n40168), .C1(
        n40156), .C2(n31300), .ZN(n8544) );
  OAI222_X1 U30100 ( .A1(n40617), .A2(n40175), .B1(n41001), .B2(n40168), .C1(
        n40156), .C2(n31299), .ZN(n8543) );
  OAI222_X1 U30101 ( .A1(n40623), .A2(n40174), .B1(n41007), .B2(n40167), .C1(
        n40156), .C2(n31298), .ZN(n8542) );
  OAI222_X1 U30102 ( .A1(n40629), .A2(n40174), .B1(n41013), .B2(n40167), .C1(
        n40156), .C2(n31297), .ZN(n8541) );
  OAI222_X1 U30103 ( .A1(n40635), .A2(n40174), .B1(n41019), .B2(n40167), .C1(
        n40156), .C2(n31296), .ZN(n8540) );
  OAI222_X1 U30104 ( .A1(n40641), .A2(n40174), .B1(n41025), .B2(n40167), .C1(
        n40156), .C2(n31295), .ZN(n8539) );
  OAI222_X1 U30105 ( .A1(n40647), .A2(n40174), .B1(n41031), .B2(n40167), .C1(
        n40156), .C2(n31294), .ZN(n8538) );
  OAI222_X1 U30106 ( .A1(n40653), .A2(n40174), .B1(n41037), .B2(n40167), .C1(
        n40156), .C2(n31293), .ZN(n8537) );
  OAI222_X1 U30107 ( .A1(n40659), .A2(n40174), .B1(n41043), .B2(n40167), .C1(
        n40156), .C2(n31292), .ZN(n8536) );
  OAI222_X1 U30108 ( .A1(n40665), .A2(n40174), .B1(n41049), .B2(n40167), .C1(
        n40156), .C2(n31291), .ZN(n8535) );
  OAI222_X1 U30109 ( .A1(n40671), .A2(n40174), .B1(n41055), .B2(n40167), .C1(
        n40157), .C2(n31290), .ZN(n8534) );
  OAI222_X1 U30110 ( .A1(n40677), .A2(n40174), .B1(n41061), .B2(n40167), .C1(
        n40157), .C2(n31289), .ZN(n8533) );
  OAI222_X1 U30111 ( .A1(n40683), .A2(n40174), .B1(n41067), .B2(n40167), .C1(
        n40157), .C2(n31288), .ZN(n8532) );
  OAI222_X1 U30112 ( .A1(n40689), .A2(n40174), .B1(n41073), .B2(n40167), .C1(
        n40158), .C2(n31287), .ZN(n8531) );
  OAI222_X1 U30113 ( .A1(n40695), .A2(n40173), .B1(n41079), .B2(n40166), .C1(
        n40157), .C2(n31286), .ZN(n8530) );
  OAI222_X1 U30114 ( .A1(n40701), .A2(n40173), .B1(n41085), .B2(n40166), .C1(
        n40157), .C2(n31285), .ZN(n8529) );
  OAI222_X1 U30115 ( .A1(n40707), .A2(n40173), .B1(n41091), .B2(n40166), .C1(
        n40157), .C2(n31284), .ZN(n8528) );
  OAI222_X1 U30116 ( .A1(n40713), .A2(n40173), .B1(n41097), .B2(n40166), .C1(
        n40157), .C2(n31283), .ZN(n8527) );
  OAI222_X1 U30117 ( .A1(n40719), .A2(n40173), .B1(n41103), .B2(n40166), .C1(
        n40157), .C2(n31282), .ZN(n8526) );
  OAI222_X1 U30118 ( .A1(n40725), .A2(n40173), .B1(n41109), .B2(n40166), .C1(
        n40157), .C2(n31281), .ZN(n8525) );
  OAI222_X1 U30119 ( .A1(n40731), .A2(n40173), .B1(n41115), .B2(n40166), .C1(
        n40157), .C2(n31280), .ZN(n8524) );
  OAI222_X1 U30120 ( .A1(n40737), .A2(n40173), .B1(n41121), .B2(n40166), .C1(
        n40157), .C2(n31279), .ZN(n8523) );
  OAI222_X1 U30121 ( .A1(n40743), .A2(n40173), .B1(n41127), .B2(n40166), .C1(
        n40157), .C2(n31278), .ZN(n8522) );
  OAI222_X1 U30122 ( .A1(n40749), .A2(n40173), .B1(n41133), .B2(n40166), .C1(
        n40158), .C2(n31277), .ZN(n8521) );
  OAI222_X1 U30123 ( .A1(n40755), .A2(n40173), .B1(n41139), .B2(n40166), .C1(
        n40158), .C2(n31276), .ZN(n8520) );
  OAI222_X1 U30124 ( .A1(n40761), .A2(n40173), .B1(n41145), .B2(n40166), .C1(
        n40158), .C2(n31275), .ZN(n8519) );
  OAI222_X1 U30125 ( .A1(n40767), .A2(n40172), .B1(n41151), .B2(n40165), .C1(
        n40158), .C2(n31274), .ZN(n8518) );
  OAI222_X1 U30126 ( .A1(n40773), .A2(n40172), .B1(n41157), .B2(n40165), .C1(
        n40158), .C2(n31273), .ZN(n8517) );
  OAI222_X1 U30127 ( .A1(n40779), .A2(n40172), .B1(n41163), .B2(n40165), .C1(
        n40158), .C2(n31272), .ZN(n8516) );
  OAI222_X1 U30128 ( .A1(n40785), .A2(n40172), .B1(n41169), .B2(n40165), .C1(
        n40158), .C2(n31271), .ZN(n8515) );
  OAI222_X1 U30129 ( .A1(n40791), .A2(n40172), .B1(n41175), .B2(n40165), .C1(
        n40158), .C2(n31270), .ZN(n8514) );
  OAI222_X1 U30130 ( .A1(n40797), .A2(n40172), .B1(n41181), .B2(n40165), .C1(
        n40158), .C2(n31269), .ZN(n8513) );
  OAI222_X1 U30131 ( .A1(n40803), .A2(n40172), .B1(n41187), .B2(n40165), .C1(
        n40158), .C2(n31268), .ZN(n8512) );
  OAI222_X1 U30132 ( .A1(n40809), .A2(n40172), .B1(n41193), .B2(n40165), .C1(
        n40158), .C2(n31267), .ZN(n8511) );
  OAI222_X1 U30133 ( .A1(n40815), .A2(n40172), .B1(n41199), .B2(n40165), .C1(
        n40159), .C2(n31266), .ZN(n8510) );
  OAI222_X1 U30134 ( .A1(n40821), .A2(n40172), .B1(n41205), .B2(n40165), .C1(
        n40159), .C2(n31265), .ZN(n8509) );
  OAI222_X1 U30135 ( .A1(n40827), .A2(n40172), .B1(n41211), .B2(n40165), .C1(
        n40159), .C2(n31264), .ZN(n8508) );
  OAI222_X1 U30136 ( .A1(n40833), .A2(n40172), .B1(n41217), .B2(n40165), .C1(
        n40159), .C2(n31263), .ZN(n8507) );
  OAI222_X1 U30137 ( .A1(n40839), .A2(n40171), .B1(n41223), .B2(n40164), .C1(
        n40159), .C2(n31262), .ZN(n8506) );
  OAI222_X1 U30138 ( .A1(n40845), .A2(n40171), .B1(n41229), .B2(n40164), .C1(
        n40159), .C2(n31261), .ZN(n8505) );
  OAI222_X1 U30139 ( .A1(n40851), .A2(n40171), .B1(n41235), .B2(n40164), .C1(
        n40159), .C2(n31260), .ZN(n8504) );
  OAI222_X1 U30140 ( .A1(n40857), .A2(n40171), .B1(n41241), .B2(n40164), .C1(
        n40159), .C2(n31259), .ZN(n8503) );
  OAI222_X1 U30141 ( .A1(n40863), .A2(n40171), .B1(n41247), .B2(n40164), .C1(
        n40159), .C2(n31258), .ZN(n8502) );
  OAI222_X1 U30142 ( .A1(n40869), .A2(n40171), .B1(n41253), .B2(n40164), .C1(
        n40159), .C2(n31257), .ZN(n8501) );
  OAI222_X1 U30143 ( .A1(n40875), .A2(n40171), .B1(n41259), .B2(n40164), .C1(
        n40159), .C2(n31256), .ZN(n8500) );
  OAI222_X1 U30144 ( .A1(n40881), .A2(n40171), .B1(n41265), .B2(n40164), .C1(
        n40159), .C2(n31255), .ZN(n8499) );
  OAI222_X1 U30145 ( .A1(n40887), .A2(n40171), .B1(n41271), .B2(n40164), .C1(
        n40160), .C2(n31254), .ZN(n8498) );
  OAI222_X1 U30146 ( .A1(n40893), .A2(n40171), .B1(n41277), .B2(n40164), .C1(
        n40160), .C2(n31253), .ZN(n8497) );
  OAI222_X1 U30147 ( .A1(n40899), .A2(n40171), .B1(n41283), .B2(n40164), .C1(
        n40160), .C2(n31252), .ZN(n8496) );
  OAI222_X1 U30148 ( .A1(n40905), .A2(n40171), .B1(n41289), .B2(n40164), .C1(
        n40160), .C2(n31251), .ZN(n8495) );
  OAI222_X1 U30149 ( .A1(n40911), .A2(n40170), .B1(n41295), .B2(n40163), .C1(
        n40160), .C2(n31250), .ZN(n8494) );
  OAI222_X1 U30150 ( .A1(n40917), .A2(n40170), .B1(n41301), .B2(n40163), .C1(
        n40160), .C2(n31249), .ZN(n8493) );
  OAI222_X1 U30151 ( .A1(n40923), .A2(n40170), .B1(n41307), .B2(n40163), .C1(
        n40160), .C2(n31248), .ZN(n8492) );
  OAI222_X1 U30152 ( .A1(n40929), .A2(n40170), .B1(n41313), .B2(n40163), .C1(
        n40160), .C2(n31247), .ZN(n8491) );
  OAI222_X1 U30153 ( .A1(n40935), .A2(n40170), .B1(n41319), .B2(n40163), .C1(
        n40160), .C2(n31246), .ZN(n8490) );
  OAI222_X1 U30154 ( .A1(n40941), .A2(n40170), .B1(n41325), .B2(n40163), .C1(
        n40160), .C2(n31245), .ZN(n8489) );
  OAI222_X1 U30155 ( .A1(n40947), .A2(n40170), .B1(n41331), .B2(n40163), .C1(
        n40160), .C2(n31244), .ZN(n8488) );
  OAI222_X1 U30156 ( .A1(n40959), .A2(n40170), .B1(n41343), .B2(n40163), .C1(
        n40160), .C2(n31242), .ZN(n8486) );
  OAI222_X1 U30157 ( .A1(n40599), .A2(n40155), .B1(n40983), .B2(n40148), .C1(
        n40136), .C2(n31238), .ZN(n8482) );
  OAI222_X1 U30158 ( .A1(n40605), .A2(n40155), .B1(n40989), .B2(n40148), .C1(
        n40136), .C2(n31237), .ZN(n8481) );
  OAI222_X1 U30159 ( .A1(n40611), .A2(n40155), .B1(n40995), .B2(n40148), .C1(
        n40136), .C2(n31236), .ZN(n8480) );
  OAI222_X1 U30160 ( .A1(n40617), .A2(n40155), .B1(n41001), .B2(n40148), .C1(
        n40136), .C2(n31235), .ZN(n8479) );
  OAI222_X1 U30161 ( .A1(n40623), .A2(n40154), .B1(n41007), .B2(n40147), .C1(
        n40136), .C2(n31234), .ZN(n8478) );
  OAI222_X1 U30162 ( .A1(n40629), .A2(n40154), .B1(n41013), .B2(n40147), .C1(
        n40136), .C2(n31233), .ZN(n8477) );
  OAI222_X1 U30163 ( .A1(n40635), .A2(n40154), .B1(n41019), .B2(n40147), .C1(
        n40136), .C2(n31232), .ZN(n8476) );
  OAI222_X1 U30164 ( .A1(n40641), .A2(n40154), .B1(n41025), .B2(n40147), .C1(
        n40136), .C2(n31231), .ZN(n8475) );
  OAI222_X1 U30165 ( .A1(n40647), .A2(n40154), .B1(n41031), .B2(n40147), .C1(
        n40136), .C2(n31230), .ZN(n8474) );
  OAI222_X1 U30166 ( .A1(n40653), .A2(n40154), .B1(n41037), .B2(n40147), .C1(
        n40136), .C2(n31229), .ZN(n8473) );
  OAI222_X1 U30167 ( .A1(n40659), .A2(n40154), .B1(n41043), .B2(n40147), .C1(
        n40136), .C2(n31228), .ZN(n8472) );
  OAI222_X1 U30168 ( .A1(n40665), .A2(n40154), .B1(n41049), .B2(n40147), .C1(
        n40136), .C2(n31227), .ZN(n8471) );
  OAI222_X1 U30169 ( .A1(n40671), .A2(n40154), .B1(n41055), .B2(n40147), .C1(
        n40137), .C2(n31226), .ZN(n8470) );
  OAI222_X1 U30170 ( .A1(n40677), .A2(n40154), .B1(n41061), .B2(n40147), .C1(
        n40137), .C2(n31225), .ZN(n8469) );
  OAI222_X1 U30171 ( .A1(n40683), .A2(n40154), .B1(n41067), .B2(n40147), .C1(
        n40137), .C2(n31224), .ZN(n8468) );
  OAI222_X1 U30172 ( .A1(n40689), .A2(n40154), .B1(n41073), .B2(n40147), .C1(
        n40138), .C2(n31223), .ZN(n8467) );
  OAI222_X1 U30173 ( .A1(n40695), .A2(n40153), .B1(n41079), .B2(n40146), .C1(
        n40137), .C2(n31222), .ZN(n8466) );
  OAI222_X1 U30174 ( .A1(n40701), .A2(n40153), .B1(n41085), .B2(n40146), .C1(
        n40137), .C2(n31221), .ZN(n8465) );
  OAI222_X1 U30175 ( .A1(n40707), .A2(n40153), .B1(n41091), .B2(n40146), .C1(
        n40137), .C2(n31220), .ZN(n8464) );
  OAI222_X1 U30176 ( .A1(n40713), .A2(n40153), .B1(n41097), .B2(n40146), .C1(
        n40137), .C2(n31219), .ZN(n8463) );
  OAI222_X1 U30177 ( .A1(n40719), .A2(n40153), .B1(n41103), .B2(n40146), .C1(
        n40137), .C2(n31218), .ZN(n8462) );
  OAI222_X1 U30178 ( .A1(n40725), .A2(n40153), .B1(n41109), .B2(n40146), .C1(
        n40137), .C2(n31217), .ZN(n8461) );
  OAI222_X1 U30179 ( .A1(n40731), .A2(n40153), .B1(n41115), .B2(n40146), .C1(
        n40137), .C2(n31216), .ZN(n8460) );
  OAI222_X1 U30180 ( .A1(n40737), .A2(n40153), .B1(n41121), .B2(n40146), .C1(
        n40137), .C2(n31215), .ZN(n8459) );
  OAI222_X1 U30181 ( .A1(n40743), .A2(n40153), .B1(n41127), .B2(n40146), .C1(
        n40137), .C2(n31214), .ZN(n8458) );
  OAI222_X1 U30182 ( .A1(n40749), .A2(n40153), .B1(n41133), .B2(n40146), .C1(
        n40138), .C2(n31213), .ZN(n8457) );
  OAI222_X1 U30183 ( .A1(n40755), .A2(n40153), .B1(n41139), .B2(n40146), .C1(
        n40138), .C2(n31212), .ZN(n8456) );
  OAI222_X1 U30184 ( .A1(n40761), .A2(n40153), .B1(n41145), .B2(n40146), .C1(
        n40138), .C2(n31211), .ZN(n8455) );
  OAI222_X1 U30185 ( .A1(n40767), .A2(n40152), .B1(n41151), .B2(n40145), .C1(
        n40138), .C2(n31210), .ZN(n8454) );
  OAI222_X1 U30186 ( .A1(n40773), .A2(n40152), .B1(n41157), .B2(n40145), .C1(
        n40138), .C2(n31209), .ZN(n8453) );
  OAI222_X1 U30187 ( .A1(n40779), .A2(n40152), .B1(n41163), .B2(n40145), .C1(
        n40138), .C2(n31208), .ZN(n8452) );
  OAI222_X1 U30188 ( .A1(n40785), .A2(n40152), .B1(n41169), .B2(n40145), .C1(
        n40138), .C2(n31207), .ZN(n8451) );
  OAI222_X1 U30189 ( .A1(n40791), .A2(n40152), .B1(n41175), .B2(n40145), .C1(
        n40138), .C2(n31206), .ZN(n8450) );
  OAI222_X1 U30190 ( .A1(n40797), .A2(n40152), .B1(n41181), .B2(n40145), .C1(
        n40138), .C2(n31205), .ZN(n8449) );
  OAI222_X1 U30191 ( .A1(n40803), .A2(n40152), .B1(n41187), .B2(n40145), .C1(
        n40138), .C2(n31204), .ZN(n8448) );
  OAI222_X1 U30192 ( .A1(n40809), .A2(n40152), .B1(n41193), .B2(n40145), .C1(
        n40138), .C2(n31203), .ZN(n8447) );
  OAI222_X1 U30193 ( .A1(n40815), .A2(n40152), .B1(n41199), .B2(n40145), .C1(
        n40139), .C2(n31202), .ZN(n8446) );
  OAI222_X1 U30194 ( .A1(n40821), .A2(n40152), .B1(n41205), .B2(n40145), .C1(
        n40139), .C2(n31201), .ZN(n8445) );
  OAI222_X1 U30195 ( .A1(n40827), .A2(n40152), .B1(n41211), .B2(n40145), .C1(
        n40139), .C2(n31200), .ZN(n8444) );
  OAI222_X1 U30196 ( .A1(n40833), .A2(n40152), .B1(n41217), .B2(n40145), .C1(
        n40139), .C2(n31199), .ZN(n8443) );
  OAI222_X1 U30197 ( .A1(n40839), .A2(n40151), .B1(n41223), .B2(n40144), .C1(
        n40139), .C2(n31198), .ZN(n8442) );
  OAI222_X1 U30198 ( .A1(n40845), .A2(n40151), .B1(n41229), .B2(n40144), .C1(
        n40139), .C2(n31197), .ZN(n8441) );
  OAI222_X1 U30199 ( .A1(n40851), .A2(n40151), .B1(n41235), .B2(n40144), .C1(
        n40139), .C2(n31196), .ZN(n8440) );
  OAI222_X1 U30200 ( .A1(n40857), .A2(n40151), .B1(n41241), .B2(n40144), .C1(
        n40139), .C2(n31195), .ZN(n8439) );
  OAI222_X1 U30201 ( .A1(n40863), .A2(n40151), .B1(n41247), .B2(n40144), .C1(
        n40139), .C2(n31194), .ZN(n8438) );
  OAI222_X1 U30202 ( .A1(n40869), .A2(n40151), .B1(n41253), .B2(n40144), .C1(
        n40139), .C2(n31193), .ZN(n8437) );
  OAI222_X1 U30203 ( .A1(n40875), .A2(n40151), .B1(n41259), .B2(n40144), .C1(
        n40139), .C2(n31192), .ZN(n8436) );
  OAI222_X1 U30204 ( .A1(n40881), .A2(n40151), .B1(n41265), .B2(n40144), .C1(
        n40139), .C2(n31191), .ZN(n8435) );
  OAI222_X1 U30205 ( .A1(n40887), .A2(n40151), .B1(n41271), .B2(n40144), .C1(
        n40140), .C2(n31190), .ZN(n8434) );
  OAI222_X1 U30206 ( .A1(n40893), .A2(n40151), .B1(n41277), .B2(n40144), .C1(
        n40140), .C2(n31189), .ZN(n8433) );
  OAI222_X1 U30207 ( .A1(n40899), .A2(n40151), .B1(n41283), .B2(n40144), .C1(
        n40140), .C2(n31188), .ZN(n8432) );
  OAI222_X1 U30208 ( .A1(n40905), .A2(n40151), .B1(n41289), .B2(n40144), .C1(
        n40140), .C2(n31187), .ZN(n8431) );
  OAI222_X1 U30209 ( .A1(n40911), .A2(n40150), .B1(n41295), .B2(n40143), .C1(
        n40140), .C2(n31186), .ZN(n8430) );
  OAI222_X1 U30210 ( .A1(n40917), .A2(n40150), .B1(n41301), .B2(n40143), .C1(
        n40140), .C2(n31185), .ZN(n8429) );
  OAI222_X1 U30211 ( .A1(n40923), .A2(n40150), .B1(n41307), .B2(n40143), .C1(
        n40140), .C2(n31184), .ZN(n8428) );
  OAI222_X1 U30212 ( .A1(n40929), .A2(n40150), .B1(n41313), .B2(n40143), .C1(
        n40140), .C2(n31183), .ZN(n8427) );
  OAI222_X1 U30213 ( .A1(n40935), .A2(n40150), .B1(n41319), .B2(n40143), .C1(
        n40140), .C2(n31182), .ZN(n8426) );
  OAI222_X1 U30214 ( .A1(n40941), .A2(n40150), .B1(n41325), .B2(n40143), .C1(
        n40140), .C2(n31181), .ZN(n8425) );
  OAI222_X1 U30215 ( .A1(n40947), .A2(n40150), .B1(n41331), .B2(n40143), .C1(
        n40140), .C2(n31180), .ZN(n8424) );
  OAI222_X1 U30216 ( .A1(n40959), .A2(n40150), .B1(n41343), .B2(n40143), .C1(
        n40140), .C2(n31178), .ZN(n8422) );
  OAI222_X1 U30217 ( .A1(n40599), .A2(n40096), .B1(n40983), .B2(n40089), .C1(
        n40077), .C2(n31056), .ZN(n8290) );
  OAI222_X1 U30218 ( .A1(n40605), .A2(n40096), .B1(n40989), .B2(n40089), .C1(
        n40077), .C2(n31055), .ZN(n8289) );
  OAI222_X1 U30219 ( .A1(n40611), .A2(n40096), .B1(n40995), .B2(n40089), .C1(
        n40077), .C2(n31054), .ZN(n8288) );
  OAI222_X1 U30220 ( .A1(n40617), .A2(n40096), .B1(n41001), .B2(n40089), .C1(
        n40077), .C2(n31053), .ZN(n8287) );
  OAI222_X1 U30221 ( .A1(n40623), .A2(n40095), .B1(n41007), .B2(n40088), .C1(
        n40077), .C2(n31052), .ZN(n8286) );
  OAI222_X1 U30222 ( .A1(n40629), .A2(n40095), .B1(n41013), .B2(n40088), .C1(
        n40077), .C2(n31051), .ZN(n8285) );
  OAI222_X1 U30223 ( .A1(n40635), .A2(n40095), .B1(n41019), .B2(n40088), .C1(
        n40077), .C2(n31050), .ZN(n8284) );
  OAI222_X1 U30224 ( .A1(n40641), .A2(n40095), .B1(n41025), .B2(n40088), .C1(
        n40077), .C2(n31049), .ZN(n8283) );
  OAI222_X1 U30225 ( .A1(n40647), .A2(n40095), .B1(n41031), .B2(n40088), .C1(
        n40077), .C2(n31048), .ZN(n8282) );
  OAI222_X1 U30226 ( .A1(n40653), .A2(n40095), .B1(n41037), .B2(n40088), .C1(
        n40077), .C2(n31047), .ZN(n8281) );
  OAI222_X1 U30227 ( .A1(n40659), .A2(n40095), .B1(n41043), .B2(n40088), .C1(
        n40077), .C2(n31046), .ZN(n8280) );
  OAI222_X1 U30228 ( .A1(n40665), .A2(n40095), .B1(n41049), .B2(n40088), .C1(
        n40077), .C2(n31045), .ZN(n8279) );
  OAI222_X1 U30229 ( .A1(n40671), .A2(n40095), .B1(n41055), .B2(n40088), .C1(
        n40078), .C2(n31044), .ZN(n8278) );
  OAI222_X1 U30230 ( .A1(n40677), .A2(n40095), .B1(n41061), .B2(n40088), .C1(
        n40078), .C2(n31043), .ZN(n8277) );
  OAI222_X1 U30231 ( .A1(n40683), .A2(n40095), .B1(n41067), .B2(n40088), .C1(
        n40078), .C2(n31042), .ZN(n8276) );
  OAI222_X1 U30232 ( .A1(n40689), .A2(n40095), .B1(n41073), .B2(n40088), .C1(
        n40079), .C2(n31041), .ZN(n8275) );
  OAI222_X1 U30233 ( .A1(n40695), .A2(n40094), .B1(n41079), .B2(n40087), .C1(
        n40078), .C2(n31040), .ZN(n8274) );
  OAI222_X1 U30234 ( .A1(n40701), .A2(n40094), .B1(n41085), .B2(n40087), .C1(
        n40078), .C2(n31039), .ZN(n8273) );
  OAI222_X1 U30235 ( .A1(n40707), .A2(n40094), .B1(n41091), .B2(n40087), .C1(
        n40078), .C2(n31038), .ZN(n8272) );
  OAI222_X1 U30236 ( .A1(n40713), .A2(n40094), .B1(n41097), .B2(n40087), .C1(
        n40078), .C2(n31037), .ZN(n8271) );
  OAI222_X1 U30237 ( .A1(n40719), .A2(n40094), .B1(n41103), .B2(n40087), .C1(
        n40078), .C2(n31036), .ZN(n8270) );
  OAI222_X1 U30238 ( .A1(n40725), .A2(n40094), .B1(n41109), .B2(n40087), .C1(
        n40078), .C2(n31035), .ZN(n8269) );
  OAI222_X1 U30239 ( .A1(n40731), .A2(n40094), .B1(n41115), .B2(n40087), .C1(
        n40078), .C2(n31034), .ZN(n8268) );
  OAI222_X1 U30240 ( .A1(n40737), .A2(n40094), .B1(n41121), .B2(n40087), .C1(
        n40078), .C2(n31033), .ZN(n8267) );
  OAI222_X1 U30241 ( .A1(n40743), .A2(n40094), .B1(n41127), .B2(n40087), .C1(
        n40078), .C2(n31032), .ZN(n8266) );
  OAI222_X1 U30242 ( .A1(n40749), .A2(n40094), .B1(n41133), .B2(n40087), .C1(
        n40079), .C2(n31031), .ZN(n8265) );
  OAI222_X1 U30243 ( .A1(n40755), .A2(n40094), .B1(n41139), .B2(n40087), .C1(
        n40079), .C2(n31030), .ZN(n8264) );
  OAI222_X1 U30244 ( .A1(n40761), .A2(n40094), .B1(n41145), .B2(n40087), .C1(
        n40079), .C2(n31029), .ZN(n8263) );
  OAI222_X1 U30245 ( .A1(n40767), .A2(n40093), .B1(n41151), .B2(n40086), .C1(
        n40079), .C2(n31028), .ZN(n8262) );
  OAI222_X1 U30246 ( .A1(n40773), .A2(n40093), .B1(n41157), .B2(n40086), .C1(
        n40079), .C2(n31027), .ZN(n8261) );
  OAI222_X1 U30247 ( .A1(n40779), .A2(n40093), .B1(n41163), .B2(n40086), .C1(
        n40079), .C2(n31026), .ZN(n8260) );
  OAI222_X1 U30248 ( .A1(n40785), .A2(n40093), .B1(n41169), .B2(n40086), .C1(
        n40079), .C2(n31025), .ZN(n8259) );
  OAI222_X1 U30249 ( .A1(n40791), .A2(n40093), .B1(n41175), .B2(n40086), .C1(
        n40079), .C2(n31024), .ZN(n8258) );
  OAI222_X1 U30250 ( .A1(n40797), .A2(n40093), .B1(n41181), .B2(n40086), .C1(
        n40079), .C2(n31023), .ZN(n8257) );
  OAI222_X1 U30251 ( .A1(n40803), .A2(n40093), .B1(n41187), .B2(n40086), .C1(
        n40079), .C2(n31022), .ZN(n8256) );
  OAI222_X1 U30252 ( .A1(n40809), .A2(n40093), .B1(n41193), .B2(n40086), .C1(
        n40079), .C2(n31021), .ZN(n8255) );
  OAI222_X1 U30253 ( .A1(n40815), .A2(n40093), .B1(n41199), .B2(n40086), .C1(
        n40080), .C2(n31020), .ZN(n8254) );
  OAI222_X1 U30254 ( .A1(n40821), .A2(n40093), .B1(n41205), .B2(n40086), .C1(
        n40080), .C2(n31019), .ZN(n8253) );
  OAI222_X1 U30255 ( .A1(n40827), .A2(n40093), .B1(n41211), .B2(n40086), .C1(
        n40080), .C2(n31018), .ZN(n8252) );
  OAI222_X1 U30256 ( .A1(n40833), .A2(n40093), .B1(n41217), .B2(n40086), .C1(
        n40080), .C2(n31017), .ZN(n8251) );
  OAI222_X1 U30257 ( .A1(n40839), .A2(n40092), .B1(n41223), .B2(n40085), .C1(
        n40080), .C2(n31016), .ZN(n8250) );
  OAI222_X1 U30258 ( .A1(n40845), .A2(n40092), .B1(n41229), .B2(n40085), .C1(
        n40080), .C2(n31015), .ZN(n8249) );
  OAI222_X1 U30259 ( .A1(n40851), .A2(n40092), .B1(n41235), .B2(n40085), .C1(
        n40080), .C2(n31014), .ZN(n8248) );
  OAI222_X1 U30260 ( .A1(n40857), .A2(n40092), .B1(n41241), .B2(n40085), .C1(
        n40080), .C2(n31013), .ZN(n8247) );
  OAI222_X1 U30261 ( .A1(n40863), .A2(n40092), .B1(n41247), .B2(n40085), .C1(
        n40080), .C2(n31012), .ZN(n8246) );
  OAI222_X1 U30262 ( .A1(n40869), .A2(n40092), .B1(n41253), .B2(n40085), .C1(
        n40080), .C2(n31011), .ZN(n8245) );
  OAI222_X1 U30263 ( .A1(n40875), .A2(n40092), .B1(n41259), .B2(n40085), .C1(
        n40080), .C2(n31010), .ZN(n8244) );
  OAI222_X1 U30264 ( .A1(n40881), .A2(n40092), .B1(n41265), .B2(n40085), .C1(
        n40080), .C2(n31009), .ZN(n8243) );
  OAI222_X1 U30265 ( .A1(n40887), .A2(n40092), .B1(n41271), .B2(n40085), .C1(
        n40081), .C2(n31008), .ZN(n8242) );
  OAI222_X1 U30266 ( .A1(n40893), .A2(n40092), .B1(n41277), .B2(n40085), .C1(
        n40081), .C2(n31007), .ZN(n8241) );
  OAI222_X1 U30267 ( .A1(n40899), .A2(n40092), .B1(n41283), .B2(n40085), .C1(
        n40081), .C2(n31006), .ZN(n8240) );
  OAI222_X1 U30268 ( .A1(n40905), .A2(n40092), .B1(n41289), .B2(n40085), .C1(
        n40081), .C2(n31005), .ZN(n8239) );
  OAI222_X1 U30269 ( .A1(n40911), .A2(n40091), .B1(n41295), .B2(n40084), .C1(
        n40081), .C2(n31004), .ZN(n8238) );
  OAI222_X1 U30270 ( .A1(n40917), .A2(n40091), .B1(n41301), .B2(n40084), .C1(
        n40081), .C2(n31003), .ZN(n8237) );
  OAI222_X1 U30271 ( .A1(n40923), .A2(n40091), .B1(n41307), .B2(n40084), .C1(
        n40081), .C2(n31002), .ZN(n8236) );
  OAI222_X1 U30272 ( .A1(n40929), .A2(n40091), .B1(n41313), .B2(n40084), .C1(
        n40081), .C2(n31001), .ZN(n8235) );
  OAI222_X1 U30273 ( .A1(n40935), .A2(n40091), .B1(n41319), .B2(n40084), .C1(
        n40081), .C2(n31000), .ZN(n8234) );
  OAI222_X1 U30274 ( .A1(n40941), .A2(n40091), .B1(n41325), .B2(n40084), .C1(
        n40081), .C2(n30999), .ZN(n8233) );
  OAI222_X1 U30275 ( .A1(n40947), .A2(n40091), .B1(n41331), .B2(n40084), .C1(
        n40081), .C2(n30998), .ZN(n8232) );
  OAI222_X1 U30276 ( .A1(n40959), .A2(n40091), .B1(n41343), .B2(n40084), .C1(
        n40081), .C2(n30996), .ZN(n8230) );
  OAI222_X1 U30277 ( .A1(n40599), .A2(n40076), .B1(n40983), .B2(n40069), .C1(
        n40057), .C2(n30992), .ZN(n8226) );
  OAI222_X1 U30278 ( .A1(n40605), .A2(n40076), .B1(n40989), .B2(n40069), .C1(
        n40057), .C2(n30991), .ZN(n8225) );
  OAI222_X1 U30279 ( .A1(n40611), .A2(n40076), .B1(n40995), .B2(n40069), .C1(
        n40057), .C2(n30990), .ZN(n8224) );
  OAI222_X1 U30280 ( .A1(n40617), .A2(n40076), .B1(n41001), .B2(n40069), .C1(
        n40057), .C2(n30989), .ZN(n8223) );
  OAI222_X1 U30281 ( .A1(n40623), .A2(n40075), .B1(n41007), .B2(n40068), .C1(
        n40057), .C2(n30988), .ZN(n8222) );
  OAI222_X1 U30282 ( .A1(n40629), .A2(n40075), .B1(n41013), .B2(n40068), .C1(
        n40057), .C2(n30987), .ZN(n8221) );
  OAI222_X1 U30283 ( .A1(n40635), .A2(n40075), .B1(n41019), .B2(n40068), .C1(
        n40057), .C2(n30986), .ZN(n8220) );
  OAI222_X1 U30284 ( .A1(n40641), .A2(n40075), .B1(n41025), .B2(n40068), .C1(
        n40057), .C2(n30985), .ZN(n8219) );
  OAI222_X1 U30285 ( .A1(n40647), .A2(n40075), .B1(n41031), .B2(n40068), .C1(
        n40057), .C2(n30984), .ZN(n8218) );
  OAI222_X1 U30286 ( .A1(n40653), .A2(n40075), .B1(n41037), .B2(n40068), .C1(
        n40057), .C2(n30983), .ZN(n8217) );
  OAI222_X1 U30287 ( .A1(n40659), .A2(n40075), .B1(n41043), .B2(n40068), .C1(
        n40057), .C2(n30982), .ZN(n8216) );
  OAI222_X1 U30288 ( .A1(n40665), .A2(n40075), .B1(n41049), .B2(n40068), .C1(
        n40057), .C2(n30981), .ZN(n8215) );
  OAI222_X1 U30289 ( .A1(n40671), .A2(n40075), .B1(n41055), .B2(n40068), .C1(
        n40058), .C2(n30980), .ZN(n8214) );
  OAI222_X1 U30290 ( .A1(n40677), .A2(n40075), .B1(n41061), .B2(n40068), .C1(
        n40058), .C2(n30979), .ZN(n8213) );
  OAI222_X1 U30291 ( .A1(n40683), .A2(n40075), .B1(n41067), .B2(n40068), .C1(
        n40058), .C2(n30978), .ZN(n8212) );
  OAI222_X1 U30292 ( .A1(n40689), .A2(n40075), .B1(n41073), .B2(n40068), .C1(
        n40059), .C2(n30977), .ZN(n8211) );
  OAI222_X1 U30293 ( .A1(n40695), .A2(n40074), .B1(n41079), .B2(n40067), .C1(
        n40058), .C2(n30976), .ZN(n8210) );
  OAI222_X1 U30294 ( .A1(n40701), .A2(n40074), .B1(n41085), .B2(n40067), .C1(
        n40058), .C2(n30975), .ZN(n8209) );
  OAI222_X1 U30295 ( .A1(n40707), .A2(n40074), .B1(n41091), .B2(n40067), .C1(
        n40058), .C2(n30974), .ZN(n8208) );
  OAI222_X1 U30296 ( .A1(n40713), .A2(n40074), .B1(n41097), .B2(n40067), .C1(
        n40058), .C2(n30973), .ZN(n8207) );
  OAI222_X1 U30297 ( .A1(n40719), .A2(n40074), .B1(n41103), .B2(n40067), .C1(
        n40058), .C2(n30972), .ZN(n8206) );
  OAI222_X1 U30298 ( .A1(n40725), .A2(n40074), .B1(n41109), .B2(n40067), .C1(
        n40058), .C2(n30971), .ZN(n8205) );
  OAI222_X1 U30299 ( .A1(n40731), .A2(n40074), .B1(n41115), .B2(n40067), .C1(
        n40058), .C2(n30970), .ZN(n8204) );
  OAI222_X1 U30300 ( .A1(n40737), .A2(n40074), .B1(n41121), .B2(n40067), .C1(
        n40058), .C2(n30969), .ZN(n8203) );
  OAI222_X1 U30301 ( .A1(n40743), .A2(n40074), .B1(n41127), .B2(n40067), .C1(
        n40058), .C2(n30968), .ZN(n8202) );
  OAI222_X1 U30302 ( .A1(n40749), .A2(n40074), .B1(n41133), .B2(n40067), .C1(
        n40059), .C2(n30967), .ZN(n8201) );
  OAI222_X1 U30303 ( .A1(n40755), .A2(n40074), .B1(n41139), .B2(n40067), .C1(
        n40059), .C2(n30966), .ZN(n8200) );
  OAI222_X1 U30304 ( .A1(n40761), .A2(n40074), .B1(n41145), .B2(n40067), .C1(
        n40059), .C2(n30965), .ZN(n8199) );
  OAI222_X1 U30305 ( .A1(n40767), .A2(n40073), .B1(n41151), .B2(n40066), .C1(
        n40059), .C2(n30964), .ZN(n8198) );
  OAI222_X1 U30306 ( .A1(n40773), .A2(n40073), .B1(n41157), .B2(n40066), .C1(
        n40059), .C2(n30963), .ZN(n8197) );
  OAI222_X1 U30307 ( .A1(n40779), .A2(n40073), .B1(n41163), .B2(n40066), .C1(
        n40059), .C2(n30962), .ZN(n8196) );
  OAI222_X1 U30308 ( .A1(n40785), .A2(n40073), .B1(n41169), .B2(n40066), .C1(
        n40059), .C2(n30961), .ZN(n8195) );
  OAI222_X1 U30309 ( .A1(n40791), .A2(n40073), .B1(n41175), .B2(n40066), .C1(
        n40059), .C2(n30960), .ZN(n8194) );
  OAI222_X1 U30310 ( .A1(n40797), .A2(n40073), .B1(n41181), .B2(n40066), .C1(
        n40059), .C2(n30959), .ZN(n8193) );
  OAI222_X1 U30311 ( .A1(n40803), .A2(n40073), .B1(n41187), .B2(n40066), .C1(
        n40059), .C2(n30958), .ZN(n8192) );
  OAI222_X1 U30312 ( .A1(n40809), .A2(n40073), .B1(n41193), .B2(n40066), .C1(
        n40059), .C2(n30957), .ZN(n8191) );
  OAI222_X1 U30313 ( .A1(n40815), .A2(n40073), .B1(n41199), .B2(n40066), .C1(
        n40060), .C2(n30956), .ZN(n8190) );
  OAI222_X1 U30314 ( .A1(n40821), .A2(n40073), .B1(n41205), .B2(n40066), .C1(
        n40060), .C2(n30955), .ZN(n8189) );
  OAI222_X1 U30315 ( .A1(n40827), .A2(n40073), .B1(n41211), .B2(n40066), .C1(
        n40060), .C2(n30954), .ZN(n8188) );
  OAI222_X1 U30316 ( .A1(n40833), .A2(n40073), .B1(n41217), .B2(n40066), .C1(
        n40060), .C2(n30953), .ZN(n8187) );
  OAI222_X1 U30317 ( .A1(n40839), .A2(n40072), .B1(n41223), .B2(n40065), .C1(
        n40060), .C2(n30952), .ZN(n8186) );
  OAI222_X1 U30318 ( .A1(n40845), .A2(n40072), .B1(n41229), .B2(n40065), .C1(
        n40060), .C2(n30951), .ZN(n8185) );
  OAI222_X1 U30319 ( .A1(n40851), .A2(n40072), .B1(n41235), .B2(n40065), .C1(
        n40060), .C2(n30950), .ZN(n8184) );
  OAI222_X1 U30320 ( .A1(n40857), .A2(n40072), .B1(n41241), .B2(n40065), .C1(
        n40060), .C2(n30949), .ZN(n8183) );
  OAI222_X1 U30321 ( .A1(n40863), .A2(n40072), .B1(n41247), .B2(n40065), .C1(
        n40060), .C2(n30948), .ZN(n8182) );
  OAI222_X1 U30322 ( .A1(n40869), .A2(n40072), .B1(n41253), .B2(n40065), .C1(
        n40060), .C2(n30947), .ZN(n8181) );
  OAI222_X1 U30323 ( .A1(n40875), .A2(n40072), .B1(n41259), .B2(n40065), .C1(
        n40060), .C2(n30946), .ZN(n8180) );
  OAI222_X1 U30324 ( .A1(n40881), .A2(n40072), .B1(n41265), .B2(n40065), .C1(
        n40060), .C2(n30945), .ZN(n8179) );
  OAI222_X1 U30325 ( .A1(n40887), .A2(n40072), .B1(n41271), .B2(n40065), .C1(
        n40061), .C2(n30944), .ZN(n8178) );
  OAI222_X1 U30326 ( .A1(n40893), .A2(n40072), .B1(n41277), .B2(n40065), .C1(
        n40061), .C2(n30943), .ZN(n8177) );
  OAI222_X1 U30327 ( .A1(n40899), .A2(n40072), .B1(n41283), .B2(n40065), .C1(
        n40061), .C2(n30942), .ZN(n8176) );
  OAI222_X1 U30328 ( .A1(n40905), .A2(n40072), .B1(n41289), .B2(n40065), .C1(
        n40061), .C2(n30941), .ZN(n8175) );
  OAI222_X1 U30329 ( .A1(n40911), .A2(n40071), .B1(n41295), .B2(n40064), .C1(
        n40061), .C2(n30940), .ZN(n8174) );
  OAI222_X1 U30330 ( .A1(n40917), .A2(n40071), .B1(n41301), .B2(n40064), .C1(
        n40061), .C2(n30939), .ZN(n8173) );
  OAI222_X1 U30331 ( .A1(n40923), .A2(n40071), .B1(n41307), .B2(n40064), .C1(
        n40061), .C2(n30938), .ZN(n8172) );
  OAI222_X1 U30332 ( .A1(n40929), .A2(n40071), .B1(n41313), .B2(n40064), .C1(
        n40061), .C2(n30937), .ZN(n8171) );
  OAI222_X1 U30333 ( .A1(n40935), .A2(n40071), .B1(n41319), .B2(n40064), .C1(
        n40061), .C2(n30936), .ZN(n8170) );
  OAI222_X1 U30334 ( .A1(n40941), .A2(n40071), .B1(n41325), .B2(n40064), .C1(
        n40061), .C2(n30935), .ZN(n8169) );
  OAI222_X1 U30335 ( .A1(n40947), .A2(n40071), .B1(n41331), .B2(n40064), .C1(
        n40061), .C2(n30934), .ZN(n8168) );
  OAI222_X1 U30336 ( .A1(n40959), .A2(n40071), .B1(n41343), .B2(n40064), .C1(
        n40061), .C2(n30932), .ZN(n8166) );
  OAI222_X1 U30337 ( .A1(n40599), .A2(n40056), .B1(n40983), .B2(n40049), .C1(
        n40037), .C2(n30928), .ZN(n8162) );
  OAI222_X1 U30338 ( .A1(n40605), .A2(n40056), .B1(n40989), .B2(n40049), .C1(
        n40037), .C2(n30927), .ZN(n8161) );
  OAI222_X1 U30339 ( .A1(n40611), .A2(n40056), .B1(n40995), .B2(n40049), .C1(
        n40037), .C2(n30926), .ZN(n8160) );
  OAI222_X1 U30340 ( .A1(n40617), .A2(n40056), .B1(n41001), .B2(n40049), .C1(
        n40037), .C2(n30925), .ZN(n8159) );
  OAI222_X1 U30341 ( .A1(n40623), .A2(n40055), .B1(n41007), .B2(n40048), .C1(
        n40037), .C2(n30924), .ZN(n8158) );
  OAI222_X1 U30342 ( .A1(n40629), .A2(n40055), .B1(n41013), .B2(n40048), .C1(
        n40037), .C2(n30923), .ZN(n8157) );
  OAI222_X1 U30343 ( .A1(n40635), .A2(n40055), .B1(n41019), .B2(n40048), .C1(
        n40037), .C2(n30922), .ZN(n8156) );
  OAI222_X1 U30344 ( .A1(n40641), .A2(n40055), .B1(n41025), .B2(n40048), .C1(
        n40037), .C2(n30921), .ZN(n8155) );
  OAI222_X1 U30345 ( .A1(n40647), .A2(n40055), .B1(n41031), .B2(n40048), .C1(
        n40037), .C2(n30920), .ZN(n8154) );
  OAI222_X1 U30346 ( .A1(n40653), .A2(n40055), .B1(n41037), .B2(n40048), .C1(
        n40037), .C2(n30919), .ZN(n8153) );
  OAI222_X1 U30347 ( .A1(n40659), .A2(n40055), .B1(n41043), .B2(n40048), .C1(
        n40037), .C2(n30918), .ZN(n8152) );
  OAI222_X1 U30348 ( .A1(n40665), .A2(n40055), .B1(n41049), .B2(n40048), .C1(
        n40037), .C2(n30917), .ZN(n8151) );
  OAI222_X1 U30349 ( .A1(n40671), .A2(n40055), .B1(n41055), .B2(n40048), .C1(
        n40038), .C2(n30916), .ZN(n8150) );
  OAI222_X1 U30350 ( .A1(n40677), .A2(n40055), .B1(n41061), .B2(n40048), .C1(
        n40038), .C2(n30915), .ZN(n8149) );
  OAI222_X1 U30351 ( .A1(n40683), .A2(n40055), .B1(n41067), .B2(n40048), .C1(
        n40038), .C2(n30914), .ZN(n8148) );
  OAI222_X1 U30352 ( .A1(n40689), .A2(n40055), .B1(n41073), .B2(n40048), .C1(
        n40039), .C2(n30913), .ZN(n8147) );
  OAI222_X1 U30353 ( .A1(n40695), .A2(n40054), .B1(n41079), .B2(n40047), .C1(
        n40038), .C2(n30912), .ZN(n8146) );
  OAI222_X1 U30354 ( .A1(n40701), .A2(n40054), .B1(n41085), .B2(n40047), .C1(
        n40038), .C2(n30911), .ZN(n8145) );
  OAI222_X1 U30355 ( .A1(n40707), .A2(n40054), .B1(n41091), .B2(n40047), .C1(
        n40038), .C2(n30910), .ZN(n8144) );
  OAI222_X1 U30356 ( .A1(n40713), .A2(n40054), .B1(n41097), .B2(n40047), .C1(
        n40038), .C2(n30909), .ZN(n8143) );
  OAI222_X1 U30357 ( .A1(n40719), .A2(n40054), .B1(n41103), .B2(n40047), .C1(
        n40038), .C2(n30908), .ZN(n8142) );
  OAI222_X1 U30358 ( .A1(n40725), .A2(n40054), .B1(n41109), .B2(n40047), .C1(
        n40038), .C2(n30907), .ZN(n8141) );
  OAI222_X1 U30359 ( .A1(n40731), .A2(n40054), .B1(n41115), .B2(n40047), .C1(
        n40038), .C2(n30906), .ZN(n8140) );
  OAI222_X1 U30360 ( .A1(n40737), .A2(n40054), .B1(n41121), .B2(n40047), .C1(
        n40038), .C2(n30905), .ZN(n8139) );
  OAI222_X1 U30361 ( .A1(n40743), .A2(n40054), .B1(n41127), .B2(n40047), .C1(
        n40038), .C2(n30904), .ZN(n8138) );
  OAI222_X1 U30362 ( .A1(n40749), .A2(n40054), .B1(n41133), .B2(n40047), .C1(
        n40039), .C2(n30903), .ZN(n8137) );
  OAI222_X1 U30363 ( .A1(n40755), .A2(n40054), .B1(n41139), .B2(n40047), .C1(
        n40039), .C2(n30902), .ZN(n8136) );
  OAI222_X1 U30364 ( .A1(n40761), .A2(n40054), .B1(n41145), .B2(n40047), .C1(
        n40039), .C2(n30901), .ZN(n8135) );
  OAI222_X1 U30365 ( .A1(n40767), .A2(n40053), .B1(n41151), .B2(n40046), .C1(
        n40039), .C2(n30900), .ZN(n8134) );
  OAI222_X1 U30366 ( .A1(n40773), .A2(n40053), .B1(n41157), .B2(n40046), .C1(
        n40039), .C2(n30899), .ZN(n8133) );
  OAI222_X1 U30367 ( .A1(n40779), .A2(n40053), .B1(n41163), .B2(n40046), .C1(
        n40039), .C2(n30898), .ZN(n8132) );
  OAI222_X1 U30368 ( .A1(n40785), .A2(n40053), .B1(n41169), .B2(n40046), .C1(
        n40039), .C2(n30897), .ZN(n8131) );
  OAI222_X1 U30369 ( .A1(n40791), .A2(n40053), .B1(n41175), .B2(n40046), .C1(
        n40039), .C2(n30896), .ZN(n8130) );
  OAI222_X1 U30370 ( .A1(n40797), .A2(n40053), .B1(n41181), .B2(n40046), .C1(
        n40039), .C2(n30895), .ZN(n8129) );
  OAI222_X1 U30371 ( .A1(n40803), .A2(n40053), .B1(n41187), .B2(n40046), .C1(
        n40039), .C2(n30894), .ZN(n8128) );
  OAI222_X1 U30372 ( .A1(n40809), .A2(n40053), .B1(n41193), .B2(n40046), .C1(
        n40039), .C2(n30893), .ZN(n8127) );
  OAI222_X1 U30373 ( .A1(n40815), .A2(n40053), .B1(n41199), .B2(n40046), .C1(
        n40040), .C2(n30892), .ZN(n8126) );
  OAI222_X1 U30374 ( .A1(n40821), .A2(n40053), .B1(n41205), .B2(n40046), .C1(
        n40040), .C2(n30891), .ZN(n8125) );
  OAI222_X1 U30375 ( .A1(n40827), .A2(n40053), .B1(n41211), .B2(n40046), .C1(
        n40040), .C2(n30890), .ZN(n8124) );
  OAI222_X1 U30376 ( .A1(n40833), .A2(n40053), .B1(n41217), .B2(n40046), .C1(
        n40040), .C2(n30889), .ZN(n8123) );
  OAI222_X1 U30377 ( .A1(n40839), .A2(n40052), .B1(n41223), .B2(n40045), .C1(
        n40040), .C2(n30888), .ZN(n8122) );
  OAI222_X1 U30378 ( .A1(n40845), .A2(n40052), .B1(n41229), .B2(n40045), .C1(
        n40040), .C2(n30887), .ZN(n8121) );
  OAI222_X1 U30379 ( .A1(n40851), .A2(n40052), .B1(n41235), .B2(n40045), .C1(
        n40040), .C2(n30886), .ZN(n8120) );
  OAI222_X1 U30380 ( .A1(n40857), .A2(n40052), .B1(n41241), .B2(n40045), .C1(
        n40040), .C2(n30885), .ZN(n8119) );
  OAI222_X1 U30381 ( .A1(n40863), .A2(n40052), .B1(n41247), .B2(n40045), .C1(
        n40040), .C2(n30884), .ZN(n8118) );
  OAI222_X1 U30382 ( .A1(n40869), .A2(n40052), .B1(n41253), .B2(n40045), .C1(
        n40040), .C2(n30883), .ZN(n8117) );
  OAI222_X1 U30383 ( .A1(n40875), .A2(n40052), .B1(n41259), .B2(n40045), .C1(
        n40040), .C2(n30882), .ZN(n8116) );
  OAI222_X1 U30384 ( .A1(n40881), .A2(n40052), .B1(n41265), .B2(n40045), .C1(
        n40040), .C2(n30881), .ZN(n8115) );
  OAI222_X1 U30385 ( .A1(n40887), .A2(n40052), .B1(n41271), .B2(n40045), .C1(
        n40041), .C2(n30880), .ZN(n8114) );
  OAI222_X1 U30386 ( .A1(n40893), .A2(n40052), .B1(n41277), .B2(n40045), .C1(
        n40041), .C2(n30879), .ZN(n8113) );
  OAI222_X1 U30387 ( .A1(n40899), .A2(n40052), .B1(n41283), .B2(n40045), .C1(
        n40041), .C2(n30878), .ZN(n8112) );
  OAI222_X1 U30388 ( .A1(n40905), .A2(n40052), .B1(n41289), .B2(n40045), .C1(
        n40041), .C2(n30877), .ZN(n8111) );
  OAI222_X1 U30389 ( .A1(n40911), .A2(n40051), .B1(n41295), .B2(n40044), .C1(
        n40041), .C2(n30876), .ZN(n8110) );
  OAI222_X1 U30390 ( .A1(n40917), .A2(n40051), .B1(n41301), .B2(n40044), .C1(
        n40041), .C2(n30875), .ZN(n8109) );
  OAI222_X1 U30391 ( .A1(n40923), .A2(n40051), .B1(n41307), .B2(n40044), .C1(
        n40041), .C2(n30874), .ZN(n8108) );
  OAI222_X1 U30392 ( .A1(n40929), .A2(n40051), .B1(n41313), .B2(n40044), .C1(
        n40041), .C2(n30873), .ZN(n8107) );
  OAI222_X1 U30393 ( .A1(n40935), .A2(n40051), .B1(n41319), .B2(n40044), .C1(
        n40041), .C2(n30872), .ZN(n8106) );
  OAI222_X1 U30394 ( .A1(n40941), .A2(n40051), .B1(n41325), .B2(n40044), .C1(
        n40041), .C2(n30871), .ZN(n8105) );
  OAI222_X1 U30395 ( .A1(n40947), .A2(n40051), .B1(n41331), .B2(n40044), .C1(
        n40041), .C2(n30870), .ZN(n8104) );
  OAI222_X1 U30396 ( .A1(n40959), .A2(n40051), .B1(n41343), .B2(n40044), .C1(
        n40041), .C2(n30868), .ZN(n8102) );
  OAI222_X1 U30397 ( .A1(n40598), .A2(n39998), .B1(n40982), .B2(n39991), .C1(
        n39979), .C2(n30864), .ZN(n7970) );
  OAI222_X1 U30398 ( .A1(n40604), .A2(n39998), .B1(n40988), .B2(n39991), .C1(
        n39979), .C2(n30863), .ZN(n7969) );
  OAI222_X1 U30399 ( .A1(n40610), .A2(n39998), .B1(n40994), .B2(n39991), .C1(
        n39979), .C2(n30862), .ZN(n7968) );
  OAI222_X1 U30400 ( .A1(n40616), .A2(n39998), .B1(n41000), .B2(n39991), .C1(
        n39979), .C2(n30861), .ZN(n7967) );
  OAI222_X1 U30401 ( .A1(n40622), .A2(n39997), .B1(n41006), .B2(n39990), .C1(
        n39979), .C2(n30860), .ZN(n7966) );
  OAI222_X1 U30402 ( .A1(n40628), .A2(n39997), .B1(n41012), .B2(n39990), .C1(
        n39979), .C2(n30859), .ZN(n7965) );
  OAI222_X1 U30403 ( .A1(n40634), .A2(n39997), .B1(n41018), .B2(n39990), .C1(
        n39979), .C2(n30858), .ZN(n7964) );
  OAI222_X1 U30404 ( .A1(n40640), .A2(n39997), .B1(n41024), .B2(n39990), .C1(
        n39979), .C2(n30857), .ZN(n7963) );
  OAI222_X1 U30405 ( .A1(n40646), .A2(n39997), .B1(n41030), .B2(n39990), .C1(
        n39979), .C2(n30856), .ZN(n7962) );
  OAI222_X1 U30406 ( .A1(n40652), .A2(n39997), .B1(n41036), .B2(n39990), .C1(
        n39979), .C2(n30855), .ZN(n7961) );
  OAI222_X1 U30407 ( .A1(n40658), .A2(n39997), .B1(n41042), .B2(n39990), .C1(
        n39979), .C2(n30854), .ZN(n7960) );
  OAI222_X1 U30408 ( .A1(n40664), .A2(n39997), .B1(n41048), .B2(n39990), .C1(
        n39979), .C2(n30853), .ZN(n7959) );
  OAI222_X1 U30409 ( .A1(n40670), .A2(n39997), .B1(n41054), .B2(n39990), .C1(
        n39980), .C2(n30852), .ZN(n7958) );
  OAI222_X1 U30410 ( .A1(n40676), .A2(n39997), .B1(n41060), .B2(n39990), .C1(
        n39980), .C2(n30851), .ZN(n7957) );
  OAI222_X1 U30411 ( .A1(n40682), .A2(n39997), .B1(n41066), .B2(n39990), .C1(
        n39980), .C2(n30850), .ZN(n7956) );
  OAI222_X1 U30412 ( .A1(n40688), .A2(n39997), .B1(n41072), .B2(n39990), .C1(
        n39981), .C2(n30849), .ZN(n7955) );
  OAI222_X1 U30413 ( .A1(n40694), .A2(n39996), .B1(n41078), .B2(n39989), .C1(
        n39980), .C2(n30848), .ZN(n7954) );
  OAI222_X1 U30414 ( .A1(n40700), .A2(n39996), .B1(n41084), .B2(n39989), .C1(
        n39980), .C2(n30847), .ZN(n7953) );
  OAI222_X1 U30415 ( .A1(n40706), .A2(n39996), .B1(n41090), .B2(n39989), .C1(
        n39980), .C2(n30846), .ZN(n7952) );
  OAI222_X1 U30416 ( .A1(n40712), .A2(n39996), .B1(n41096), .B2(n39989), .C1(
        n39980), .C2(n30845), .ZN(n7951) );
  OAI222_X1 U30417 ( .A1(n40718), .A2(n39996), .B1(n41102), .B2(n39989), .C1(
        n39980), .C2(n30844), .ZN(n7950) );
  OAI222_X1 U30418 ( .A1(n40724), .A2(n39996), .B1(n41108), .B2(n39989), .C1(
        n39980), .C2(n30843), .ZN(n7949) );
  OAI222_X1 U30419 ( .A1(n40730), .A2(n39996), .B1(n41114), .B2(n39989), .C1(
        n39980), .C2(n30842), .ZN(n7948) );
  OAI222_X1 U30420 ( .A1(n40736), .A2(n39996), .B1(n41120), .B2(n39989), .C1(
        n39980), .C2(n30841), .ZN(n7947) );
  OAI222_X1 U30421 ( .A1(n40742), .A2(n39996), .B1(n41126), .B2(n39989), .C1(
        n39980), .C2(n30840), .ZN(n7946) );
  OAI222_X1 U30422 ( .A1(n40748), .A2(n39996), .B1(n41132), .B2(n39989), .C1(
        n39981), .C2(n30839), .ZN(n7945) );
  OAI222_X1 U30423 ( .A1(n40754), .A2(n39996), .B1(n41138), .B2(n39989), .C1(
        n39981), .C2(n30838), .ZN(n7944) );
  OAI222_X1 U30424 ( .A1(n40760), .A2(n39996), .B1(n41144), .B2(n39989), .C1(
        n39981), .C2(n30837), .ZN(n7943) );
  OAI222_X1 U30425 ( .A1(n40766), .A2(n39995), .B1(n41150), .B2(n39988), .C1(
        n39981), .C2(n30836), .ZN(n7942) );
  OAI222_X1 U30426 ( .A1(n40772), .A2(n39995), .B1(n41156), .B2(n39988), .C1(
        n39981), .C2(n30835), .ZN(n7941) );
  OAI222_X1 U30427 ( .A1(n40778), .A2(n39995), .B1(n41162), .B2(n39988), .C1(
        n39981), .C2(n30834), .ZN(n7940) );
  OAI222_X1 U30428 ( .A1(n40784), .A2(n39995), .B1(n41168), .B2(n39988), .C1(
        n39981), .C2(n30833), .ZN(n7939) );
  OAI222_X1 U30429 ( .A1(n40790), .A2(n39995), .B1(n41174), .B2(n39988), .C1(
        n39981), .C2(n30832), .ZN(n7938) );
  OAI222_X1 U30430 ( .A1(n40796), .A2(n39995), .B1(n41180), .B2(n39988), .C1(
        n39981), .C2(n30831), .ZN(n7937) );
  OAI222_X1 U30431 ( .A1(n40802), .A2(n39995), .B1(n41186), .B2(n39988), .C1(
        n39981), .C2(n30830), .ZN(n7936) );
  OAI222_X1 U30432 ( .A1(n40808), .A2(n39995), .B1(n41192), .B2(n39988), .C1(
        n39981), .C2(n30829), .ZN(n7935) );
  OAI222_X1 U30433 ( .A1(n40814), .A2(n39995), .B1(n41198), .B2(n39988), .C1(
        n39982), .C2(n30828), .ZN(n7934) );
  OAI222_X1 U30434 ( .A1(n40820), .A2(n39995), .B1(n41204), .B2(n39988), .C1(
        n39982), .C2(n30827), .ZN(n7933) );
  OAI222_X1 U30435 ( .A1(n40826), .A2(n39995), .B1(n41210), .B2(n39988), .C1(
        n39982), .C2(n30826), .ZN(n7932) );
  OAI222_X1 U30436 ( .A1(n40832), .A2(n39995), .B1(n41216), .B2(n39988), .C1(
        n39982), .C2(n30825), .ZN(n7931) );
  OAI222_X1 U30437 ( .A1(n40838), .A2(n39994), .B1(n41222), .B2(n39987), .C1(
        n39982), .C2(n30824), .ZN(n7930) );
  OAI222_X1 U30438 ( .A1(n40844), .A2(n39994), .B1(n41228), .B2(n39987), .C1(
        n39982), .C2(n30823), .ZN(n7929) );
  OAI222_X1 U30439 ( .A1(n40850), .A2(n39994), .B1(n41234), .B2(n39987), .C1(
        n39982), .C2(n30822), .ZN(n7928) );
  OAI222_X1 U30440 ( .A1(n40856), .A2(n39994), .B1(n41240), .B2(n39987), .C1(
        n39982), .C2(n30821), .ZN(n7927) );
  OAI222_X1 U30441 ( .A1(n40862), .A2(n39994), .B1(n41246), .B2(n39987), .C1(
        n39982), .C2(n30820), .ZN(n7926) );
  OAI222_X1 U30442 ( .A1(n40868), .A2(n39994), .B1(n41252), .B2(n39987), .C1(
        n39982), .C2(n30819), .ZN(n7925) );
  OAI222_X1 U30443 ( .A1(n40874), .A2(n39994), .B1(n41258), .B2(n39987), .C1(
        n39982), .C2(n30818), .ZN(n7924) );
  OAI222_X1 U30444 ( .A1(n40880), .A2(n39994), .B1(n41264), .B2(n39987), .C1(
        n39982), .C2(n30817), .ZN(n7923) );
  OAI222_X1 U30445 ( .A1(n40886), .A2(n39994), .B1(n41270), .B2(n39987), .C1(
        n39983), .C2(n30816), .ZN(n7922) );
  OAI222_X1 U30446 ( .A1(n40892), .A2(n39994), .B1(n41276), .B2(n39987), .C1(
        n39983), .C2(n30815), .ZN(n7921) );
  OAI222_X1 U30447 ( .A1(n40898), .A2(n39994), .B1(n41282), .B2(n39987), .C1(
        n39983), .C2(n30814), .ZN(n7920) );
  OAI222_X1 U30448 ( .A1(n40904), .A2(n39994), .B1(n41288), .B2(n39987), .C1(
        n39983), .C2(n30813), .ZN(n7919) );
  OAI222_X1 U30449 ( .A1(n40910), .A2(n39993), .B1(n41294), .B2(n39986), .C1(
        n39983), .C2(n30812), .ZN(n7918) );
  OAI222_X1 U30450 ( .A1(n40916), .A2(n39993), .B1(n41300), .B2(n39986), .C1(
        n39983), .C2(n30811), .ZN(n7917) );
  OAI222_X1 U30451 ( .A1(n40922), .A2(n39993), .B1(n41306), .B2(n39986), .C1(
        n39983), .C2(n30810), .ZN(n7916) );
  OAI222_X1 U30452 ( .A1(n40928), .A2(n39993), .B1(n41312), .B2(n39986), .C1(
        n39983), .C2(n30809), .ZN(n7915) );
  OAI222_X1 U30453 ( .A1(n40934), .A2(n39993), .B1(n41318), .B2(n39986), .C1(
        n39983), .C2(n30808), .ZN(n7914) );
  OAI222_X1 U30454 ( .A1(n40940), .A2(n39993), .B1(n41324), .B2(n39986), .C1(
        n39983), .C2(n30807), .ZN(n7913) );
  OAI222_X1 U30455 ( .A1(n40946), .A2(n39993), .B1(n41330), .B2(n39986), .C1(
        n39983), .C2(n30806), .ZN(n7912) );
  OAI222_X1 U30456 ( .A1(n40958), .A2(n39993), .B1(n41342), .B2(n39986), .C1(
        n39983), .C2(n30804), .ZN(n7910) );
  OAI222_X1 U30457 ( .A1(n40598), .A2(n39978), .B1(n40982), .B2(n39971), .C1(
        n39959), .C2(n30800), .ZN(n7906) );
  OAI222_X1 U30458 ( .A1(n40604), .A2(n39978), .B1(n40988), .B2(n39971), .C1(
        n39959), .C2(n30799), .ZN(n7905) );
  OAI222_X1 U30459 ( .A1(n40610), .A2(n39978), .B1(n40994), .B2(n39971), .C1(
        n39959), .C2(n30798), .ZN(n7904) );
  OAI222_X1 U30460 ( .A1(n40616), .A2(n39978), .B1(n41000), .B2(n39971), .C1(
        n39959), .C2(n30797), .ZN(n7903) );
  OAI222_X1 U30461 ( .A1(n40622), .A2(n39977), .B1(n41006), .B2(n39970), .C1(
        n39959), .C2(n30796), .ZN(n7902) );
  OAI222_X1 U30462 ( .A1(n40628), .A2(n39977), .B1(n41012), .B2(n39970), .C1(
        n39959), .C2(n30795), .ZN(n7901) );
  OAI222_X1 U30463 ( .A1(n40634), .A2(n39977), .B1(n41018), .B2(n39970), .C1(
        n39959), .C2(n30794), .ZN(n7900) );
  OAI222_X1 U30464 ( .A1(n40640), .A2(n39977), .B1(n41024), .B2(n39970), .C1(
        n39959), .C2(n30793), .ZN(n7899) );
  OAI222_X1 U30465 ( .A1(n40646), .A2(n39977), .B1(n41030), .B2(n39970), .C1(
        n39959), .C2(n30792), .ZN(n7898) );
  OAI222_X1 U30466 ( .A1(n40652), .A2(n39977), .B1(n41036), .B2(n39970), .C1(
        n39959), .C2(n30791), .ZN(n7897) );
  OAI222_X1 U30467 ( .A1(n40658), .A2(n39977), .B1(n41042), .B2(n39970), .C1(
        n39959), .C2(n30790), .ZN(n7896) );
  OAI222_X1 U30468 ( .A1(n40664), .A2(n39977), .B1(n41048), .B2(n39970), .C1(
        n39959), .C2(n30789), .ZN(n7895) );
  OAI222_X1 U30469 ( .A1(n40670), .A2(n39977), .B1(n41054), .B2(n39970), .C1(
        n39960), .C2(n30788), .ZN(n7894) );
  OAI222_X1 U30470 ( .A1(n40676), .A2(n39977), .B1(n41060), .B2(n39970), .C1(
        n39960), .C2(n30787), .ZN(n7893) );
  OAI222_X1 U30471 ( .A1(n40682), .A2(n39977), .B1(n41066), .B2(n39970), .C1(
        n39960), .C2(n30786), .ZN(n7892) );
  OAI222_X1 U30472 ( .A1(n40688), .A2(n39977), .B1(n41072), .B2(n39970), .C1(
        n39961), .C2(n30785), .ZN(n7891) );
  OAI222_X1 U30473 ( .A1(n40694), .A2(n39976), .B1(n41078), .B2(n39969), .C1(
        n39960), .C2(n30784), .ZN(n7890) );
  OAI222_X1 U30474 ( .A1(n40700), .A2(n39976), .B1(n41084), .B2(n39969), .C1(
        n39960), .C2(n30783), .ZN(n7889) );
  OAI222_X1 U30475 ( .A1(n40706), .A2(n39976), .B1(n41090), .B2(n39969), .C1(
        n39960), .C2(n30782), .ZN(n7888) );
  OAI222_X1 U30476 ( .A1(n40712), .A2(n39976), .B1(n41096), .B2(n39969), .C1(
        n39960), .C2(n30781), .ZN(n7887) );
  OAI222_X1 U30477 ( .A1(n40718), .A2(n39976), .B1(n41102), .B2(n39969), .C1(
        n39960), .C2(n30780), .ZN(n7886) );
  OAI222_X1 U30478 ( .A1(n40724), .A2(n39976), .B1(n41108), .B2(n39969), .C1(
        n39960), .C2(n30779), .ZN(n7885) );
  OAI222_X1 U30479 ( .A1(n40730), .A2(n39976), .B1(n41114), .B2(n39969), .C1(
        n39960), .C2(n30778), .ZN(n7884) );
  OAI222_X1 U30480 ( .A1(n40736), .A2(n39976), .B1(n41120), .B2(n39969), .C1(
        n39960), .C2(n30777), .ZN(n7883) );
  OAI222_X1 U30481 ( .A1(n40742), .A2(n39976), .B1(n41126), .B2(n39969), .C1(
        n39960), .C2(n30776), .ZN(n7882) );
  OAI222_X1 U30482 ( .A1(n40748), .A2(n39976), .B1(n41132), .B2(n39969), .C1(
        n39961), .C2(n30775), .ZN(n7881) );
  OAI222_X1 U30483 ( .A1(n40754), .A2(n39976), .B1(n41138), .B2(n39969), .C1(
        n39961), .C2(n30774), .ZN(n7880) );
  OAI222_X1 U30484 ( .A1(n40760), .A2(n39976), .B1(n41144), .B2(n39969), .C1(
        n39961), .C2(n30773), .ZN(n7879) );
  OAI222_X1 U30485 ( .A1(n40766), .A2(n39975), .B1(n41150), .B2(n39968), .C1(
        n39961), .C2(n30772), .ZN(n7878) );
  OAI222_X1 U30486 ( .A1(n40772), .A2(n39975), .B1(n41156), .B2(n39968), .C1(
        n39961), .C2(n30771), .ZN(n7877) );
  OAI222_X1 U30487 ( .A1(n40778), .A2(n39975), .B1(n41162), .B2(n39968), .C1(
        n39961), .C2(n30770), .ZN(n7876) );
  OAI222_X1 U30488 ( .A1(n40784), .A2(n39975), .B1(n41168), .B2(n39968), .C1(
        n39961), .C2(n30769), .ZN(n7875) );
  OAI222_X1 U30489 ( .A1(n40790), .A2(n39975), .B1(n41174), .B2(n39968), .C1(
        n39961), .C2(n30768), .ZN(n7874) );
  OAI222_X1 U30490 ( .A1(n40796), .A2(n39975), .B1(n41180), .B2(n39968), .C1(
        n39961), .C2(n30767), .ZN(n7873) );
  OAI222_X1 U30491 ( .A1(n40802), .A2(n39975), .B1(n41186), .B2(n39968), .C1(
        n39961), .C2(n30766), .ZN(n7872) );
  OAI222_X1 U30492 ( .A1(n40808), .A2(n39975), .B1(n41192), .B2(n39968), .C1(
        n39961), .C2(n30765), .ZN(n7871) );
  OAI222_X1 U30493 ( .A1(n40814), .A2(n39975), .B1(n41198), .B2(n39968), .C1(
        n39962), .C2(n30764), .ZN(n7870) );
  OAI222_X1 U30494 ( .A1(n40820), .A2(n39975), .B1(n41204), .B2(n39968), .C1(
        n39962), .C2(n30763), .ZN(n7869) );
  OAI222_X1 U30495 ( .A1(n40826), .A2(n39975), .B1(n41210), .B2(n39968), .C1(
        n39962), .C2(n30762), .ZN(n7868) );
  OAI222_X1 U30496 ( .A1(n40832), .A2(n39975), .B1(n41216), .B2(n39968), .C1(
        n39962), .C2(n30761), .ZN(n7867) );
  OAI222_X1 U30497 ( .A1(n40838), .A2(n39974), .B1(n41222), .B2(n39967), .C1(
        n39962), .C2(n30760), .ZN(n7866) );
  OAI222_X1 U30498 ( .A1(n40844), .A2(n39974), .B1(n41228), .B2(n39967), .C1(
        n39962), .C2(n30759), .ZN(n7865) );
  OAI222_X1 U30499 ( .A1(n40850), .A2(n39974), .B1(n41234), .B2(n39967), .C1(
        n39962), .C2(n30758), .ZN(n7864) );
  OAI222_X1 U30500 ( .A1(n40856), .A2(n39974), .B1(n41240), .B2(n39967), .C1(
        n39962), .C2(n30757), .ZN(n7863) );
  OAI222_X1 U30501 ( .A1(n40862), .A2(n39974), .B1(n41246), .B2(n39967), .C1(
        n39962), .C2(n30756), .ZN(n7862) );
  OAI222_X1 U30502 ( .A1(n40868), .A2(n39974), .B1(n41252), .B2(n39967), .C1(
        n39962), .C2(n30755), .ZN(n7861) );
  OAI222_X1 U30503 ( .A1(n40874), .A2(n39974), .B1(n41258), .B2(n39967), .C1(
        n39962), .C2(n30754), .ZN(n7860) );
  OAI222_X1 U30504 ( .A1(n40880), .A2(n39974), .B1(n41264), .B2(n39967), .C1(
        n39962), .C2(n30753), .ZN(n7859) );
  OAI222_X1 U30505 ( .A1(n40886), .A2(n39974), .B1(n41270), .B2(n39967), .C1(
        n39963), .C2(n30752), .ZN(n7858) );
  OAI222_X1 U30506 ( .A1(n40892), .A2(n39974), .B1(n41276), .B2(n39967), .C1(
        n39963), .C2(n30751), .ZN(n7857) );
  OAI222_X1 U30507 ( .A1(n40898), .A2(n39974), .B1(n41282), .B2(n39967), .C1(
        n39963), .C2(n30750), .ZN(n7856) );
  OAI222_X1 U30508 ( .A1(n40904), .A2(n39974), .B1(n41288), .B2(n39967), .C1(
        n39963), .C2(n30749), .ZN(n7855) );
  OAI222_X1 U30509 ( .A1(n40910), .A2(n39973), .B1(n41294), .B2(n39966), .C1(
        n39963), .C2(n30748), .ZN(n7854) );
  OAI222_X1 U30510 ( .A1(n40916), .A2(n39973), .B1(n41300), .B2(n39966), .C1(
        n39963), .C2(n30747), .ZN(n7853) );
  OAI222_X1 U30511 ( .A1(n40922), .A2(n39973), .B1(n41306), .B2(n39966), .C1(
        n39963), .C2(n30746), .ZN(n7852) );
  OAI222_X1 U30512 ( .A1(n40928), .A2(n39973), .B1(n41312), .B2(n39966), .C1(
        n39963), .C2(n30745), .ZN(n7851) );
  OAI222_X1 U30513 ( .A1(n40934), .A2(n39973), .B1(n41318), .B2(n39966), .C1(
        n39963), .C2(n30744), .ZN(n7850) );
  OAI222_X1 U30514 ( .A1(n40940), .A2(n39973), .B1(n41324), .B2(n39966), .C1(
        n39963), .C2(n30743), .ZN(n7849) );
  OAI222_X1 U30515 ( .A1(n40946), .A2(n39973), .B1(n41330), .B2(n39966), .C1(
        n39963), .C2(n30742), .ZN(n7848) );
  OAI222_X1 U30516 ( .A1(n40958), .A2(n39973), .B1(n41342), .B2(n39966), .C1(
        n39963), .C2(n30740), .ZN(n7846) );
  OAI222_X1 U30517 ( .A1(n40598), .A2(n39958), .B1(n40982), .B2(n39951), .C1(
        n39939), .C2(n30736), .ZN(n7842) );
  OAI222_X1 U30518 ( .A1(n40604), .A2(n39958), .B1(n40988), .B2(n39951), .C1(
        n39939), .C2(n30735), .ZN(n7841) );
  OAI222_X1 U30519 ( .A1(n40610), .A2(n39958), .B1(n40994), .B2(n39951), .C1(
        n39939), .C2(n30734), .ZN(n7840) );
  OAI222_X1 U30520 ( .A1(n40616), .A2(n39958), .B1(n41000), .B2(n39951), .C1(
        n39939), .C2(n30733), .ZN(n7839) );
  OAI222_X1 U30521 ( .A1(n40622), .A2(n39957), .B1(n41006), .B2(n39950), .C1(
        n39939), .C2(n30732), .ZN(n7838) );
  OAI222_X1 U30522 ( .A1(n40628), .A2(n39957), .B1(n41012), .B2(n39950), .C1(
        n39939), .C2(n30731), .ZN(n7837) );
  OAI222_X1 U30523 ( .A1(n40634), .A2(n39957), .B1(n41018), .B2(n39950), .C1(
        n39939), .C2(n30730), .ZN(n7836) );
  OAI222_X1 U30524 ( .A1(n40640), .A2(n39957), .B1(n41024), .B2(n39950), .C1(
        n39939), .C2(n30729), .ZN(n7835) );
  OAI222_X1 U30525 ( .A1(n40646), .A2(n39957), .B1(n41030), .B2(n39950), .C1(
        n39939), .C2(n30728), .ZN(n7834) );
  OAI222_X1 U30526 ( .A1(n40652), .A2(n39957), .B1(n41036), .B2(n39950), .C1(
        n39939), .C2(n30727), .ZN(n7833) );
  OAI222_X1 U30527 ( .A1(n40658), .A2(n39957), .B1(n41042), .B2(n39950), .C1(
        n39939), .C2(n30726), .ZN(n7832) );
  OAI222_X1 U30528 ( .A1(n40664), .A2(n39957), .B1(n41048), .B2(n39950), .C1(
        n39939), .C2(n30725), .ZN(n7831) );
  OAI222_X1 U30529 ( .A1(n40670), .A2(n39957), .B1(n41054), .B2(n39950), .C1(
        n39940), .C2(n30724), .ZN(n7830) );
  OAI222_X1 U30530 ( .A1(n40676), .A2(n39957), .B1(n41060), .B2(n39950), .C1(
        n39940), .C2(n30723), .ZN(n7829) );
  OAI222_X1 U30531 ( .A1(n40682), .A2(n39957), .B1(n41066), .B2(n39950), .C1(
        n39940), .C2(n30722), .ZN(n7828) );
  OAI222_X1 U30532 ( .A1(n40688), .A2(n39957), .B1(n41072), .B2(n39950), .C1(
        n39941), .C2(n30721), .ZN(n7827) );
  OAI222_X1 U30533 ( .A1(n40694), .A2(n39956), .B1(n41078), .B2(n39949), .C1(
        n39940), .C2(n30720), .ZN(n7826) );
  OAI222_X1 U30534 ( .A1(n40700), .A2(n39956), .B1(n41084), .B2(n39949), .C1(
        n39940), .C2(n30719), .ZN(n7825) );
  OAI222_X1 U30535 ( .A1(n40706), .A2(n39956), .B1(n41090), .B2(n39949), .C1(
        n39940), .C2(n30718), .ZN(n7824) );
  OAI222_X1 U30536 ( .A1(n40712), .A2(n39956), .B1(n41096), .B2(n39949), .C1(
        n39940), .C2(n30717), .ZN(n7823) );
  OAI222_X1 U30537 ( .A1(n40718), .A2(n39956), .B1(n41102), .B2(n39949), .C1(
        n39940), .C2(n30716), .ZN(n7822) );
  OAI222_X1 U30538 ( .A1(n40724), .A2(n39956), .B1(n41108), .B2(n39949), .C1(
        n39940), .C2(n30715), .ZN(n7821) );
  OAI222_X1 U30539 ( .A1(n40730), .A2(n39956), .B1(n41114), .B2(n39949), .C1(
        n39940), .C2(n30714), .ZN(n7820) );
  OAI222_X1 U30540 ( .A1(n40736), .A2(n39956), .B1(n41120), .B2(n39949), .C1(
        n39940), .C2(n30713), .ZN(n7819) );
  OAI222_X1 U30541 ( .A1(n40742), .A2(n39956), .B1(n41126), .B2(n39949), .C1(
        n39940), .C2(n30712), .ZN(n7818) );
  OAI222_X1 U30542 ( .A1(n40748), .A2(n39956), .B1(n41132), .B2(n39949), .C1(
        n39941), .C2(n30711), .ZN(n7817) );
  OAI222_X1 U30543 ( .A1(n40754), .A2(n39956), .B1(n41138), .B2(n39949), .C1(
        n39941), .C2(n30710), .ZN(n7816) );
  OAI222_X1 U30544 ( .A1(n40760), .A2(n39956), .B1(n41144), .B2(n39949), .C1(
        n39941), .C2(n30709), .ZN(n7815) );
  OAI222_X1 U30545 ( .A1(n40766), .A2(n39955), .B1(n41150), .B2(n39948), .C1(
        n39941), .C2(n30708), .ZN(n7814) );
  OAI222_X1 U30546 ( .A1(n40772), .A2(n39955), .B1(n41156), .B2(n39948), .C1(
        n39941), .C2(n30707), .ZN(n7813) );
  OAI222_X1 U30547 ( .A1(n40778), .A2(n39955), .B1(n41162), .B2(n39948), .C1(
        n39941), .C2(n30706), .ZN(n7812) );
  OAI222_X1 U30548 ( .A1(n40784), .A2(n39955), .B1(n41168), .B2(n39948), .C1(
        n39941), .C2(n30705), .ZN(n7811) );
  OAI222_X1 U30549 ( .A1(n40790), .A2(n39955), .B1(n41174), .B2(n39948), .C1(
        n39941), .C2(n30704), .ZN(n7810) );
  OAI222_X1 U30550 ( .A1(n40796), .A2(n39955), .B1(n41180), .B2(n39948), .C1(
        n39941), .C2(n30703), .ZN(n7809) );
  OAI222_X1 U30551 ( .A1(n40802), .A2(n39955), .B1(n41186), .B2(n39948), .C1(
        n39941), .C2(n30702), .ZN(n7808) );
  OAI222_X1 U30552 ( .A1(n40808), .A2(n39955), .B1(n41192), .B2(n39948), .C1(
        n39941), .C2(n30701), .ZN(n7807) );
  OAI222_X1 U30553 ( .A1(n40814), .A2(n39955), .B1(n41198), .B2(n39948), .C1(
        n39942), .C2(n30700), .ZN(n7806) );
  OAI222_X1 U30554 ( .A1(n40820), .A2(n39955), .B1(n41204), .B2(n39948), .C1(
        n39942), .C2(n30699), .ZN(n7805) );
  OAI222_X1 U30555 ( .A1(n40826), .A2(n39955), .B1(n41210), .B2(n39948), .C1(
        n39942), .C2(n30698), .ZN(n7804) );
  OAI222_X1 U30556 ( .A1(n40832), .A2(n39955), .B1(n41216), .B2(n39948), .C1(
        n39942), .C2(n30697), .ZN(n7803) );
  OAI222_X1 U30557 ( .A1(n40838), .A2(n39954), .B1(n41222), .B2(n39947), .C1(
        n39942), .C2(n30696), .ZN(n7802) );
  OAI222_X1 U30558 ( .A1(n40844), .A2(n39954), .B1(n41228), .B2(n39947), .C1(
        n39942), .C2(n30695), .ZN(n7801) );
  OAI222_X1 U30559 ( .A1(n40850), .A2(n39954), .B1(n41234), .B2(n39947), .C1(
        n39942), .C2(n30694), .ZN(n7800) );
  OAI222_X1 U30560 ( .A1(n40856), .A2(n39954), .B1(n41240), .B2(n39947), .C1(
        n39942), .C2(n30693), .ZN(n7799) );
  OAI222_X1 U30561 ( .A1(n40862), .A2(n39954), .B1(n41246), .B2(n39947), .C1(
        n39942), .C2(n30692), .ZN(n7798) );
  OAI222_X1 U30562 ( .A1(n40868), .A2(n39954), .B1(n41252), .B2(n39947), .C1(
        n39942), .C2(n30691), .ZN(n7797) );
  OAI222_X1 U30563 ( .A1(n40874), .A2(n39954), .B1(n41258), .B2(n39947), .C1(
        n39942), .C2(n30690), .ZN(n7796) );
  OAI222_X1 U30564 ( .A1(n40880), .A2(n39954), .B1(n41264), .B2(n39947), .C1(
        n39942), .C2(n30689), .ZN(n7795) );
  OAI222_X1 U30565 ( .A1(n40886), .A2(n39954), .B1(n41270), .B2(n39947), .C1(
        n39943), .C2(n30688), .ZN(n7794) );
  OAI222_X1 U30566 ( .A1(n40892), .A2(n39954), .B1(n41276), .B2(n39947), .C1(
        n39943), .C2(n30687), .ZN(n7793) );
  OAI222_X1 U30567 ( .A1(n40898), .A2(n39954), .B1(n41282), .B2(n39947), .C1(
        n39943), .C2(n30686), .ZN(n7792) );
  OAI222_X1 U30568 ( .A1(n40904), .A2(n39954), .B1(n41288), .B2(n39947), .C1(
        n39943), .C2(n30685), .ZN(n7791) );
  OAI222_X1 U30569 ( .A1(n40910), .A2(n39953), .B1(n41294), .B2(n39946), .C1(
        n39943), .C2(n30684), .ZN(n7790) );
  OAI222_X1 U30570 ( .A1(n40916), .A2(n39953), .B1(n41300), .B2(n39946), .C1(
        n39943), .C2(n30683), .ZN(n7789) );
  OAI222_X1 U30571 ( .A1(n40922), .A2(n39953), .B1(n41306), .B2(n39946), .C1(
        n39943), .C2(n30682), .ZN(n7788) );
  OAI222_X1 U30572 ( .A1(n40928), .A2(n39953), .B1(n41312), .B2(n39946), .C1(
        n39943), .C2(n30681), .ZN(n7787) );
  OAI222_X1 U30573 ( .A1(n40934), .A2(n39953), .B1(n41318), .B2(n39946), .C1(
        n39943), .C2(n30680), .ZN(n7786) );
  OAI222_X1 U30574 ( .A1(n40940), .A2(n39953), .B1(n41324), .B2(n39946), .C1(
        n39943), .C2(n30679), .ZN(n7785) );
  OAI222_X1 U30575 ( .A1(n40946), .A2(n39953), .B1(n41330), .B2(n39946), .C1(
        n39943), .C2(n30678), .ZN(n7784) );
  OAI222_X1 U30576 ( .A1(n40958), .A2(n39953), .B1(n41342), .B2(n39946), .C1(
        n39943), .C2(n30676), .ZN(n7782) );
  OAI222_X1 U30577 ( .A1(n40598), .A2(n39900), .B1(n40982), .B2(n39893), .C1(
        n39881), .C2(n30672), .ZN(n7650) );
  OAI222_X1 U30578 ( .A1(n40604), .A2(n39900), .B1(n40988), .B2(n39893), .C1(
        n39881), .C2(n30671), .ZN(n7649) );
  OAI222_X1 U30579 ( .A1(n40610), .A2(n39900), .B1(n40994), .B2(n39893), .C1(
        n39881), .C2(n30670), .ZN(n7648) );
  OAI222_X1 U30580 ( .A1(n40616), .A2(n39900), .B1(n41000), .B2(n39893), .C1(
        n39881), .C2(n30669), .ZN(n7647) );
  OAI222_X1 U30581 ( .A1(n40622), .A2(n39899), .B1(n41006), .B2(n39892), .C1(
        n39881), .C2(n30668), .ZN(n7646) );
  OAI222_X1 U30582 ( .A1(n40628), .A2(n39899), .B1(n41012), .B2(n39892), .C1(
        n39881), .C2(n30667), .ZN(n7645) );
  OAI222_X1 U30583 ( .A1(n40634), .A2(n39899), .B1(n41018), .B2(n39892), .C1(
        n39881), .C2(n30666), .ZN(n7644) );
  OAI222_X1 U30584 ( .A1(n40640), .A2(n39899), .B1(n41024), .B2(n39892), .C1(
        n39881), .C2(n30665), .ZN(n7643) );
  OAI222_X1 U30585 ( .A1(n40646), .A2(n39899), .B1(n41030), .B2(n39892), .C1(
        n39881), .C2(n30664), .ZN(n7642) );
  OAI222_X1 U30586 ( .A1(n40652), .A2(n39899), .B1(n41036), .B2(n39892), .C1(
        n39881), .C2(n30663), .ZN(n7641) );
  OAI222_X1 U30587 ( .A1(n40658), .A2(n39899), .B1(n41042), .B2(n39892), .C1(
        n39881), .C2(n30662), .ZN(n7640) );
  OAI222_X1 U30588 ( .A1(n40664), .A2(n39899), .B1(n41048), .B2(n39892), .C1(
        n39881), .C2(n30661), .ZN(n7639) );
  OAI222_X1 U30589 ( .A1(n40670), .A2(n39899), .B1(n41054), .B2(n39892), .C1(
        n39882), .C2(n30660), .ZN(n7638) );
  OAI222_X1 U30590 ( .A1(n40676), .A2(n39899), .B1(n41060), .B2(n39892), .C1(
        n39882), .C2(n30659), .ZN(n7637) );
  OAI222_X1 U30591 ( .A1(n40682), .A2(n39899), .B1(n41066), .B2(n39892), .C1(
        n39882), .C2(n30658), .ZN(n7636) );
  OAI222_X1 U30592 ( .A1(n40688), .A2(n39899), .B1(n41072), .B2(n39892), .C1(
        n39883), .C2(n30657), .ZN(n7635) );
  OAI222_X1 U30593 ( .A1(n40694), .A2(n39898), .B1(n41078), .B2(n39891), .C1(
        n39882), .C2(n30656), .ZN(n7634) );
  OAI222_X1 U30594 ( .A1(n40700), .A2(n39898), .B1(n41084), .B2(n39891), .C1(
        n39882), .C2(n30655), .ZN(n7633) );
  OAI222_X1 U30595 ( .A1(n40706), .A2(n39898), .B1(n41090), .B2(n39891), .C1(
        n39882), .C2(n30654), .ZN(n7632) );
  OAI222_X1 U30596 ( .A1(n40712), .A2(n39898), .B1(n41096), .B2(n39891), .C1(
        n39882), .C2(n30653), .ZN(n7631) );
  OAI222_X1 U30597 ( .A1(n40718), .A2(n39898), .B1(n41102), .B2(n39891), .C1(
        n39882), .C2(n30652), .ZN(n7630) );
  OAI222_X1 U30598 ( .A1(n40724), .A2(n39898), .B1(n41108), .B2(n39891), .C1(
        n39882), .C2(n30651), .ZN(n7629) );
  OAI222_X1 U30599 ( .A1(n40730), .A2(n39898), .B1(n41114), .B2(n39891), .C1(
        n39882), .C2(n30650), .ZN(n7628) );
  OAI222_X1 U30600 ( .A1(n40736), .A2(n39898), .B1(n41120), .B2(n39891), .C1(
        n39882), .C2(n30649), .ZN(n7627) );
  OAI222_X1 U30601 ( .A1(n40742), .A2(n39898), .B1(n41126), .B2(n39891), .C1(
        n39882), .C2(n30648), .ZN(n7626) );
  OAI222_X1 U30602 ( .A1(n40748), .A2(n39898), .B1(n41132), .B2(n39891), .C1(
        n39883), .C2(n30647), .ZN(n7625) );
  OAI222_X1 U30603 ( .A1(n40754), .A2(n39898), .B1(n41138), .B2(n39891), .C1(
        n39883), .C2(n30646), .ZN(n7624) );
  OAI222_X1 U30604 ( .A1(n40760), .A2(n39898), .B1(n41144), .B2(n39891), .C1(
        n39883), .C2(n30645), .ZN(n7623) );
  OAI222_X1 U30605 ( .A1(n40766), .A2(n39897), .B1(n41150), .B2(n39890), .C1(
        n39883), .C2(n30644), .ZN(n7622) );
  OAI222_X1 U30606 ( .A1(n40772), .A2(n39897), .B1(n41156), .B2(n39890), .C1(
        n39883), .C2(n30643), .ZN(n7621) );
  OAI222_X1 U30607 ( .A1(n40778), .A2(n39897), .B1(n41162), .B2(n39890), .C1(
        n39883), .C2(n30642), .ZN(n7620) );
  OAI222_X1 U30608 ( .A1(n40784), .A2(n39897), .B1(n41168), .B2(n39890), .C1(
        n39883), .C2(n30641), .ZN(n7619) );
  OAI222_X1 U30609 ( .A1(n40790), .A2(n39897), .B1(n41174), .B2(n39890), .C1(
        n39883), .C2(n30640), .ZN(n7618) );
  OAI222_X1 U30610 ( .A1(n40796), .A2(n39897), .B1(n41180), .B2(n39890), .C1(
        n39883), .C2(n30639), .ZN(n7617) );
  OAI222_X1 U30611 ( .A1(n40802), .A2(n39897), .B1(n41186), .B2(n39890), .C1(
        n39883), .C2(n30638), .ZN(n7616) );
  OAI222_X1 U30612 ( .A1(n40808), .A2(n39897), .B1(n41192), .B2(n39890), .C1(
        n39883), .C2(n30637), .ZN(n7615) );
  OAI222_X1 U30613 ( .A1(n40814), .A2(n39897), .B1(n41198), .B2(n39890), .C1(
        n39884), .C2(n30636), .ZN(n7614) );
  OAI222_X1 U30614 ( .A1(n40820), .A2(n39897), .B1(n41204), .B2(n39890), .C1(
        n39884), .C2(n30635), .ZN(n7613) );
  OAI222_X1 U30615 ( .A1(n40826), .A2(n39897), .B1(n41210), .B2(n39890), .C1(
        n39884), .C2(n30634), .ZN(n7612) );
  OAI222_X1 U30616 ( .A1(n40832), .A2(n39897), .B1(n41216), .B2(n39890), .C1(
        n39884), .C2(n30633), .ZN(n7611) );
  OAI222_X1 U30617 ( .A1(n40838), .A2(n39896), .B1(n41222), .B2(n39889), .C1(
        n39884), .C2(n30632), .ZN(n7610) );
  OAI222_X1 U30618 ( .A1(n40844), .A2(n39896), .B1(n41228), .B2(n39889), .C1(
        n39884), .C2(n30631), .ZN(n7609) );
  OAI222_X1 U30619 ( .A1(n40850), .A2(n39896), .B1(n41234), .B2(n39889), .C1(
        n39884), .C2(n30630), .ZN(n7608) );
  OAI222_X1 U30620 ( .A1(n40856), .A2(n39896), .B1(n41240), .B2(n39889), .C1(
        n39884), .C2(n30629), .ZN(n7607) );
  OAI222_X1 U30621 ( .A1(n40862), .A2(n39896), .B1(n41246), .B2(n39889), .C1(
        n39884), .C2(n30628), .ZN(n7606) );
  OAI222_X1 U30622 ( .A1(n40868), .A2(n39896), .B1(n41252), .B2(n39889), .C1(
        n39884), .C2(n30627), .ZN(n7605) );
  OAI222_X1 U30623 ( .A1(n40874), .A2(n39896), .B1(n41258), .B2(n39889), .C1(
        n39884), .C2(n30626), .ZN(n7604) );
  OAI222_X1 U30624 ( .A1(n40880), .A2(n39896), .B1(n41264), .B2(n39889), .C1(
        n39884), .C2(n30625), .ZN(n7603) );
  OAI222_X1 U30625 ( .A1(n40886), .A2(n39896), .B1(n41270), .B2(n39889), .C1(
        n39885), .C2(n30624), .ZN(n7602) );
  OAI222_X1 U30626 ( .A1(n40892), .A2(n39896), .B1(n41276), .B2(n39889), .C1(
        n39885), .C2(n30623), .ZN(n7601) );
  OAI222_X1 U30627 ( .A1(n40898), .A2(n39896), .B1(n41282), .B2(n39889), .C1(
        n39885), .C2(n30622), .ZN(n7600) );
  OAI222_X1 U30628 ( .A1(n40904), .A2(n39896), .B1(n41288), .B2(n39889), .C1(
        n39885), .C2(n30621), .ZN(n7599) );
  OAI222_X1 U30629 ( .A1(n40910), .A2(n39895), .B1(n41294), .B2(n39888), .C1(
        n39885), .C2(n30620), .ZN(n7598) );
  OAI222_X1 U30630 ( .A1(n40916), .A2(n39895), .B1(n41300), .B2(n39888), .C1(
        n39885), .C2(n30619), .ZN(n7597) );
  OAI222_X1 U30631 ( .A1(n40922), .A2(n39895), .B1(n41306), .B2(n39888), .C1(
        n39885), .C2(n30618), .ZN(n7596) );
  OAI222_X1 U30632 ( .A1(n40928), .A2(n39895), .B1(n41312), .B2(n39888), .C1(
        n39885), .C2(n30617), .ZN(n7595) );
  OAI222_X1 U30633 ( .A1(n40934), .A2(n39895), .B1(n41318), .B2(n39888), .C1(
        n39885), .C2(n30616), .ZN(n7594) );
  OAI222_X1 U30634 ( .A1(n40940), .A2(n39895), .B1(n41324), .B2(n39888), .C1(
        n39885), .C2(n30615), .ZN(n7593) );
  OAI222_X1 U30635 ( .A1(n40946), .A2(n39895), .B1(n41330), .B2(n39888), .C1(
        n39885), .C2(n30614), .ZN(n7592) );
  OAI222_X1 U30636 ( .A1(n40958), .A2(n39895), .B1(n41342), .B2(n39888), .C1(
        n39885), .C2(n30612), .ZN(n7590) );
  OAI222_X1 U30637 ( .A1(n40598), .A2(n39880), .B1(n40982), .B2(n39873), .C1(
        n39861), .C2(n30608), .ZN(n7586) );
  OAI222_X1 U30638 ( .A1(n40604), .A2(n39880), .B1(n40988), .B2(n39873), .C1(
        n39861), .C2(n30607), .ZN(n7585) );
  OAI222_X1 U30639 ( .A1(n40610), .A2(n39880), .B1(n40994), .B2(n39873), .C1(
        n39861), .C2(n30606), .ZN(n7584) );
  OAI222_X1 U30640 ( .A1(n40616), .A2(n39880), .B1(n41000), .B2(n39873), .C1(
        n39861), .C2(n30605), .ZN(n7583) );
  OAI222_X1 U30641 ( .A1(n40622), .A2(n39879), .B1(n41006), .B2(n39872), .C1(
        n39861), .C2(n30604), .ZN(n7582) );
  OAI222_X1 U30642 ( .A1(n40628), .A2(n39879), .B1(n41012), .B2(n39872), .C1(
        n39861), .C2(n30603), .ZN(n7581) );
  OAI222_X1 U30643 ( .A1(n40634), .A2(n39879), .B1(n41018), .B2(n39872), .C1(
        n39861), .C2(n30602), .ZN(n7580) );
  OAI222_X1 U30644 ( .A1(n40640), .A2(n39879), .B1(n41024), .B2(n39872), .C1(
        n39861), .C2(n30601), .ZN(n7579) );
  OAI222_X1 U30645 ( .A1(n40646), .A2(n39879), .B1(n41030), .B2(n39872), .C1(
        n39861), .C2(n30600), .ZN(n7578) );
  OAI222_X1 U30646 ( .A1(n40652), .A2(n39879), .B1(n41036), .B2(n39872), .C1(
        n39861), .C2(n30599), .ZN(n7577) );
  OAI222_X1 U30647 ( .A1(n40658), .A2(n39879), .B1(n41042), .B2(n39872), .C1(
        n39861), .C2(n30598), .ZN(n7576) );
  OAI222_X1 U30648 ( .A1(n40664), .A2(n39879), .B1(n41048), .B2(n39872), .C1(
        n39861), .C2(n30597), .ZN(n7575) );
  OAI222_X1 U30649 ( .A1(n40670), .A2(n39879), .B1(n41054), .B2(n39872), .C1(
        n39862), .C2(n30596), .ZN(n7574) );
  OAI222_X1 U30650 ( .A1(n40676), .A2(n39879), .B1(n41060), .B2(n39872), .C1(
        n39862), .C2(n30595), .ZN(n7573) );
  OAI222_X1 U30651 ( .A1(n40682), .A2(n39879), .B1(n41066), .B2(n39872), .C1(
        n39862), .C2(n30594), .ZN(n7572) );
  OAI222_X1 U30652 ( .A1(n40688), .A2(n39879), .B1(n41072), .B2(n39872), .C1(
        n39863), .C2(n30593), .ZN(n7571) );
  OAI222_X1 U30653 ( .A1(n40694), .A2(n39878), .B1(n41078), .B2(n39871), .C1(
        n39862), .C2(n30592), .ZN(n7570) );
  OAI222_X1 U30654 ( .A1(n40700), .A2(n39878), .B1(n41084), .B2(n39871), .C1(
        n39862), .C2(n30591), .ZN(n7569) );
  OAI222_X1 U30655 ( .A1(n40706), .A2(n39878), .B1(n41090), .B2(n39871), .C1(
        n39862), .C2(n30590), .ZN(n7568) );
  OAI222_X1 U30656 ( .A1(n40712), .A2(n39878), .B1(n41096), .B2(n39871), .C1(
        n39862), .C2(n30589), .ZN(n7567) );
  OAI222_X1 U30657 ( .A1(n40718), .A2(n39878), .B1(n41102), .B2(n39871), .C1(
        n39862), .C2(n30588), .ZN(n7566) );
  OAI222_X1 U30658 ( .A1(n40724), .A2(n39878), .B1(n41108), .B2(n39871), .C1(
        n39862), .C2(n30587), .ZN(n7565) );
  OAI222_X1 U30659 ( .A1(n40730), .A2(n39878), .B1(n41114), .B2(n39871), .C1(
        n39862), .C2(n30586), .ZN(n7564) );
  OAI222_X1 U30660 ( .A1(n40736), .A2(n39878), .B1(n41120), .B2(n39871), .C1(
        n39862), .C2(n30585), .ZN(n7563) );
  OAI222_X1 U30661 ( .A1(n40742), .A2(n39878), .B1(n41126), .B2(n39871), .C1(
        n39862), .C2(n30584), .ZN(n7562) );
  OAI222_X1 U30662 ( .A1(n40748), .A2(n39878), .B1(n41132), .B2(n39871), .C1(
        n39863), .C2(n30583), .ZN(n7561) );
  OAI222_X1 U30663 ( .A1(n40754), .A2(n39878), .B1(n41138), .B2(n39871), .C1(
        n39863), .C2(n30582), .ZN(n7560) );
  OAI222_X1 U30664 ( .A1(n40760), .A2(n39878), .B1(n41144), .B2(n39871), .C1(
        n39863), .C2(n30581), .ZN(n7559) );
  OAI222_X1 U30665 ( .A1(n40766), .A2(n39877), .B1(n41150), .B2(n39870), .C1(
        n39863), .C2(n30580), .ZN(n7558) );
  OAI222_X1 U30666 ( .A1(n40772), .A2(n39877), .B1(n41156), .B2(n39870), .C1(
        n39863), .C2(n30579), .ZN(n7557) );
  OAI222_X1 U30667 ( .A1(n40778), .A2(n39877), .B1(n41162), .B2(n39870), .C1(
        n39863), .C2(n30578), .ZN(n7556) );
  OAI222_X1 U30668 ( .A1(n40784), .A2(n39877), .B1(n41168), .B2(n39870), .C1(
        n39863), .C2(n30577), .ZN(n7555) );
  OAI222_X1 U30669 ( .A1(n40790), .A2(n39877), .B1(n41174), .B2(n39870), .C1(
        n39863), .C2(n30576), .ZN(n7554) );
  OAI222_X1 U30670 ( .A1(n40796), .A2(n39877), .B1(n41180), .B2(n39870), .C1(
        n39863), .C2(n30575), .ZN(n7553) );
  OAI222_X1 U30671 ( .A1(n40802), .A2(n39877), .B1(n41186), .B2(n39870), .C1(
        n39863), .C2(n30574), .ZN(n7552) );
  OAI222_X1 U30672 ( .A1(n40808), .A2(n39877), .B1(n41192), .B2(n39870), .C1(
        n39863), .C2(n30573), .ZN(n7551) );
  OAI222_X1 U30673 ( .A1(n40814), .A2(n39877), .B1(n41198), .B2(n39870), .C1(
        n39864), .C2(n30572), .ZN(n7550) );
  OAI222_X1 U30674 ( .A1(n40820), .A2(n39877), .B1(n41204), .B2(n39870), .C1(
        n39864), .C2(n30571), .ZN(n7549) );
  OAI222_X1 U30675 ( .A1(n40826), .A2(n39877), .B1(n41210), .B2(n39870), .C1(
        n39864), .C2(n30570), .ZN(n7548) );
  OAI222_X1 U30676 ( .A1(n40832), .A2(n39877), .B1(n41216), .B2(n39870), .C1(
        n39864), .C2(n30569), .ZN(n7547) );
  OAI222_X1 U30677 ( .A1(n40838), .A2(n39876), .B1(n41222), .B2(n39869), .C1(
        n39864), .C2(n30568), .ZN(n7546) );
  OAI222_X1 U30678 ( .A1(n40844), .A2(n39876), .B1(n41228), .B2(n39869), .C1(
        n39864), .C2(n30567), .ZN(n7545) );
  OAI222_X1 U30679 ( .A1(n40850), .A2(n39876), .B1(n41234), .B2(n39869), .C1(
        n39864), .C2(n30566), .ZN(n7544) );
  OAI222_X1 U30680 ( .A1(n40856), .A2(n39876), .B1(n41240), .B2(n39869), .C1(
        n39864), .C2(n30565), .ZN(n7543) );
  OAI222_X1 U30681 ( .A1(n40862), .A2(n39876), .B1(n41246), .B2(n39869), .C1(
        n39864), .C2(n30564), .ZN(n7542) );
  OAI222_X1 U30682 ( .A1(n40868), .A2(n39876), .B1(n41252), .B2(n39869), .C1(
        n39864), .C2(n30563), .ZN(n7541) );
  OAI222_X1 U30683 ( .A1(n40874), .A2(n39876), .B1(n41258), .B2(n39869), .C1(
        n39864), .C2(n30562), .ZN(n7540) );
  OAI222_X1 U30684 ( .A1(n40880), .A2(n39876), .B1(n41264), .B2(n39869), .C1(
        n39864), .C2(n30561), .ZN(n7539) );
  OAI222_X1 U30685 ( .A1(n40886), .A2(n39876), .B1(n41270), .B2(n39869), .C1(
        n39865), .C2(n30560), .ZN(n7538) );
  OAI222_X1 U30686 ( .A1(n40892), .A2(n39876), .B1(n41276), .B2(n39869), .C1(
        n39865), .C2(n30559), .ZN(n7537) );
  OAI222_X1 U30687 ( .A1(n40898), .A2(n39876), .B1(n41282), .B2(n39869), .C1(
        n39865), .C2(n30558), .ZN(n7536) );
  OAI222_X1 U30688 ( .A1(n40904), .A2(n39876), .B1(n41288), .B2(n39869), .C1(
        n39865), .C2(n30557), .ZN(n7535) );
  OAI222_X1 U30689 ( .A1(n40910), .A2(n39875), .B1(n41294), .B2(n39868), .C1(
        n39865), .C2(n30556), .ZN(n7534) );
  OAI222_X1 U30690 ( .A1(n40916), .A2(n39875), .B1(n41300), .B2(n39868), .C1(
        n39865), .C2(n30555), .ZN(n7533) );
  OAI222_X1 U30691 ( .A1(n40922), .A2(n39875), .B1(n41306), .B2(n39868), .C1(
        n39865), .C2(n30554), .ZN(n7532) );
  OAI222_X1 U30692 ( .A1(n40928), .A2(n39875), .B1(n41312), .B2(n39868), .C1(
        n39865), .C2(n30553), .ZN(n7531) );
  OAI222_X1 U30693 ( .A1(n40934), .A2(n39875), .B1(n41318), .B2(n39868), .C1(
        n39865), .C2(n30552), .ZN(n7530) );
  OAI222_X1 U30694 ( .A1(n40940), .A2(n39875), .B1(n41324), .B2(n39868), .C1(
        n39865), .C2(n30551), .ZN(n7529) );
  OAI222_X1 U30695 ( .A1(n40946), .A2(n39875), .B1(n41330), .B2(n39868), .C1(
        n39865), .C2(n30550), .ZN(n7528) );
  OAI222_X1 U30696 ( .A1(n40958), .A2(n39875), .B1(n41342), .B2(n39868), .C1(
        n39865), .C2(n30548), .ZN(n7526) );
  OAI222_X1 U30697 ( .A1(n40598), .A2(n39860), .B1(n40982), .B2(n39853), .C1(
        n39841), .C2(n30544), .ZN(n7522) );
  OAI222_X1 U30698 ( .A1(n40604), .A2(n39860), .B1(n40988), .B2(n39853), .C1(
        n39841), .C2(n30543), .ZN(n7521) );
  OAI222_X1 U30699 ( .A1(n40610), .A2(n39860), .B1(n40994), .B2(n39853), .C1(
        n39841), .C2(n30542), .ZN(n7520) );
  OAI222_X1 U30700 ( .A1(n40616), .A2(n39860), .B1(n41000), .B2(n39853), .C1(
        n39841), .C2(n30541), .ZN(n7519) );
  OAI222_X1 U30701 ( .A1(n40622), .A2(n39859), .B1(n41006), .B2(n39852), .C1(
        n39841), .C2(n30540), .ZN(n7518) );
  OAI222_X1 U30702 ( .A1(n40628), .A2(n39859), .B1(n41012), .B2(n39852), .C1(
        n39841), .C2(n30539), .ZN(n7517) );
  OAI222_X1 U30703 ( .A1(n40634), .A2(n39859), .B1(n41018), .B2(n39852), .C1(
        n39841), .C2(n30538), .ZN(n7516) );
  OAI222_X1 U30704 ( .A1(n40640), .A2(n39859), .B1(n41024), .B2(n39852), .C1(
        n39841), .C2(n30537), .ZN(n7515) );
  OAI222_X1 U30705 ( .A1(n40646), .A2(n39859), .B1(n41030), .B2(n39852), .C1(
        n39841), .C2(n30536), .ZN(n7514) );
  OAI222_X1 U30706 ( .A1(n40652), .A2(n39859), .B1(n41036), .B2(n39852), .C1(
        n39841), .C2(n30535), .ZN(n7513) );
  OAI222_X1 U30707 ( .A1(n40658), .A2(n39859), .B1(n41042), .B2(n39852), .C1(
        n39841), .C2(n30534), .ZN(n7512) );
  OAI222_X1 U30708 ( .A1(n40664), .A2(n39859), .B1(n41048), .B2(n39852), .C1(
        n39841), .C2(n30533), .ZN(n7511) );
  OAI222_X1 U30709 ( .A1(n40670), .A2(n39859), .B1(n41054), .B2(n39852), .C1(
        n39842), .C2(n30532), .ZN(n7510) );
  OAI222_X1 U30710 ( .A1(n40676), .A2(n39859), .B1(n41060), .B2(n39852), .C1(
        n39842), .C2(n30531), .ZN(n7509) );
  OAI222_X1 U30711 ( .A1(n40682), .A2(n39859), .B1(n41066), .B2(n39852), .C1(
        n39842), .C2(n30530), .ZN(n7508) );
  OAI222_X1 U30712 ( .A1(n40688), .A2(n39859), .B1(n41072), .B2(n39852), .C1(
        n39843), .C2(n30529), .ZN(n7507) );
  OAI222_X1 U30713 ( .A1(n40694), .A2(n39858), .B1(n41078), .B2(n39851), .C1(
        n39842), .C2(n30528), .ZN(n7506) );
  OAI222_X1 U30714 ( .A1(n40700), .A2(n39858), .B1(n41084), .B2(n39851), .C1(
        n39842), .C2(n30527), .ZN(n7505) );
  OAI222_X1 U30715 ( .A1(n40706), .A2(n39858), .B1(n41090), .B2(n39851), .C1(
        n39842), .C2(n30526), .ZN(n7504) );
  OAI222_X1 U30716 ( .A1(n40712), .A2(n39858), .B1(n41096), .B2(n39851), .C1(
        n39842), .C2(n30525), .ZN(n7503) );
  OAI222_X1 U30717 ( .A1(n40718), .A2(n39858), .B1(n41102), .B2(n39851), .C1(
        n39842), .C2(n30524), .ZN(n7502) );
  OAI222_X1 U30718 ( .A1(n40724), .A2(n39858), .B1(n41108), .B2(n39851), .C1(
        n39842), .C2(n30523), .ZN(n7501) );
  OAI222_X1 U30719 ( .A1(n40730), .A2(n39858), .B1(n41114), .B2(n39851), .C1(
        n39842), .C2(n30522), .ZN(n7500) );
  OAI222_X1 U30720 ( .A1(n40736), .A2(n39858), .B1(n41120), .B2(n39851), .C1(
        n39842), .C2(n30521), .ZN(n7499) );
  OAI222_X1 U30721 ( .A1(n40742), .A2(n39858), .B1(n41126), .B2(n39851), .C1(
        n39842), .C2(n30520), .ZN(n7498) );
  OAI222_X1 U30722 ( .A1(n40748), .A2(n39858), .B1(n41132), .B2(n39851), .C1(
        n39843), .C2(n30519), .ZN(n7497) );
  OAI222_X1 U30723 ( .A1(n40754), .A2(n39858), .B1(n41138), .B2(n39851), .C1(
        n39843), .C2(n30518), .ZN(n7496) );
  OAI222_X1 U30724 ( .A1(n40760), .A2(n39858), .B1(n41144), .B2(n39851), .C1(
        n39843), .C2(n30517), .ZN(n7495) );
  OAI222_X1 U30725 ( .A1(n40766), .A2(n39857), .B1(n41150), .B2(n39850), .C1(
        n39843), .C2(n30516), .ZN(n7494) );
  OAI222_X1 U30726 ( .A1(n40772), .A2(n39857), .B1(n41156), .B2(n39850), .C1(
        n39843), .C2(n30515), .ZN(n7493) );
  OAI222_X1 U30727 ( .A1(n40778), .A2(n39857), .B1(n41162), .B2(n39850), .C1(
        n39843), .C2(n30514), .ZN(n7492) );
  OAI222_X1 U30728 ( .A1(n40784), .A2(n39857), .B1(n41168), .B2(n39850), .C1(
        n39843), .C2(n30513), .ZN(n7491) );
  OAI222_X1 U30729 ( .A1(n40790), .A2(n39857), .B1(n41174), .B2(n39850), .C1(
        n39843), .C2(n30512), .ZN(n7490) );
  OAI222_X1 U30730 ( .A1(n40796), .A2(n39857), .B1(n41180), .B2(n39850), .C1(
        n39843), .C2(n30511), .ZN(n7489) );
  OAI222_X1 U30731 ( .A1(n40802), .A2(n39857), .B1(n41186), .B2(n39850), .C1(
        n39843), .C2(n30510), .ZN(n7488) );
  OAI222_X1 U30732 ( .A1(n40808), .A2(n39857), .B1(n41192), .B2(n39850), .C1(
        n39843), .C2(n30509), .ZN(n7487) );
  OAI222_X1 U30733 ( .A1(n40814), .A2(n39857), .B1(n41198), .B2(n39850), .C1(
        n39844), .C2(n30508), .ZN(n7486) );
  OAI222_X1 U30734 ( .A1(n40820), .A2(n39857), .B1(n41204), .B2(n39850), .C1(
        n39844), .C2(n30507), .ZN(n7485) );
  OAI222_X1 U30735 ( .A1(n40826), .A2(n39857), .B1(n41210), .B2(n39850), .C1(
        n39844), .C2(n30506), .ZN(n7484) );
  OAI222_X1 U30736 ( .A1(n40832), .A2(n39857), .B1(n41216), .B2(n39850), .C1(
        n39844), .C2(n30505), .ZN(n7483) );
  OAI222_X1 U30737 ( .A1(n40838), .A2(n39856), .B1(n41222), .B2(n39849), .C1(
        n39844), .C2(n30504), .ZN(n7482) );
  OAI222_X1 U30738 ( .A1(n40844), .A2(n39856), .B1(n41228), .B2(n39849), .C1(
        n39844), .C2(n30503), .ZN(n7481) );
  OAI222_X1 U30739 ( .A1(n40850), .A2(n39856), .B1(n41234), .B2(n39849), .C1(
        n39844), .C2(n30502), .ZN(n7480) );
  OAI222_X1 U30740 ( .A1(n40856), .A2(n39856), .B1(n41240), .B2(n39849), .C1(
        n39844), .C2(n30501), .ZN(n7479) );
  OAI222_X1 U30741 ( .A1(n40862), .A2(n39856), .B1(n41246), .B2(n39849), .C1(
        n39844), .C2(n30500), .ZN(n7478) );
  OAI222_X1 U30742 ( .A1(n40868), .A2(n39856), .B1(n41252), .B2(n39849), .C1(
        n39844), .C2(n30499), .ZN(n7477) );
  OAI222_X1 U30743 ( .A1(n40874), .A2(n39856), .B1(n41258), .B2(n39849), .C1(
        n39844), .C2(n30498), .ZN(n7476) );
  OAI222_X1 U30744 ( .A1(n40880), .A2(n39856), .B1(n41264), .B2(n39849), .C1(
        n39844), .C2(n30497), .ZN(n7475) );
  OAI222_X1 U30745 ( .A1(n40886), .A2(n39856), .B1(n41270), .B2(n39849), .C1(
        n39845), .C2(n30496), .ZN(n7474) );
  OAI222_X1 U30746 ( .A1(n40892), .A2(n39856), .B1(n41276), .B2(n39849), .C1(
        n39845), .C2(n30495), .ZN(n7473) );
  OAI222_X1 U30747 ( .A1(n40898), .A2(n39856), .B1(n41282), .B2(n39849), .C1(
        n39845), .C2(n30494), .ZN(n7472) );
  OAI222_X1 U30748 ( .A1(n40904), .A2(n39856), .B1(n41288), .B2(n39849), .C1(
        n39845), .C2(n30493), .ZN(n7471) );
  OAI222_X1 U30749 ( .A1(n40910), .A2(n39855), .B1(n41294), .B2(n39848), .C1(
        n39845), .C2(n30492), .ZN(n7470) );
  OAI222_X1 U30750 ( .A1(n40916), .A2(n39855), .B1(n41300), .B2(n39848), .C1(
        n39845), .C2(n30491), .ZN(n7469) );
  OAI222_X1 U30751 ( .A1(n40922), .A2(n39855), .B1(n41306), .B2(n39848), .C1(
        n39845), .C2(n30490), .ZN(n7468) );
  OAI222_X1 U30752 ( .A1(n40928), .A2(n39855), .B1(n41312), .B2(n39848), .C1(
        n39845), .C2(n30489), .ZN(n7467) );
  OAI222_X1 U30753 ( .A1(n40934), .A2(n39855), .B1(n41318), .B2(n39848), .C1(
        n39845), .C2(n30488), .ZN(n7466) );
  OAI222_X1 U30754 ( .A1(n40940), .A2(n39855), .B1(n41324), .B2(n39848), .C1(
        n39845), .C2(n30487), .ZN(n7465) );
  OAI222_X1 U30755 ( .A1(n40946), .A2(n39855), .B1(n41330), .B2(n39848), .C1(
        n39845), .C2(n30486), .ZN(n7464) );
  OAI222_X1 U30756 ( .A1(n40958), .A2(n39855), .B1(n41342), .B2(n39848), .C1(
        n39845), .C2(n30484), .ZN(n7462) );
  AOI221_X1 U30757 ( .B1(n39102), .B2(n33031), .C1(n39096), .C2(n32983), .A(
        n37026), .ZN(n37021) );
  OAI222_X1 U30758 ( .A1(n30789), .A2(n39090), .B1(n30853), .B2(n39084), .C1(
        n30725), .C2(n39078), .ZN(n37026) );
  AOI221_X1 U30759 ( .B1(n39103), .B2(n33030), .C1(n39097), .C2(n32982), .A(
        n37007), .ZN(n37002) );
  OAI222_X1 U30760 ( .A1(n30788), .A2(n39091), .B1(n30852), .B2(n39085), .C1(
        n30724), .C2(n39079), .ZN(n37007) );
  AOI221_X1 U30761 ( .B1(n39103), .B2(n33029), .C1(n39097), .C2(n32981), .A(
        n36988), .ZN(n36983) );
  OAI222_X1 U30762 ( .A1(n30787), .A2(n39091), .B1(n30851), .B2(n39085), .C1(
        n30723), .C2(n39079), .ZN(n36988) );
  AOI221_X1 U30763 ( .B1(n39103), .B2(n33028), .C1(n39097), .C2(n32980), .A(
        n36969), .ZN(n36964) );
  OAI222_X1 U30764 ( .A1(n30786), .A2(n39091), .B1(n30850), .B2(n39085), .C1(
        n30722), .C2(n39079), .ZN(n36969) );
  AOI221_X1 U30765 ( .B1(n39103), .B2(n33027), .C1(n39097), .C2(n32979), .A(
        n36950), .ZN(n36945) );
  OAI222_X1 U30766 ( .A1(n30785), .A2(n39091), .B1(n30849), .B2(n39085), .C1(
        n30721), .C2(n39079), .ZN(n36950) );
  AOI221_X1 U30767 ( .B1(n39103), .B2(n33026), .C1(n39097), .C2(n32978), .A(
        n36931), .ZN(n36926) );
  OAI222_X1 U30768 ( .A1(n30784), .A2(n39091), .B1(n30848), .B2(n39085), .C1(
        n30720), .C2(n39079), .ZN(n36931) );
  AOI221_X1 U30769 ( .B1(n39103), .B2(n33025), .C1(n39097), .C2(n32977), .A(
        n36912), .ZN(n36907) );
  OAI222_X1 U30770 ( .A1(n30783), .A2(n39091), .B1(n30847), .B2(n39085), .C1(
        n30719), .C2(n39079), .ZN(n36912) );
  AOI221_X1 U30771 ( .B1(n39103), .B2(n33024), .C1(n39097), .C2(n32976), .A(
        n36893), .ZN(n36888) );
  OAI222_X1 U30772 ( .A1(n30782), .A2(n39091), .B1(n30846), .B2(n39085), .C1(
        n30718), .C2(n39079), .ZN(n36893) );
  AOI221_X1 U30773 ( .B1(n39103), .B2(n33023), .C1(n39097), .C2(n32975), .A(
        n36874), .ZN(n36869) );
  OAI222_X1 U30774 ( .A1(n30781), .A2(n39091), .B1(n30845), .B2(n39085), .C1(
        n30717), .C2(n39079), .ZN(n36874) );
  AOI221_X1 U30775 ( .B1(n39103), .B2(n33022), .C1(n39097), .C2(n32974), .A(
        n36855), .ZN(n36850) );
  OAI222_X1 U30776 ( .A1(n30780), .A2(n39091), .B1(n30844), .B2(n39085), .C1(
        n30716), .C2(n39079), .ZN(n36855) );
  AOI221_X1 U30777 ( .B1(n39103), .B2(n33021), .C1(n39097), .C2(n32973), .A(
        n36836), .ZN(n36831) );
  OAI222_X1 U30778 ( .A1(n30779), .A2(n39091), .B1(n30843), .B2(n39085), .C1(
        n30715), .C2(n39079), .ZN(n36836) );
  AOI221_X1 U30779 ( .B1(n39103), .B2(n33020), .C1(n39097), .C2(n32972), .A(
        n36817), .ZN(n36812) );
  OAI222_X1 U30780 ( .A1(n30778), .A2(n39091), .B1(n30842), .B2(n39085), .C1(
        n30714), .C2(n39079), .ZN(n36817) );
  AOI221_X1 U30781 ( .B1(n39103), .B2(n33019), .C1(n39097), .C2(n32971), .A(
        n36798), .ZN(n36793) );
  OAI222_X1 U30782 ( .A1(n30777), .A2(n39091), .B1(n30841), .B2(n39085), .C1(
        n30713), .C2(n39079), .ZN(n36798) );
  AOI221_X1 U30783 ( .B1(n39104), .B2(n33018), .C1(n39098), .C2(n32970), .A(
        n36779), .ZN(n36774) );
  OAI222_X1 U30784 ( .A1(n30776), .A2(n39092), .B1(n30840), .B2(n39086), .C1(
        n30712), .C2(n39080), .ZN(n36779) );
  AOI221_X1 U30785 ( .B1(n39104), .B2(n33017), .C1(n39098), .C2(n32969), .A(
        n36760), .ZN(n36755) );
  OAI222_X1 U30786 ( .A1(n30775), .A2(n39092), .B1(n30839), .B2(n39086), .C1(
        n30711), .C2(n39080), .ZN(n36760) );
  AOI221_X1 U30787 ( .B1(n39104), .B2(n33016), .C1(n39098), .C2(n32968), .A(
        n36741), .ZN(n36736) );
  OAI222_X1 U30788 ( .A1(n30774), .A2(n39092), .B1(n30838), .B2(n39086), .C1(
        n30710), .C2(n39080), .ZN(n36741) );
  AOI221_X1 U30789 ( .B1(n39104), .B2(n33015), .C1(n39098), .C2(n32967), .A(
        n36722), .ZN(n36717) );
  OAI222_X1 U30790 ( .A1(n30773), .A2(n39092), .B1(n30837), .B2(n39086), .C1(
        n30709), .C2(n39080), .ZN(n36722) );
  AOI221_X1 U30791 ( .B1(n39104), .B2(n33014), .C1(n39098), .C2(n32966), .A(
        n36703), .ZN(n36698) );
  OAI222_X1 U30792 ( .A1(n30772), .A2(n39092), .B1(n30836), .B2(n39086), .C1(
        n30708), .C2(n39080), .ZN(n36703) );
  AOI221_X1 U30793 ( .B1(n39104), .B2(n33013), .C1(n39098), .C2(n32965), .A(
        n36684), .ZN(n36679) );
  OAI222_X1 U30794 ( .A1(n30771), .A2(n39092), .B1(n30835), .B2(n39086), .C1(
        n30707), .C2(n39080), .ZN(n36684) );
  AOI221_X1 U30795 ( .B1(n39104), .B2(n33012), .C1(n39098), .C2(n32964), .A(
        n36665), .ZN(n36660) );
  OAI222_X1 U30796 ( .A1(n30770), .A2(n39092), .B1(n30834), .B2(n39086), .C1(
        n30706), .C2(n39080), .ZN(n36665) );
  AOI221_X1 U30797 ( .B1(n39104), .B2(n33011), .C1(n39098), .C2(n32963), .A(
        n36646), .ZN(n36641) );
  OAI222_X1 U30798 ( .A1(n30769), .A2(n39092), .B1(n30833), .B2(n39086), .C1(
        n30705), .C2(n39080), .ZN(n36646) );
  AOI221_X1 U30799 ( .B1(n39104), .B2(n33010), .C1(n39098), .C2(n32962), .A(
        n36627), .ZN(n36622) );
  OAI222_X1 U30800 ( .A1(n30768), .A2(n39092), .B1(n30832), .B2(n39086), .C1(
        n30704), .C2(n39080), .ZN(n36627) );
  AOI221_X1 U30801 ( .B1(n39104), .B2(n33009), .C1(n39098), .C2(n32961), .A(
        n36608), .ZN(n36603) );
  OAI222_X1 U30802 ( .A1(n30767), .A2(n39092), .B1(n30831), .B2(n39086), .C1(
        n30703), .C2(n39080), .ZN(n36608) );
  AOI221_X1 U30803 ( .B1(n39104), .B2(n33008), .C1(n39098), .C2(n32960), .A(
        n36589), .ZN(n36584) );
  OAI222_X1 U30804 ( .A1(n30766), .A2(n39092), .B1(n30830), .B2(n39086), .C1(
        n30702), .C2(n39080), .ZN(n36589) );
  AOI221_X1 U30805 ( .B1(n39104), .B2(n33007), .C1(n39098), .C2(n32959), .A(
        n36570), .ZN(n36565) );
  OAI222_X1 U30806 ( .A1(n30765), .A2(n39092), .B1(n30829), .B2(n39086), .C1(
        n30701), .C2(n39080), .ZN(n36570) );
  AOI221_X1 U30807 ( .B1(n39105), .B2(n33006), .C1(n39099), .C2(n32958), .A(
        n36551), .ZN(n36546) );
  OAI222_X1 U30808 ( .A1(n30764), .A2(n39093), .B1(n30828), .B2(n39087), .C1(
        n30700), .C2(n39081), .ZN(n36551) );
  AOI221_X1 U30809 ( .B1(n39105), .B2(n33005), .C1(n39099), .C2(n32957), .A(
        n36532), .ZN(n36527) );
  OAI222_X1 U30810 ( .A1(n30763), .A2(n39093), .B1(n30827), .B2(n39087), .C1(
        n30699), .C2(n39081), .ZN(n36532) );
  AOI221_X1 U30811 ( .B1(n39105), .B2(n33004), .C1(n39099), .C2(n32956), .A(
        n36513), .ZN(n36508) );
  OAI222_X1 U30812 ( .A1(n30762), .A2(n39093), .B1(n30826), .B2(n39087), .C1(
        n30698), .C2(n39081), .ZN(n36513) );
  AOI221_X1 U30813 ( .B1(n39105), .B2(n33003), .C1(n39099), .C2(n32955), .A(
        n36494), .ZN(n36489) );
  OAI222_X1 U30814 ( .A1(n30761), .A2(n39093), .B1(n30825), .B2(n39087), .C1(
        n30697), .C2(n39081), .ZN(n36494) );
  AOI221_X1 U30815 ( .B1(n39105), .B2(n33002), .C1(n39099), .C2(n32954), .A(
        n36475), .ZN(n36470) );
  OAI222_X1 U30816 ( .A1(n30760), .A2(n39093), .B1(n30824), .B2(n39087), .C1(
        n30696), .C2(n39081), .ZN(n36475) );
  AOI221_X1 U30817 ( .B1(n39105), .B2(n33001), .C1(n39099), .C2(n32953), .A(
        n36456), .ZN(n36451) );
  OAI222_X1 U30818 ( .A1(n30759), .A2(n39093), .B1(n30823), .B2(n39087), .C1(
        n30695), .C2(n39081), .ZN(n36456) );
  AOI221_X1 U30819 ( .B1(n39105), .B2(n33000), .C1(n39099), .C2(n32952), .A(
        n36437), .ZN(n36432) );
  OAI222_X1 U30820 ( .A1(n30758), .A2(n39093), .B1(n30822), .B2(n39087), .C1(
        n30694), .C2(n39081), .ZN(n36437) );
  AOI221_X1 U30821 ( .B1(n39105), .B2(n32999), .C1(n39099), .C2(n32951), .A(
        n36418), .ZN(n36413) );
  OAI222_X1 U30822 ( .A1(n30757), .A2(n39093), .B1(n30821), .B2(n39087), .C1(
        n30693), .C2(n39081), .ZN(n36418) );
  AOI221_X1 U30823 ( .B1(n39105), .B2(n32998), .C1(n39099), .C2(n32950), .A(
        n36399), .ZN(n36394) );
  OAI222_X1 U30824 ( .A1(n30756), .A2(n39093), .B1(n30820), .B2(n39087), .C1(
        n30692), .C2(n39081), .ZN(n36399) );
  AOI221_X1 U30825 ( .B1(n39105), .B2(n32997), .C1(n39099), .C2(n32949), .A(
        n36380), .ZN(n36375) );
  OAI222_X1 U30826 ( .A1(n30755), .A2(n39093), .B1(n30819), .B2(n39087), .C1(
        n30691), .C2(n39081), .ZN(n36380) );
  AOI221_X1 U30827 ( .B1(n39105), .B2(n32996), .C1(n39099), .C2(n32948), .A(
        n36361), .ZN(n36356) );
  OAI222_X1 U30828 ( .A1(n30754), .A2(n39093), .B1(n30818), .B2(n39087), .C1(
        n30690), .C2(n39081), .ZN(n36361) );
  AOI221_X1 U30829 ( .B1(n39105), .B2(n32995), .C1(n39099), .C2(n32947), .A(
        n36342), .ZN(n36337) );
  OAI222_X1 U30830 ( .A1(n30753), .A2(n39093), .B1(n30817), .B2(n39087), .C1(
        n30689), .C2(n39081), .ZN(n36342) );
  AOI221_X1 U30831 ( .B1(n39106), .B2(n32994), .C1(n39100), .C2(n32946), .A(
        n36323), .ZN(n36318) );
  OAI222_X1 U30832 ( .A1(n30752), .A2(n39094), .B1(n30816), .B2(n39088), .C1(
        n30688), .C2(n39082), .ZN(n36323) );
  AOI221_X1 U30833 ( .B1(n39106), .B2(n32993), .C1(n39100), .C2(n32945), .A(
        n36304), .ZN(n36299) );
  OAI222_X1 U30834 ( .A1(n30751), .A2(n39094), .B1(n30815), .B2(n39088), .C1(
        n30687), .C2(n39082), .ZN(n36304) );
  AOI221_X1 U30835 ( .B1(n39106), .B2(n32992), .C1(n39100), .C2(n32944), .A(
        n36285), .ZN(n36280) );
  OAI222_X1 U30836 ( .A1(n30750), .A2(n39094), .B1(n30814), .B2(n39088), .C1(
        n30686), .C2(n39082), .ZN(n36285) );
  AOI221_X1 U30837 ( .B1(n39106), .B2(n32991), .C1(n39100), .C2(n32943), .A(
        n36266), .ZN(n36261) );
  OAI222_X1 U30838 ( .A1(n30749), .A2(n39094), .B1(n30813), .B2(n39088), .C1(
        n30685), .C2(n39082), .ZN(n36266) );
  AOI221_X1 U30839 ( .B1(n39106), .B2(n33134), .C1(n39100), .C2(n33122), .A(
        n36247), .ZN(n36242) );
  OAI222_X1 U30840 ( .A1(n30748), .A2(n39094), .B1(n30812), .B2(n39088), .C1(
        n30684), .C2(n39082), .ZN(n36247) );
  AOI221_X1 U30841 ( .B1(n39106), .B2(n33133), .C1(n39100), .C2(n33121), .A(
        n36228), .ZN(n36223) );
  OAI222_X1 U30842 ( .A1(n30747), .A2(n39094), .B1(n30811), .B2(n39088), .C1(
        n30683), .C2(n39082), .ZN(n36228) );
  AOI221_X1 U30843 ( .B1(n39102), .B2(n32490), .C1(n39096), .C2(n32486), .A(
        n37216), .ZN(n37211) );
  OAI222_X1 U30844 ( .A1(n30799), .A2(n39090), .B1(n30863), .B2(n39084), .C1(
        n30735), .C2(n39078), .ZN(n37216) );
  AOI221_X1 U30845 ( .B1(n39102), .B2(n32489), .C1(n39096), .C2(n32485), .A(
        n37197), .ZN(n37192) );
  OAI222_X1 U30846 ( .A1(n30798), .A2(n39090), .B1(n30862), .B2(n39084), .C1(
        n30734), .C2(n39078), .ZN(n37197) );
  AOI221_X1 U30847 ( .B1(n39102), .B2(n32488), .C1(n39096), .C2(n32484), .A(
        n37178), .ZN(n37173) );
  OAI222_X1 U30848 ( .A1(n30797), .A2(n39090), .B1(n30861), .B2(n39084), .C1(
        n30733), .C2(n39078), .ZN(n37178) );
  AOI221_X1 U30849 ( .B1(n39102), .B2(n33038), .C1(n39096), .C2(n32990), .A(
        n37159), .ZN(n37154) );
  OAI222_X1 U30850 ( .A1(n30796), .A2(n39090), .B1(n30860), .B2(n39084), .C1(
        n30732), .C2(n39078), .ZN(n37159) );
  AOI221_X1 U30851 ( .B1(n39102), .B2(n33037), .C1(n39096), .C2(n32989), .A(
        n37140), .ZN(n37135) );
  OAI222_X1 U30852 ( .A1(n30795), .A2(n39090), .B1(n30859), .B2(n39084), .C1(
        n30731), .C2(n39078), .ZN(n37140) );
  AOI221_X1 U30853 ( .B1(n39107), .B2(n33126), .C1(n39101), .C2(n33114), .A(
        n36095), .ZN(n36090) );
  OAI222_X1 U30854 ( .A1(n30740), .A2(n39095), .B1(n30804), .B2(n39089), .C1(
        n30676), .C2(n39083), .ZN(n36095) );
  AOI221_X1 U30855 ( .B1(n39107), .B2(n33125), .C1(n39101), .C2(n33113), .A(
        n36076), .ZN(n36071) );
  OAI222_X1 U30856 ( .A1(n30739), .A2(n39095), .B1(n30803), .B2(n39089), .C1(
        n30675), .C2(n39083), .ZN(n36076) );
  AOI221_X1 U30857 ( .B1(n39107), .B2(n33124), .C1(n39101), .C2(n33112), .A(
        n36057), .ZN(n36052) );
  OAI222_X1 U30858 ( .A1(n30738), .A2(n39095), .B1(n30802), .B2(n39089), .C1(
        n30674), .C2(n39083), .ZN(n36057) );
  AOI221_X1 U30859 ( .B1(n39107), .B2(n33123), .C1(n39101), .C2(n33111), .A(
        n36030), .ZN(n36013) );
  OAI222_X1 U30860 ( .A1(n30737), .A2(n39095), .B1(n30801), .B2(n39089), .C1(
        n30673), .C2(n39083), .ZN(n36030) );
  AOI221_X1 U30861 ( .B1(n39102), .B2(n32491), .C1(n39096), .C2(n32487), .A(
        n37248), .ZN(n37242) );
  OAI222_X1 U30862 ( .A1(n30800), .A2(n39090), .B1(n30864), .B2(n39084), .C1(
        n30736), .C2(n39078), .ZN(n37248) );
  AOI221_X1 U30863 ( .B1(n39102), .B2(n33036), .C1(n39096), .C2(n32988), .A(
        n37121), .ZN(n37116) );
  OAI222_X1 U30864 ( .A1(n30794), .A2(n39090), .B1(n30858), .B2(n39084), .C1(
        n30730), .C2(n39078), .ZN(n37121) );
  AOI221_X1 U30865 ( .B1(n39102), .B2(n33035), .C1(n39096), .C2(n32987), .A(
        n37102), .ZN(n37097) );
  OAI222_X1 U30866 ( .A1(n30793), .A2(n39090), .B1(n30857), .B2(n39084), .C1(
        n30729), .C2(n39078), .ZN(n37102) );
  AOI221_X1 U30867 ( .B1(n39102), .B2(n33034), .C1(n39096), .C2(n32986), .A(
        n37083), .ZN(n37078) );
  OAI222_X1 U30868 ( .A1(n30792), .A2(n39090), .B1(n30856), .B2(n39084), .C1(
        n30728), .C2(n39078), .ZN(n37083) );
  AOI221_X1 U30869 ( .B1(n39102), .B2(n33033), .C1(n39096), .C2(n32985), .A(
        n37064), .ZN(n37059) );
  OAI222_X1 U30870 ( .A1(n30791), .A2(n39090), .B1(n30855), .B2(n39084), .C1(
        n30727), .C2(n39078), .ZN(n37064) );
  AOI221_X1 U30871 ( .B1(n39102), .B2(n33032), .C1(n39096), .C2(n32984), .A(
        n37045), .ZN(n37040) );
  OAI222_X1 U30872 ( .A1(n30790), .A2(n39090), .B1(n30854), .B2(n39084), .C1(
        n30726), .C2(n39078), .ZN(n37045) );
  AOI221_X1 U30873 ( .B1(n39106), .B2(n33132), .C1(n39100), .C2(n33120), .A(
        n36209), .ZN(n36204) );
  OAI222_X1 U30874 ( .A1(n30746), .A2(n39094), .B1(n30810), .B2(n39088), .C1(
        n30682), .C2(n39082), .ZN(n36209) );
  AOI221_X1 U30875 ( .B1(n39106), .B2(n33131), .C1(n39100), .C2(n33119), .A(
        n36190), .ZN(n36185) );
  OAI222_X1 U30876 ( .A1(n30745), .A2(n39094), .B1(n30809), .B2(n39088), .C1(
        n30681), .C2(n39082), .ZN(n36190) );
  AOI221_X1 U30877 ( .B1(n39106), .B2(n33130), .C1(n39100), .C2(n33118), .A(
        n36171), .ZN(n36166) );
  OAI222_X1 U30878 ( .A1(n30744), .A2(n39094), .B1(n30808), .B2(n39088), .C1(
        n30680), .C2(n39082), .ZN(n36171) );
  AOI221_X1 U30879 ( .B1(n39106), .B2(n33129), .C1(n39100), .C2(n33117), .A(
        n36152), .ZN(n36147) );
  OAI222_X1 U30880 ( .A1(n30743), .A2(n39094), .B1(n30807), .B2(n39088), .C1(
        n30679), .C2(n39082), .ZN(n36152) );
  AOI221_X1 U30881 ( .B1(n39106), .B2(n33128), .C1(n39100), .C2(n33116), .A(
        n36133), .ZN(n36128) );
  OAI222_X1 U30882 ( .A1(n30742), .A2(n39094), .B1(n30806), .B2(n39088), .C1(
        n30678), .C2(n39082), .ZN(n36133) );
  AOI221_X1 U30883 ( .B1(n39106), .B2(n33127), .C1(n39100), .C2(n33115), .A(
        n36114), .ZN(n36109) );
  OAI222_X1 U30884 ( .A1(n30741), .A2(n39094), .B1(n30805), .B2(n39088), .C1(
        n30677), .C2(n39082), .ZN(n36114) );
  AOI221_X1 U30885 ( .B1(n39609), .B2(n32491), .C1(n39603), .C2(n32487), .A(
        n33475), .ZN(n33458) );
  OAI222_X1 U30886 ( .A1(n30800), .A2(n39597), .B1(n30864), .B2(n39591), .C1(
        n30736), .C2(n39585), .ZN(n33475) );
  AOI221_X1 U30887 ( .B1(n39357), .B2(n32491), .C1(n39351), .C2(n32487), .A(
        n34749), .ZN(n34732) );
  OAI222_X1 U30888 ( .A1(n30800), .A2(n39345), .B1(n30864), .B2(n39339), .C1(
        n30736), .C2(n39333), .ZN(n34749) );
  AOI221_X1 U30889 ( .B1(n39609), .B2(n32490), .C1(n39603), .C2(n32486), .A(
        n33502), .ZN(n33497) );
  OAI222_X1 U30890 ( .A1(n30799), .A2(n39597), .B1(n30863), .B2(n39591), .C1(
        n30735), .C2(n39585), .ZN(n33502) );
  AOI221_X1 U30891 ( .B1(n39357), .B2(n32490), .C1(n39351), .C2(n32486), .A(
        n34776), .ZN(n34771) );
  OAI222_X1 U30892 ( .A1(n30799), .A2(n39345), .B1(n30863), .B2(n39339), .C1(
        n30735), .C2(n39333), .ZN(n34776) );
  AOI221_X1 U30893 ( .B1(n39609), .B2(n32489), .C1(n39603), .C2(n32485), .A(
        n33521), .ZN(n33516) );
  OAI222_X1 U30894 ( .A1(n30798), .A2(n39597), .B1(n30862), .B2(n39591), .C1(
        n30734), .C2(n39585), .ZN(n33521) );
  AOI221_X1 U30895 ( .B1(n39357), .B2(n32489), .C1(n39351), .C2(n32485), .A(
        n34795), .ZN(n34790) );
  OAI222_X1 U30896 ( .A1(n30798), .A2(n39345), .B1(n30862), .B2(n39339), .C1(
        n30734), .C2(n39333), .ZN(n34795) );
  AOI221_X1 U30897 ( .B1(n39609), .B2(n32488), .C1(n39603), .C2(n32484), .A(
        n33540), .ZN(n33535) );
  OAI222_X1 U30898 ( .A1(n30797), .A2(n39597), .B1(n30861), .B2(n39591), .C1(
        n30733), .C2(n39585), .ZN(n33540) );
  AOI221_X1 U30899 ( .B1(n39357), .B2(n32488), .C1(n39351), .C2(n32484), .A(
        n34814), .ZN(n34809) );
  OAI222_X1 U30900 ( .A1(n30797), .A2(n39345), .B1(n30861), .B2(n39339), .C1(
        n30733), .C2(n39333), .ZN(n34814) );
  AOI221_X1 U30901 ( .B1(n39608), .B2(n33038), .C1(n39602), .C2(n32990), .A(
        n33559), .ZN(n33554) );
  OAI222_X1 U30902 ( .A1(n30796), .A2(n39596), .B1(n30860), .B2(n39590), .C1(
        n30732), .C2(n39584), .ZN(n33559) );
  AOI221_X1 U30903 ( .B1(n39356), .B2(n33038), .C1(n39350), .C2(n32990), .A(
        n34833), .ZN(n34828) );
  OAI222_X1 U30904 ( .A1(n30796), .A2(n39344), .B1(n30860), .B2(n39338), .C1(
        n30732), .C2(n39332), .ZN(n34833) );
  AOI221_X1 U30905 ( .B1(n39608), .B2(n33037), .C1(n39602), .C2(n32989), .A(
        n33578), .ZN(n33573) );
  OAI222_X1 U30906 ( .A1(n30795), .A2(n39596), .B1(n30859), .B2(n39590), .C1(
        n30731), .C2(n39584), .ZN(n33578) );
  AOI221_X1 U30907 ( .B1(n39356), .B2(n33037), .C1(n39350), .C2(n32989), .A(
        n34852), .ZN(n34847) );
  OAI222_X1 U30908 ( .A1(n30795), .A2(n39344), .B1(n30859), .B2(n39338), .C1(
        n30731), .C2(n39332), .ZN(n34852) );
  AOI221_X1 U30909 ( .B1(n39608), .B2(n33036), .C1(n39602), .C2(n32988), .A(
        n33597), .ZN(n33592) );
  OAI222_X1 U30910 ( .A1(n30794), .A2(n39596), .B1(n30858), .B2(n39590), .C1(
        n30730), .C2(n39584), .ZN(n33597) );
  AOI221_X1 U30911 ( .B1(n39356), .B2(n33036), .C1(n39350), .C2(n32988), .A(
        n34871), .ZN(n34866) );
  OAI222_X1 U30912 ( .A1(n30794), .A2(n39344), .B1(n30858), .B2(n39338), .C1(
        n30730), .C2(n39332), .ZN(n34871) );
  AOI221_X1 U30913 ( .B1(n39608), .B2(n33035), .C1(n39602), .C2(n32987), .A(
        n33616), .ZN(n33611) );
  OAI222_X1 U30914 ( .A1(n30793), .A2(n39596), .B1(n30857), .B2(n39590), .C1(
        n30729), .C2(n39584), .ZN(n33616) );
  AOI221_X1 U30915 ( .B1(n39356), .B2(n33035), .C1(n39350), .C2(n32987), .A(
        n34890), .ZN(n34885) );
  OAI222_X1 U30916 ( .A1(n30793), .A2(n39344), .B1(n30857), .B2(n39338), .C1(
        n30729), .C2(n39332), .ZN(n34890) );
  AOI221_X1 U30917 ( .B1(n39608), .B2(n33034), .C1(n39602), .C2(n32986), .A(
        n33635), .ZN(n33630) );
  OAI222_X1 U30918 ( .A1(n30792), .A2(n39596), .B1(n30856), .B2(n39590), .C1(
        n30728), .C2(n39584), .ZN(n33635) );
  AOI221_X1 U30919 ( .B1(n39356), .B2(n33034), .C1(n39350), .C2(n32986), .A(
        n34909), .ZN(n34904) );
  OAI222_X1 U30920 ( .A1(n30792), .A2(n39344), .B1(n30856), .B2(n39338), .C1(
        n30728), .C2(n39332), .ZN(n34909) );
  AOI221_X1 U30921 ( .B1(n39608), .B2(n33033), .C1(n39602), .C2(n32985), .A(
        n33654), .ZN(n33649) );
  OAI222_X1 U30922 ( .A1(n30791), .A2(n39596), .B1(n30855), .B2(n39590), .C1(
        n30727), .C2(n39584), .ZN(n33654) );
  AOI221_X1 U30923 ( .B1(n39356), .B2(n33033), .C1(n39350), .C2(n32985), .A(
        n34928), .ZN(n34923) );
  OAI222_X1 U30924 ( .A1(n30791), .A2(n39344), .B1(n30855), .B2(n39338), .C1(
        n30727), .C2(n39332), .ZN(n34928) );
  AOI221_X1 U30925 ( .B1(n39608), .B2(n33032), .C1(n39602), .C2(n32984), .A(
        n33673), .ZN(n33668) );
  OAI222_X1 U30926 ( .A1(n30790), .A2(n39596), .B1(n30854), .B2(n39590), .C1(
        n30726), .C2(n39584), .ZN(n33673) );
  AOI221_X1 U30927 ( .B1(n39356), .B2(n33032), .C1(n39350), .C2(n32984), .A(
        n34947), .ZN(n34942) );
  OAI222_X1 U30928 ( .A1(n30790), .A2(n39344), .B1(n30854), .B2(n39338), .C1(
        n30726), .C2(n39332), .ZN(n34947) );
  AOI221_X1 U30929 ( .B1(n39608), .B2(n33031), .C1(n39602), .C2(n32983), .A(
        n33692), .ZN(n33687) );
  OAI222_X1 U30930 ( .A1(n30789), .A2(n39596), .B1(n30853), .B2(n39590), .C1(
        n30725), .C2(n39584), .ZN(n33692) );
  AOI221_X1 U30931 ( .B1(n39356), .B2(n33031), .C1(n39350), .C2(n32983), .A(
        n34966), .ZN(n34961) );
  OAI222_X1 U30932 ( .A1(n30789), .A2(n39344), .B1(n30853), .B2(n39338), .C1(
        n30725), .C2(n39332), .ZN(n34966) );
  AOI221_X1 U30933 ( .B1(n39608), .B2(n33030), .C1(n39602), .C2(n32982), .A(
        n33711), .ZN(n33706) );
  OAI222_X1 U30934 ( .A1(n30788), .A2(n39596), .B1(n30852), .B2(n39590), .C1(
        n30724), .C2(n39584), .ZN(n33711) );
  AOI221_X1 U30935 ( .B1(n39356), .B2(n33030), .C1(n39350), .C2(n32982), .A(
        n34985), .ZN(n34980) );
  OAI222_X1 U30936 ( .A1(n30788), .A2(n39344), .B1(n30852), .B2(n39338), .C1(
        n30724), .C2(n39332), .ZN(n34985) );
  AOI221_X1 U30937 ( .B1(n39608), .B2(n33029), .C1(n39602), .C2(n32981), .A(
        n33730), .ZN(n33725) );
  OAI222_X1 U30938 ( .A1(n30787), .A2(n39596), .B1(n30851), .B2(n39590), .C1(
        n30723), .C2(n39584), .ZN(n33730) );
  AOI221_X1 U30939 ( .B1(n39356), .B2(n33029), .C1(n39350), .C2(n32981), .A(
        n35004), .ZN(n34999) );
  OAI222_X1 U30940 ( .A1(n30787), .A2(n39344), .B1(n30851), .B2(n39338), .C1(
        n30723), .C2(n39332), .ZN(n35004) );
  AOI221_X1 U30941 ( .B1(n39608), .B2(n33028), .C1(n39602), .C2(n32980), .A(
        n33749), .ZN(n33744) );
  OAI222_X1 U30942 ( .A1(n30786), .A2(n39596), .B1(n30850), .B2(n39590), .C1(
        n30722), .C2(n39584), .ZN(n33749) );
  AOI221_X1 U30943 ( .B1(n39356), .B2(n33028), .C1(n39350), .C2(n32980), .A(
        n35023), .ZN(n35018) );
  OAI222_X1 U30944 ( .A1(n30786), .A2(n39344), .B1(n30850), .B2(n39338), .C1(
        n30722), .C2(n39332), .ZN(n35023) );
  AOI221_X1 U30945 ( .B1(n39608), .B2(n33027), .C1(n39602), .C2(n32979), .A(
        n33768), .ZN(n33763) );
  OAI222_X1 U30946 ( .A1(n30785), .A2(n39596), .B1(n30849), .B2(n39590), .C1(
        n30721), .C2(n39584), .ZN(n33768) );
  AOI221_X1 U30947 ( .B1(n39356), .B2(n33027), .C1(n39350), .C2(n32979), .A(
        n35042), .ZN(n35037) );
  OAI222_X1 U30948 ( .A1(n30785), .A2(n39344), .B1(n30849), .B2(n39338), .C1(
        n30721), .C2(n39332), .ZN(n35042) );
  AOI221_X1 U30949 ( .B1(n39607), .B2(n33026), .C1(n39601), .C2(n32978), .A(
        n33787), .ZN(n33782) );
  OAI222_X1 U30950 ( .A1(n30784), .A2(n39595), .B1(n30848), .B2(n39589), .C1(
        n30720), .C2(n39583), .ZN(n33787) );
  AOI221_X1 U30951 ( .B1(n39355), .B2(n33026), .C1(n39349), .C2(n32978), .A(
        n35061), .ZN(n35056) );
  OAI222_X1 U30952 ( .A1(n30784), .A2(n39343), .B1(n30848), .B2(n39337), .C1(
        n30720), .C2(n39331), .ZN(n35061) );
  AOI221_X1 U30953 ( .B1(n39607), .B2(n33025), .C1(n39601), .C2(n32977), .A(
        n33806), .ZN(n33801) );
  OAI222_X1 U30954 ( .A1(n30783), .A2(n39595), .B1(n30847), .B2(n39589), .C1(
        n30719), .C2(n39583), .ZN(n33806) );
  AOI221_X1 U30955 ( .B1(n39355), .B2(n33025), .C1(n39349), .C2(n32977), .A(
        n35080), .ZN(n35075) );
  OAI222_X1 U30956 ( .A1(n30783), .A2(n39343), .B1(n30847), .B2(n39337), .C1(
        n30719), .C2(n39331), .ZN(n35080) );
  AOI221_X1 U30957 ( .B1(n39607), .B2(n33024), .C1(n39601), .C2(n32976), .A(
        n33825), .ZN(n33820) );
  OAI222_X1 U30958 ( .A1(n30782), .A2(n39595), .B1(n30846), .B2(n39589), .C1(
        n30718), .C2(n39583), .ZN(n33825) );
  AOI221_X1 U30959 ( .B1(n39355), .B2(n33024), .C1(n39349), .C2(n32976), .A(
        n35099), .ZN(n35094) );
  OAI222_X1 U30960 ( .A1(n30782), .A2(n39343), .B1(n30846), .B2(n39337), .C1(
        n30718), .C2(n39331), .ZN(n35099) );
  AOI221_X1 U30961 ( .B1(n39607), .B2(n33023), .C1(n39601), .C2(n32975), .A(
        n33844), .ZN(n33839) );
  OAI222_X1 U30962 ( .A1(n30781), .A2(n39595), .B1(n30845), .B2(n39589), .C1(
        n30717), .C2(n39583), .ZN(n33844) );
  AOI221_X1 U30963 ( .B1(n39355), .B2(n33023), .C1(n39349), .C2(n32975), .A(
        n35118), .ZN(n35113) );
  OAI222_X1 U30964 ( .A1(n30781), .A2(n39343), .B1(n30845), .B2(n39337), .C1(
        n30717), .C2(n39331), .ZN(n35118) );
  AOI221_X1 U30965 ( .B1(n39607), .B2(n33022), .C1(n39601), .C2(n32974), .A(
        n33863), .ZN(n33858) );
  OAI222_X1 U30966 ( .A1(n30780), .A2(n39595), .B1(n30844), .B2(n39589), .C1(
        n30716), .C2(n39583), .ZN(n33863) );
  AOI221_X1 U30967 ( .B1(n39355), .B2(n33022), .C1(n39349), .C2(n32974), .A(
        n35137), .ZN(n35132) );
  OAI222_X1 U30968 ( .A1(n30780), .A2(n39343), .B1(n30844), .B2(n39337), .C1(
        n30716), .C2(n39331), .ZN(n35137) );
  AOI221_X1 U30969 ( .B1(n39607), .B2(n33021), .C1(n39601), .C2(n32973), .A(
        n33882), .ZN(n33877) );
  OAI222_X1 U30970 ( .A1(n30779), .A2(n39595), .B1(n30843), .B2(n39589), .C1(
        n30715), .C2(n39583), .ZN(n33882) );
  AOI221_X1 U30971 ( .B1(n39355), .B2(n33021), .C1(n39349), .C2(n32973), .A(
        n35156), .ZN(n35151) );
  OAI222_X1 U30972 ( .A1(n30779), .A2(n39343), .B1(n30843), .B2(n39337), .C1(
        n30715), .C2(n39331), .ZN(n35156) );
  AOI221_X1 U30973 ( .B1(n39607), .B2(n33020), .C1(n39601), .C2(n32972), .A(
        n33901), .ZN(n33896) );
  OAI222_X1 U30974 ( .A1(n30778), .A2(n39595), .B1(n30842), .B2(n39589), .C1(
        n30714), .C2(n39583), .ZN(n33901) );
  AOI221_X1 U30975 ( .B1(n39355), .B2(n33020), .C1(n39349), .C2(n32972), .A(
        n35175), .ZN(n35170) );
  OAI222_X1 U30976 ( .A1(n30778), .A2(n39343), .B1(n30842), .B2(n39337), .C1(
        n30714), .C2(n39331), .ZN(n35175) );
  AOI221_X1 U30977 ( .B1(n39607), .B2(n33019), .C1(n39601), .C2(n32971), .A(
        n33920), .ZN(n33915) );
  OAI222_X1 U30978 ( .A1(n30777), .A2(n39595), .B1(n30841), .B2(n39589), .C1(
        n30713), .C2(n39583), .ZN(n33920) );
  AOI221_X1 U30979 ( .B1(n39355), .B2(n33019), .C1(n39349), .C2(n32971), .A(
        n35194), .ZN(n35189) );
  OAI222_X1 U30980 ( .A1(n30777), .A2(n39343), .B1(n30841), .B2(n39337), .C1(
        n30713), .C2(n39331), .ZN(n35194) );
  AOI221_X1 U30981 ( .B1(n39607), .B2(n33018), .C1(n39601), .C2(n32970), .A(
        n33939), .ZN(n33934) );
  OAI222_X1 U30982 ( .A1(n30776), .A2(n39595), .B1(n30840), .B2(n39589), .C1(
        n30712), .C2(n39583), .ZN(n33939) );
  AOI221_X1 U30983 ( .B1(n39355), .B2(n33018), .C1(n39349), .C2(n32970), .A(
        n35213), .ZN(n35208) );
  OAI222_X1 U30984 ( .A1(n30776), .A2(n39343), .B1(n30840), .B2(n39337), .C1(
        n30712), .C2(n39331), .ZN(n35213) );
  AOI221_X1 U30985 ( .B1(n39607), .B2(n33017), .C1(n39601), .C2(n32969), .A(
        n33958), .ZN(n33953) );
  OAI222_X1 U30986 ( .A1(n30775), .A2(n39595), .B1(n30839), .B2(n39589), .C1(
        n30711), .C2(n39583), .ZN(n33958) );
  AOI221_X1 U30987 ( .B1(n39355), .B2(n33017), .C1(n39349), .C2(n32969), .A(
        n35232), .ZN(n35227) );
  OAI222_X1 U30988 ( .A1(n30775), .A2(n39343), .B1(n30839), .B2(n39337), .C1(
        n30711), .C2(n39331), .ZN(n35232) );
  AOI221_X1 U30989 ( .B1(n39607), .B2(n33016), .C1(n39601), .C2(n32968), .A(
        n33977), .ZN(n33972) );
  OAI222_X1 U30990 ( .A1(n30774), .A2(n39595), .B1(n30838), .B2(n39589), .C1(
        n30710), .C2(n39583), .ZN(n33977) );
  AOI221_X1 U30991 ( .B1(n39355), .B2(n33016), .C1(n39349), .C2(n32968), .A(
        n35251), .ZN(n35246) );
  OAI222_X1 U30992 ( .A1(n30774), .A2(n39343), .B1(n30838), .B2(n39337), .C1(
        n30710), .C2(n39331), .ZN(n35251) );
  AOI221_X1 U30993 ( .B1(n39607), .B2(n33015), .C1(n39601), .C2(n32967), .A(
        n33996), .ZN(n33991) );
  OAI222_X1 U30994 ( .A1(n30773), .A2(n39595), .B1(n30837), .B2(n39589), .C1(
        n30709), .C2(n39583), .ZN(n33996) );
  AOI221_X1 U30995 ( .B1(n39355), .B2(n33015), .C1(n39349), .C2(n32967), .A(
        n35270), .ZN(n35265) );
  OAI222_X1 U30996 ( .A1(n30773), .A2(n39343), .B1(n30837), .B2(n39337), .C1(
        n30709), .C2(n39331), .ZN(n35270) );
  AOI221_X1 U30997 ( .B1(n39606), .B2(n33014), .C1(n39600), .C2(n32966), .A(
        n34015), .ZN(n34010) );
  OAI222_X1 U30998 ( .A1(n30772), .A2(n39594), .B1(n30836), .B2(n39588), .C1(
        n30708), .C2(n39582), .ZN(n34015) );
  AOI221_X1 U30999 ( .B1(n39354), .B2(n33014), .C1(n39348), .C2(n32966), .A(
        n35289), .ZN(n35284) );
  OAI222_X1 U31000 ( .A1(n30772), .A2(n39342), .B1(n30836), .B2(n39336), .C1(
        n30708), .C2(n39330), .ZN(n35289) );
  AOI221_X1 U31001 ( .B1(n39606), .B2(n33013), .C1(n39600), .C2(n32965), .A(
        n34034), .ZN(n34029) );
  OAI222_X1 U31002 ( .A1(n30771), .A2(n39594), .B1(n30835), .B2(n39588), .C1(
        n30707), .C2(n39582), .ZN(n34034) );
  AOI221_X1 U31003 ( .B1(n39354), .B2(n33013), .C1(n39348), .C2(n32965), .A(
        n35308), .ZN(n35303) );
  OAI222_X1 U31004 ( .A1(n30771), .A2(n39342), .B1(n30835), .B2(n39336), .C1(
        n30707), .C2(n39330), .ZN(n35308) );
  AOI221_X1 U31005 ( .B1(n39606), .B2(n33012), .C1(n39600), .C2(n32964), .A(
        n34053), .ZN(n34048) );
  OAI222_X1 U31006 ( .A1(n30770), .A2(n39594), .B1(n30834), .B2(n39588), .C1(
        n30706), .C2(n39582), .ZN(n34053) );
  AOI221_X1 U31007 ( .B1(n39354), .B2(n33012), .C1(n39348), .C2(n32964), .A(
        n35327), .ZN(n35322) );
  OAI222_X1 U31008 ( .A1(n30770), .A2(n39342), .B1(n30834), .B2(n39336), .C1(
        n30706), .C2(n39330), .ZN(n35327) );
  AOI221_X1 U31009 ( .B1(n39606), .B2(n33011), .C1(n39600), .C2(n32963), .A(
        n34072), .ZN(n34067) );
  OAI222_X1 U31010 ( .A1(n30769), .A2(n39594), .B1(n30833), .B2(n39588), .C1(
        n30705), .C2(n39582), .ZN(n34072) );
  AOI221_X1 U31011 ( .B1(n39354), .B2(n33011), .C1(n39348), .C2(n32963), .A(
        n35346), .ZN(n35341) );
  OAI222_X1 U31012 ( .A1(n30769), .A2(n39342), .B1(n30833), .B2(n39336), .C1(
        n30705), .C2(n39330), .ZN(n35346) );
  AOI221_X1 U31013 ( .B1(n39606), .B2(n33010), .C1(n39600), .C2(n32962), .A(
        n34091), .ZN(n34086) );
  OAI222_X1 U31014 ( .A1(n30768), .A2(n39594), .B1(n30832), .B2(n39588), .C1(
        n30704), .C2(n39582), .ZN(n34091) );
  AOI221_X1 U31015 ( .B1(n39354), .B2(n33010), .C1(n39348), .C2(n32962), .A(
        n35365), .ZN(n35360) );
  OAI222_X1 U31016 ( .A1(n30768), .A2(n39342), .B1(n30832), .B2(n39336), .C1(
        n30704), .C2(n39330), .ZN(n35365) );
  AOI221_X1 U31017 ( .B1(n39606), .B2(n33009), .C1(n39600), .C2(n32961), .A(
        n34110), .ZN(n34105) );
  OAI222_X1 U31018 ( .A1(n30767), .A2(n39594), .B1(n30831), .B2(n39588), .C1(
        n30703), .C2(n39582), .ZN(n34110) );
  AOI221_X1 U31019 ( .B1(n39354), .B2(n33009), .C1(n39348), .C2(n32961), .A(
        n35384), .ZN(n35379) );
  OAI222_X1 U31020 ( .A1(n30767), .A2(n39342), .B1(n30831), .B2(n39336), .C1(
        n30703), .C2(n39330), .ZN(n35384) );
  AOI221_X1 U31021 ( .B1(n39606), .B2(n33008), .C1(n39600), .C2(n32960), .A(
        n34129), .ZN(n34124) );
  OAI222_X1 U31022 ( .A1(n30766), .A2(n39594), .B1(n30830), .B2(n39588), .C1(
        n30702), .C2(n39582), .ZN(n34129) );
  AOI221_X1 U31023 ( .B1(n39354), .B2(n33008), .C1(n39348), .C2(n32960), .A(
        n35403), .ZN(n35398) );
  OAI222_X1 U31024 ( .A1(n30766), .A2(n39342), .B1(n30830), .B2(n39336), .C1(
        n30702), .C2(n39330), .ZN(n35403) );
  AOI221_X1 U31025 ( .B1(n39606), .B2(n33007), .C1(n39600), .C2(n32959), .A(
        n34148), .ZN(n34143) );
  OAI222_X1 U31026 ( .A1(n30765), .A2(n39594), .B1(n30829), .B2(n39588), .C1(
        n30701), .C2(n39582), .ZN(n34148) );
  AOI221_X1 U31027 ( .B1(n39354), .B2(n33007), .C1(n39348), .C2(n32959), .A(
        n35422), .ZN(n35417) );
  OAI222_X1 U31028 ( .A1(n30765), .A2(n39342), .B1(n30829), .B2(n39336), .C1(
        n30701), .C2(n39330), .ZN(n35422) );
  AOI221_X1 U31029 ( .B1(n39606), .B2(n33006), .C1(n39600), .C2(n32958), .A(
        n34167), .ZN(n34162) );
  OAI222_X1 U31030 ( .A1(n30764), .A2(n39594), .B1(n30828), .B2(n39588), .C1(
        n30700), .C2(n39582), .ZN(n34167) );
  AOI221_X1 U31031 ( .B1(n39354), .B2(n33006), .C1(n39348), .C2(n32958), .A(
        n35441), .ZN(n35436) );
  OAI222_X1 U31032 ( .A1(n30764), .A2(n39342), .B1(n30828), .B2(n39336), .C1(
        n30700), .C2(n39330), .ZN(n35441) );
  AOI221_X1 U31033 ( .B1(n39606), .B2(n33005), .C1(n39600), .C2(n32957), .A(
        n34186), .ZN(n34181) );
  OAI222_X1 U31034 ( .A1(n30763), .A2(n39594), .B1(n30827), .B2(n39588), .C1(
        n30699), .C2(n39582), .ZN(n34186) );
  AOI221_X1 U31035 ( .B1(n39354), .B2(n33005), .C1(n39348), .C2(n32957), .A(
        n35460), .ZN(n35455) );
  OAI222_X1 U31036 ( .A1(n30763), .A2(n39342), .B1(n30827), .B2(n39336), .C1(
        n30699), .C2(n39330), .ZN(n35460) );
  AOI221_X1 U31037 ( .B1(n39606), .B2(n33004), .C1(n39600), .C2(n32956), .A(
        n34205), .ZN(n34200) );
  OAI222_X1 U31038 ( .A1(n30762), .A2(n39594), .B1(n30826), .B2(n39588), .C1(
        n30698), .C2(n39582), .ZN(n34205) );
  AOI221_X1 U31039 ( .B1(n39354), .B2(n33004), .C1(n39348), .C2(n32956), .A(
        n35479), .ZN(n35474) );
  OAI222_X1 U31040 ( .A1(n30762), .A2(n39342), .B1(n30826), .B2(n39336), .C1(
        n30698), .C2(n39330), .ZN(n35479) );
  AOI221_X1 U31041 ( .B1(n39606), .B2(n33003), .C1(n39600), .C2(n32955), .A(
        n34224), .ZN(n34219) );
  OAI222_X1 U31042 ( .A1(n30761), .A2(n39594), .B1(n30825), .B2(n39588), .C1(
        n30697), .C2(n39582), .ZN(n34224) );
  AOI221_X1 U31043 ( .B1(n39354), .B2(n33003), .C1(n39348), .C2(n32955), .A(
        n35498), .ZN(n35493) );
  OAI222_X1 U31044 ( .A1(n30761), .A2(n39342), .B1(n30825), .B2(n39336), .C1(
        n30697), .C2(n39330), .ZN(n35498) );
  AOI221_X1 U31045 ( .B1(n39605), .B2(n33002), .C1(n39599), .C2(n32954), .A(
        n34243), .ZN(n34238) );
  OAI222_X1 U31046 ( .A1(n30760), .A2(n39593), .B1(n30824), .B2(n39587), .C1(
        n30696), .C2(n39581), .ZN(n34243) );
  AOI221_X1 U31047 ( .B1(n39353), .B2(n33002), .C1(n39347), .C2(n32954), .A(
        n35517), .ZN(n35512) );
  OAI222_X1 U31048 ( .A1(n30760), .A2(n39341), .B1(n30824), .B2(n39335), .C1(
        n30696), .C2(n39329), .ZN(n35517) );
  AOI221_X1 U31049 ( .B1(n39605), .B2(n33001), .C1(n39599), .C2(n32953), .A(
        n34262), .ZN(n34257) );
  OAI222_X1 U31050 ( .A1(n30759), .A2(n39593), .B1(n30823), .B2(n39587), .C1(
        n30695), .C2(n39581), .ZN(n34262) );
  AOI221_X1 U31051 ( .B1(n39353), .B2(n33001), .C1(n39347), .C2(n32953), .A(
        n35536), .ZN(n35531) );
  OAI222_X1 U31052 ( .A1(n30759), .A2(n39341), .B1(n30823), .B2(n39335), .C1(
        n30695), .C2(n39329), .ZN(n35536) );
  AOI221_X1 U31053 ( .B1(n39605), .B2(n33000), .C1(n39599), .C2(n32952), .A(
        n34281), .ZN(n34276) );
  OAI222_X1 U31054 ( .A1(n30758), .A2(n39593), .B1(n30822), .B2(n39587), .C1(
        n30694), .C2(n39581), .ZN(n34281) );
  AOI221_X1 U31055 ( .B1(n39353), .B2(n33000), .C1(n39347), .C2(n32952), .A(
        n35555), .ZN(n35550) );
  OAI222_X1 U31056 ( .A1(n30758), .A2(n39341), .B1(n30822), .B2(n39335), .C1(
        n30694), .C2(n39329), .ZN(n35555) );
  AOI221_X1 U31057 ( .B1(n39605), .B2(n32999), .C1(n39599), .C2(n32951), .A(
        n34300), .ZN(n34295) );
  OAI222_X1 U31058 ( .A1(n30757), .A2(n39593), .B1(n30821), .B2(n39587), .C1(
        n30693), .C2(n39581), .ZN(n34300) );
  AOI221_X1 U31059 ( .B1(n39353), .B2(n32999), .C1(n39347), .C2(n32951), .A(
        n35574), .ZN(n35569) );
  OAI222_X1 U31060 ( .A1(n30757), .A2(n39341), .B1(n30821), .B2(n39335), .C1(
        n30693), .C2(n39329), .ZN(n35574) );
  AOI221_X1 U31061 ( .B1(n39605), .B2(n32998), .C1(n39599), .C2(n32950), .A(
        n34319), .ZN(n34314) );
  OAI222_X1 U31062 ( .A1(n30756), .A2(n39593), .B1(n30820), .B2(n39587), .C1(
        n30692), .C2(n39581), .ZN(n34319) );
  AOI221_X1 U31063 ( .B1(n39353), .B2(n32998), .C1(n39347), .C2(n32950), .A(
        n35593), .ZN(n35588) );
  OAI222_X1 U31064 ( .A1(n30756), .A2(n39341), .B1(n30820), .B2(n39335), .C1(
        n30692), .C2(n39329), .ZN(n35593) );
  AOI221_X1 U31065 ( .B1(n39605), .B2(n32997), .C1(n39599), .C2(n32949), .A(
        n34338), .ZN(n34333) );
  OAI222_X1 U31066 ( .A1(n30755), .A2(n39593), .B1(n30819), .B2(n39587), .C1(
        n30691), .C2(n39581), .ZN(n34338) );
  AOI221_X1 U31067 ( .B1(n39353), .B2(n32997), .C1(n39347), .C2(n32949), .A(
        n35612), .ZN(n35607) );
  OAI222_X1 U31068 ( .A1(n30755), .A2(n39341), .B1(n30819), .B2(n39335), .C1(
        n30691), .C2(n39329), .ZN(n35612) );
  AOI221_X1 U31069 ( .B1(n39605), .B2(n32996), .C1(n39599), .C2(n32948), .A(
        n34357), .ZN(n34352) );
  OAI222_X1 U31070 ( .A1(n30754), .A2(n39593), .B1(n30818), .B2(n39587), .C1(
        n30690), .C2(n39581), .ZN(n34357) );
  AOI221_X1 U31071 ( .B1(n39353), .B2(n32996), .C1(n39347), .C2(n32948), .A(
        n35631), .ZN(n35626) );
  OAI222_X1 U31072 ( .A1(n30754), .A2(n39341), .B1(n30818), .B2(n39335), .C1(
        n30690), .C2(n39329), .ZN(n35631) );
  AOI221_X1 U31073 ( .B1(n39605), .B2(n32995), .C1(n39599), .C2(n32947), .A(
        n34376), .ZN(n34371) );
  OAI222_X1 U31074 ( .A1(n30753), .A2(n39593), .B1(n30817), .B2(n39587), .C1(
        n30689), .C2(n39581), .ZN(n34376) );
  AOI221_X1 U31075 ( .B1(n39353), .B2(n32995), .C1(n39347), .C2(n32947), .A(
        n35650), .ZN(n35645) );
  OAI222_X1 U31076 ( .A1(n30753), .A2(n39341), .B1(n30817), .B2(n39335), .C1(
        n30689), .C2(n39329), .ZN(n35650) );
  AOI221_X1 U31077 ( .B1(n39605), .B2(n32994), .C1(n39599), .C2(n32946), .A(
        n34395), .ZN(n34390) );
  OAI222_X1 U31078 ( .A1(n30752), .A2(n39593), .B1(n30816), .B2(n39587), .C1(
        n30688), .C2(n39581), .ZN(n34395) );
  AOI221_X1 U31079 ( .B1(n39353), .B2(n32994), .C1(n39347), .C2(n32946), .A(
        n35669), .ZN(n35664) );
  OAI222_X1 U31080 ( .A1(n30752), .A2(n39341), .B1(n30816), .B2(n39335), .C1(
        n30688), .C2(n39329), .ZN(n35669) );
  AOI221_X1 U31081 ( .B1(n39605), .B2(n32993), .C1(n39599), .C2(n32945), .A(
        n34414), .ZN(n34409) );
  OAI222_X1 U31082 ( .A1(n30751), .A2(n39593), .B1(n30815), .B2(n39587), .C1(
        n30687), .C2(n39581), .ZN(n34414) );
  AOI221_X1 U31083 ( .B1(n39353), .B2(n32993), .C1(n39347), .C2(n32945), .A(
        n35688), .ZN(n35683) );
  OAI222_X1 U31084 ( .A1(n30751), .A2(n39341), .B1(n30815), .B2(n39335), .C1(
        n30687), .C2(n39329), .ZN(n35688) );
  AOI221_X1 U31085 ( .B1(n39605), .B2(n32992), .C1(n39599), .C2(n32944), .A(
        n34433), .ZN(n34428) );
  OAI222_X1 U31086 ( .A1(n30750), .A2(n39593), .B1(n30814), .B2(n39587), .C1(
        n30686), .C2(n39581), .ZN(n34433) );
  AOI221_X1 U31087 ( .B1(n39353), .B2(n32992), .C1(n39347), .C2(n32944), .A(
        n35707), .ZN(n35702) );
  OAI222_X1 U31088 ( .A1(n30750), .A2(n39341), .B1(n30814), .B2(n39335), .C1(
        n30686), .C2(n39329), .ZN(n35707) );
  AOI221_X1 U31089 ( .B1(n39605), .B2(n32991), .C1(n39599), .C2(n32943), .A(
        n34452), .ZN(n34447) );
  OAI222_X1 U31090 ( .A1(n30749), .A2(n39593), .B1(n30813), .B2(n39587), .C1(
        n30685), .C2(n39581), .ZN(n34452) );
  AOI221_X1 U31091 ( .B1(n39353), .B2(n32991), .C1(n39347), .C2(n32943), .A(
        n35726), .ZN(n35721) );
  OAI222_X1 U31092 ( .A1(n30749), .A2(n39341), .B1(n30813), .B2(n39335), .C1(
        n30685), .C2(n39329), .ZN(n35726) );
  AOI221_X1 U31093 ( .B1(n39604), .B2(n33134), .C1(n39598), .C2(n33122), .A(
        n34471), .ZN(n34466) );
  OAI222_X1 U31094 ( .A1(n30748), .A2(n39592), .B1(n30812), .B2(n39586), .C1(
        n30684), .C2(n39580), .ZN(n34471) );
  AOI221_X1 U31095 ( .B1(n39352), .B2(n33134), .C1(n39346), .C2(n33122), .A(
        n35745), .ZN(n35740) );
  OAI222_X1 U31096 ( .A1(n30748), .A2(n39340), .B1(n30812), .B2(n39334), .C1(
        n30684), .C2(n39328), .ZN(n35745) );
  AOI221_X1 U31097 ( .B1(n39604), .B2(n33133), .C1(n39598), .C2(n33121), .A(
        n34490), .ZN(n34485) );
  OAI222_X1 U31098 ( .A1(n30747), .A2(n39592), .B1(n30811), .B2(n39586), .C1(
        n30683), .C2(n39580), .ZN(n34490) );
  AOI221_X1 U31099 ( .B1(n39352), .B2(n33133), .C1(n39346), .C2(n33121), .A(
        n35764), .ZN(n35759) );
  OAI222_X1 U31100 ( .A1(n30747), .A2(n39340), .B1(n30811), .B2(n39334), .C1(
        n30683), .C2(n39328), .ZN(n35764) );
  AOI221_X1 U31101 ( .B1(n39604), .B2(n33132), .C1(n39598), .C2(n33120), .A(
        n34509), .ZN(n34504) );
  OAI222_X1 U31102 ( .A1(n30746), .A2(n39592), .B1(n30810), .B2(n39586), .C1(
        n30682), .C2(n39580), .ZN(n34509) );
  AOI221_X1 U31103 ( .B1(n39352), .B2(n33132), .C1(n39346), .C2(n33120), .A(
        n35783), .ZN(n35778) );
  OAI222_X1 U31104 ( .A1(n30746), .A2(n39340), .B1(n30810), .B2(n39334), .C1(
        n30682), .C2(n39328), .ZN(n35783) );
  AOI221_X1 U31105 ( .B1(n39604), .B2(n33131), .C1(n39598), .C2(n33119), .A(
        n34528), .ZN(n34523) );
  OAI222_X1 U31106 ( .A1(n30745), .A2(n39592), .B1(n30809), .B2(n39586), .C1(
        n30681), .C2(n39580), .ZN(n34528) );
  AOI221_X1 U31107 ( .B1(n39352), .B2(n33131), .C1(n39346), .C2(n33119), .A(
        n35802), .ZN(n35797) );
  OAI222_X1 U31108 ( .A1(n30745), .A2(n39340), .B1(n30809), .B2(n39334), .C1(
        n30681), .C2(n39328), .ZN(n35802) );
  AOI221_X1 U31109 ( .B1(n39604), .B2(n33130), .C1(n39598), .C2(n33118), .A(
        n34547), .ZN(n34542) );
  OAI222_X1 U31110 ( .A1(n30744), .A2(n39592), .B1(n30808), .B2(n39586), .C1(
        n30680), .C2(n39580), .ZN(n34547) );
  AOI221_X1 U31111 ( .B1(n39352), .B2(n33130), .C1(n39346), .C2(n33118), .A(
        n35821), .ZN(n35816) );
  OAI222_X1 U31112 ( .A1(n30744), .A2(n39340), .B1(n30808), .B2(n39334), .C1(
        n30680), .C2(n39328), .ZN(n35821) );
  AOI221_X1 U31113 ( .B1(n39604), .B2(n33129), .C1(n39598), .C2(n33117), .A(
        n34566), .ZN(n34561) );
  OAI222_X1 U31114 ( .A1(n30743), .A2(n39592), .B1(n30807), .B2(n39586), .C1(
        n30679), .C2(n39580), .ZN(n34566) );
  AOI221_X1 U31115 ( .B1(n39352), .B2(n33129), .C1(n39346), .C2(n33117), .A(
        n35840), .ZN(n35835) );
  OAI222_X1 U31116 ( .A1(n30743), .A2(n39340), .B1(n30807), .B2(n39334), .C1(
        n30679), .C2(n39328), .ZN(n35840) );
  AOI221_X1 U31117 ( .B1(n39604), .B2(n33128), .C1(n39598), .C2(n33116), .A(
        n34585), .ZN(n34580) );
  OAI222_X1 U31118 ( .A1(n30742), .A2(n39592), .B1(n30806), .B2(n39586), .C1(
        n30678), .C2(n39580), .ZN(n34585) );
  AOI221_X1 U31119 ( .B1(n39352), .B2(n33128), .C1(n39346), .C2(n33116), .A(
        n35859), .ZN(n35854) );
  OAI222_X1 U31120 ( .A1(n30742), .A2(n39340), .B1(n30806), .B2(n39334), .C1(
        n30678), .C2(n39328), .ZN(n35859) );
  AOI221_X1 U31121 ( .B1(n39604), .B2(n33127), .C1(n39598), .C2(n33115), .A(
        n34604), .ZN(n34599) );
  OAI222_X1 U31122 ( .A1(n30741), .A2(n39592), .B1(n30805), .B2(n39586), .C1(
        n30677), .C2(n39580), .ZN(n34604) );
  AOI221_X1 U31123 ( .B1(n39352), .B2(n33127), .C1(n39346), .C2(n33115), .A(
        n35878), .ZN(n35873) );
  OAI222_X1 U31124 ( .A1(n30741), .A2(n39340), .B1(n30805), .B2(n39334), .C1(
        n30677), .C2(n39328), .ZN(n35878) );
  AOI221_X1 U31125 ( .B1(n39604), .B2(n33126), .C1(n39598), .C2(n33114), .A(
        n34623), .ZN(n34618) );
  OAI222_X1 U31126 ( .A1(n30740), .A2(n39592), .B1(n30804), .B2(n39586), .C1(
        n30676), .C2(n39580), .ZN(n34623) );
  AOI221_X1 U31127 ( .B1(n39352), .B2(n33126), .C1(n39346), .C2(n33114), .A(
        n35897), .ZN(n35892) );
  OAI222_X1 U31128 ( .A1(n30740), .A2(n39340), .B1(n30804), .B2(n39334), .C1(
        n30676), .C2(n39328), .ZN(n35897) );
  AOI221_X1 U31129 ( .B1(n39604), .B2(n33125), .C1(n39598), .C2(n33113), .A(
        n34642), .ZN(n34637) );
  OAI222_X1 U31130 ( .A1(n30739), .A2(n39592), .B1(n30803), .B2(n39586), .C1(
        n30675), .C2(n39580), .ZN(n34642) );
  AOI221_X1 U31131 ( .B1(n39352), .B2(n33125), .C1(n39346), .C2(n33113), .A(
        n35916), .ZN(n35911) );
  OAI222_X1 U31132 ( .A1(n30739), .A2(n39340), .B1(n30803), .B2(n39334), .C1(
        n30675), .C2(n39328), .ZN(n35916) );
  AOI221_X1 U31133 ( .B1(n39604), .B2(n33124), .C1(n39598), .C2(n33112), .A(
        n34661), .ZN(n34656) );
  OAI222_X1 U31134 ( .A1(n30738), .A2(n39592), .B1(n30802), .B2(n39586), .C1(
        n30674), .C2(n39580), .ZN(n34661) );
  AOI221_X1 U31135 ( .B1(n39352), .B2(n33124), .C1(n39346), .C2(n33112), .A(
        n35935), .ZN(n35930) );
  OAI222_X1 U31136 ( .A1(n30738), .A2(n39340), .B1(n30802), .B2(n39334), .C1(
        n30674), .C2(n39328), .ZN(n35935) );
  AOI221_X1 U31137 ( .B1(n39604), .B2(n33123), .C1(n39598), .C2(n33111), .A(
        n34692), .ZN(n34686) );
  OAI222_X1 U31138 ( .A1(n30737), .A2(n39592), .B1(n30801), .B2(n39586), .C1(
        n30673), .C2(n39580), .ZN(n34692) );
  AOI221_X1 U31139 ( .B1(n39352), .B2(n33123), .C1(n39346), .C2(n33111), .A(
        n35966), .ZN(n35960) );
  OAI222_X1 U31140 ( .A1(n30737), .A2(n39340), .B1(n30801), .B2(n39334), .C1(
        n30673), .C2(n39328), .ZN(n35966) );
  NAND2_X1 U31141 ( .A1(n33330), .A2(n33294), .ZN(n33394) );
  AND2_X1 U31142 ( .A1(N6273), .A2(n32164), .ZN(n34684) );
  AND2_X1 U31143 ( .A1(N6398), .A2(n32169), .ZN(n35958) );
  INV_X1 U31144 ( .A(n33398), .ZN(n32254) );
  AND2_X1 U31145 ( .A1(N6272), .A2(N6273), .ZN(n34681) );
  AND2_X1 U31146 ( .A1(N6397), .A2(N6398), .ZN(n35955) );
  INV_X1 U31147 ( .A(n34694), .ZN(n32168) );
  INV_X1 U31148 ( .A(n35968), .ZN(n32173) );
  AND3_X1 U31149 ( .A1(N931), .A2(n32151), .A3(n33331), .ZN(n33367) );
  AND3_X1 U31150 ( .A1(N932), .A2(N931), .A3(n33331), .ZN(n33306) );
  AND3_X1 U31151 ( .A1(N932), .A2(n32152), .A3(n33331), .ZN(n33338) );
  AND3_X1 U31152 ( .A1(n33294), .A2(n32150), .A3(n33300), .ZN(n33257) );
  INV_X1 U31153 ( .A(n33402), .ZN(n32163) );
  INV_X1 U31154 ( .A(N689), .ZN(n32248) );
  INV_X1 U31155 ( .A(N6271), .ZN(n32165) );
  INV_X1 U31156 ( .A(N6396), .ZN(n32170) );
  INV_X1 U31157 ( .A(N688), .ZN(n32251) );
  INV_X1 U31158 ( .A(N6270), .ZN(n32166) );
  INV_X1 U31159 ( .A(N6395), .ZN(n32171) );
  BUF_X1 U31160 ( .A(n33272), .Z(n40522) );
  OAI211_X1 U31161 ( .C1(n33256), .C2(n33274), .A(n40521), .B(n41368), .ZN(
        n33272) );
  BUF_X1 U31162 ( .A(n33277), .Z(n40502) );
  OAI211_X1 U31163 ( .C1(n33256), .C2(n32157), .A(n40501), .B(n41367), .ZN(
        n33277) );
  BUF_X1 U31164 ( .A(n33262), .Z(n40562) );
  OAI211_X1 U31165 ( .C1(n33256), .C2(n33264), .A(n40561), .B(n41367), .ZN(
        n33262) );
  BUF_X1 U31166 ( .A(n33267), .Z(n40542) );
  OAI211_X1 U31167 ( .C1(n33256), .C2(n33269), .A(n40541), .B(n41368), .ZN(
        n33267) );
  BUF_X1 U31168 ( .A(n33282), .Z(n40482) );
  OAI211_X1 U31169 ( .C1(n33256), .C2(n32158), .A(n40481), .B(n41367), .ZN(
        n33282) );
  BUF_X1 U31170 ( .A(n33287), .Z(n40462) );
  OAI211_X1 U31171 ( .C1(n33256), .C2(n32159), .A(n40461), .B(n41367), .ZN(
        n33287) );
  BUF_X1 U31172 ( .A(n33292), .Z(n40442) );
  OAI211_X1 U31173 ( .C1(n33256), .C2(n32160), .A(n40441), .B(n41367), .ZN(
        n33292) );
  BUF_X1 U31174 ( .A(n33253), .Z(n40582) );
  OAI211_X1 U31175 ( .C1(n33255), .C2(n33256), .A(n40581), .B(n41367), .ZN(
        n33253) );
  INV_X1 U31176 ( .A(N929), .ZN(n32161) );
  INV_X1 U31177 ( .A(n37240), .ZN(n32243) );
  AND2_X1 U31178 ( .A1(n33301), .A2(n33299), .ZN(n33333) );
  INV_X1 U31179 ( .A(N931), .ZN(n32152) );
  INV_X1 U31180 ( .A(N932), .ZN(n32151) );
  INV_X1 U31181 ( .A(N812), .ZN(n32249) );
  AND2_X1 U31182 ( .A1(n33301), .A2(n33300), .ZN(n33331) );
  INV_X1 U31183 ( .A(n33362), .ZN(n32239) );
  INV_X1 U31184 ( .A(N690), .ZN(n32246) );
  INV_X1 U31185 ( .A(N6272), .ZN(n32164) );
  INV_X1 U31186 ( .A(N6397), .ZN(n32169) );
  INV_X1 U31187 ( .A(N813), .ZN(n32247) );
  NAND2_X1 U31188 ( .A1(\add_136/carry[4] ), .A2(n32242), .ZN(n37251) );
  NOR3_X1 U31189 ( .A1(n33223), .A2(n32075), .A3(n33222), .ZN(n33224) );
  INV_X1 U31190 ( .A(n39297), .ZN(n39295) );
  INV_X1 U31191 ( .A(n39297), .ZN(n39294) );
  INV_X1 U31192 ( .A(n39297), .ZN(n39296) );
  OAI21_X1 U31193 ( .B1(n33230), .B2(n33231), .A(n33232), .ZN(n33225) );
  AND3_X1 U31194 ( .A1(n33233), .A2(n41370), .A3(n33237), .ZN(n33249) );
  AND3_X1 U31195 ( .A1(n33211), .A2(n33212), .A3(n33213), .ZN(n33210) );
  NAND4_X1 U31196 ( .A1(n33218), .A2(n33212), .A3(n41367), .A4(n32083), .ZN(
        n33211) );
  OAI21_X1 U31197 ( .B1(n33216), .B2(N659), .A(n33245), .ZN(n33244) );
  NAND4_X1 U31198 ( .A1(n32241), .A2(n33239), .A3(n33245), .A4(n33218), .ZN(
        n35977) );
  INV_X1 U31199 ( .A(n33238), .ZN(n32241) );
  NAND4_X1 U31200 ( .A1(n32323), .A2(n32322), .A3(n32260), .A4(n32258), .ZN(
        n35976) );
  INV_X1 U31201 ( .A(n33233), .ZN(n32077) );
  OAI21_X1 U31202 ( .B1(n32322), .B2(n33225), .A(n33226), .ZN(n9896) );
  OAI21_X1 U31203 ( .B1(n33222), .B2(n33223), .A(n32322), .ZN(n33226) );
  NOR2_X1 U31204 ( .A1(n33224), .A2(n32260), .ZN(n9899) );
  NOR2_X1 U31205 ( .A1(n33224), .A2(n32258), .ZN(n9897) );
  INV_X1 U31206 ( .A(n33234), .ZN(n32076) );
  BUF_X1 U31207 ( .A(n32079), .Z(n41368) );
  BUF_X1 U31208 ( .A(n32079), .Z(n41369) );
  BUF_X1 U31209 ( .A(n32079), .Z(n41370) );
  BUF_X1 U31210 ( .A(n32079), .Z(n41367) );
  BUF_X1 U31211 ( .A(n32079), .Z(n41364) );
  BUF_X1 U31212 ( .A(n32079), .Z(n41366) );
  BUF_X1 U31213 ( .A(n32079), .Z(n41365) );
  BUF_X1 U31214 ( .A(n33424), .Z(n39796) );
  BUF_X1 U31215 ( .A(n34698), .Z(n39544) );
  BUF_X1 U31216 ( .A(n33424), .Z(n39800) );
  BUF_X1 U31217 ( .A(n34698), .Z(n39548) );
  BUF_X1 U31218 ( .A(n33424), .Z(n39799) );
  BUF_X1 U31219 ( .A(n34698), .Z(n39547) );
  BUF_X1 U31220 ( .A(n33424), .Z(n39798) );
  BUF_X1 U31221 ( .A(n34698), .Z(n39546) );
  BUF_X1 U31222 ( .A(n33424), .Z(n39797) );
  BUF_X1 U31223 ( .A(n34698), .Z(n39545) );
  INV_X1 U31224 ( .A(n33208), .ZN(n32167) );
  INV_X1 U31225 ( .A(n33207), .ZN(n32172) );
  INV_X1 U31226 ( .A(n33209), .ZN(n32162) );
  BUF_X1 U31227 ( .A(n32124), .Z(n41118) );
  BUF_X1 U31228 ( .A(n32214), .Z(n40734) );
  BUF_X1 U31229 ( .A(n32123), .Z(n41124) );
  BUF_X1 U31230 ( .A(n32213), .Z(n40740) );
  BUF_X1 U31231 ( .A(n32122), .Z(n41130) );
  BUF_X1 U31232 ( .A(n32212), .Z(n40746) );
  BUF_X1 U31233 ( .A(n32121), .Z(n41136) );
  BUF_X1 U31234 ( .A(n32211), .Z(n40752) );
  BUF_X1 U31235 ( .A(n32120), .Z(n41142) );
  BUF_X1 U31236 ( .A(n32210), .Z(n40758) );
  BUF_X1 U31237 ( .A(n32119), .Z(n41148) );
  BUF_X1 U31238 ( .A(n32209), .Z(n40764) );
  BUF_X1 U31239 ( .A(n32118), .Z(n41154) );
  BUF_X1 U31240 ( .A(n32208), .Z(n40770) );
  BUF_X1 U31241 ( .A(n32117), .Z(n41160) );
  BUF_X1 U31242 ( .A(n32207), .Z(n40776) );
  BUF_X1 U31243 ( .A(n32116), .Z(n41166) );
  BUF_X1 U31244 ( .A(n32206), .Z(n40782) );
  BUF_X1 U31245 ( .A(n32115), .Z(n41172) );
  BUF_X1 U31246 ( .A(n32205), .Z(n40788) );
  BUF_X1 U31247 ( .A(n32114), .Z(n41178) );
  BUF_X1 U31248 ( .A(n32204), .Z(n40794) );
  BUF_X1 U31249 ( .A(n32113), .Z(n41184) );
  BUF_X1 U31250 ( .A(n32203), .Z(n40800) );
  BUF_X1 U31251 ( .A(n32112), .Z(n41190) );
  BUF_X1 U31252 ( .A(n32202), .Z(n40806) );
  BUF_X1 U31253 ( .A(n32111), .Z(n41196) );
  BUF_X1 U31254 ( .A(n32201), .Z(n40812) );
  BUF_X1 U31255 ( .A(n32110), .Z(n41202) );
  BUF_X1 U31256 ( .A(n32200), .Z(n40818) );
  BUF_X1 U31257 ( .A(n32109), .Z(n41208) );
  BUF_X1 U31258 ( .A(n32199), .Z(n40824) );
  BUF_X1 U31259 ( .A(n32108), .Z(n41214) );
  BUF_X1 U31260 ( .A(n32198), .Z(n40830) );
  BUF_X1 U31261 ( .A(n32107), .Z(n41220) );
  BUF_X1 U31262 ( .A(n32197), .Z(n40836) );
  BUF_X1 U31263 ( .A(n32106), .Z(n41226) );
  BUF_X1 U31264 ( .A(n32196), .Z(n40842) );
  BUF_X1 U31265 ( .A(n32105), .Z(n41232) );
  BUF_X1 U31266 ( .A(n32195), .Z(n40848) );
  BUF_X1 U31267 ( .A(n32104), .Z(n41238) );
  BUF_X1 U31268 ( .A(n32194), .Z(n40854) );
  BUF_X1 U31269 ( .A(n32103), .Z(n41244) );
  BUF_X1 U31270 ( .A(n32193), .Z(n40860) );
  BUF_X1 U31271 ( .A(n32102), .Z(n41250) );
  BUF_X1 U31272 ( .A(n32192), .Z(n40866) );
  BUF_X1 U31273 ( .A(n32101), .Z(n41256) );
  BUF_X1 U31274 ( .A(n32191), .Z(n40872) );
  BUF_X1 U31275 ( .A(n32100), .Z(n41262) );
  BUF_X1 U31276 ( .A(n32190), .Z(n40878) );
  BUF_X1 U31277 ( .A(n32099), .Z(n41268) );
  BUF_X1 U31278 ( .A(n32189), .Z(n40884) );
  BUF_X1 U31279 ( .A(n32098), .Z(n41274) );
  BUF_X1 U31280 ( .A(n32188), .Z(n40890) );
  BUF_X1 U31281 ( .A(n32097), .Z(n41280) );
  BUF_X1 U31282 ( .A(n32187), .Z(n40896) );
  BUF_X1 U31283 ( .A(n32096), .Z(n41286) );
  BUF_X1 U31284 ( .A(n32186), .Z(n40902) );
  BUF_X1 U31285 ( .A(n32095), .Z(n41292) );
  BUF_X1 U31286 ( .A(n32185), .Z(n40908) );
  BUF_X1 U31287 ( .A(n32094), .Z(n41298) );
  BUF_X1 U31288 ( .A(n32184), .Z(n40914) );
  BUF_X1 U31289 ( .A(n32093), .Z(n41304) );
  BUF_X1 U31290 ( .A(n32183), .Z(n40920) );
  BUF_X1 U31291 ( .A(n32092), .Z(n41310) );
  BUF_X1 U31292 ( .A(n32182), .Z(n40926) );
  BUF_X1 U31293 ( .A(n32091), .Z(n41316) );
  BUF_X1 U31294 ( .A(n32181), .Z(n40932) );
  BUF_X1 U31295 ( .A(n32090), .Z(n41322) );
  BUF_X1 U31296 ( .A(n32180), .Z(n40938) );
  BUF_X1 U31297 ( .A(n32089), .Z(n41328) );
  BUF_X1 U31298 ( .A(n32179), .Z(n40944) );
  BUF_X1 U31299 ( .A(n32088), .Z(n41334) );
  BUF_X1 U31300 ( .A(n32178), .Z(n40950) );
  BUF_X1 U31301 ( .A(n32087), .Z(n41340) );
  BUF_X1 U31302 ( .A(n32177), .Z(n40956) );
  BUF_X1 U31303 ( .A(n32086), .Z(n41346) );
  BUF_X1 U31304 ( .A(n32176), .Z(n40962) );
  BUF_X1 U31305 ( .A(n32085), .Z(n41352) );
  BUF_X1 U31306 ( .A(n32175), .Z(n40968) );
  BUF_X1 U31307 ( .A(n32084), .Z(n41358) );
  BUF_X1 U31308 ( .A(n32174), .Z(n40974) );
  BUF_X1 U31309 ( .A(n32147), .Z(n40980) );
  BUF_X1 U31310 ( .A(n32237), .Z(n40596) );
  BUF_X1 U31311 ( .A(n32146), .Z(n40986) );
  BUF_X1 U31312 ( .A(n32236), .Z(n40602) );
  BUF_X1 U31313 ( .A(n32145), .Z(n40992) );
  BUF_X1 U31314 ( .A(n32235), .Z(n40608) );
  BUF_X1 U31315 ( .A(n32144), .Z(n40998) );
  BUF_X1 U31316 ( .A(n32234), .Z(n40614) );
  BUF_X1 U31317 ( .A(n32143), .Z(n41004) );
  BUF_X1 U31318 ( .A(n32233), .Z(n40620) );
  BUF_X1 U31319 ( .A(n32142), .Z(n41010) );
  BUF_X1 U31320 ( .A(n32232), .Z(n40626) );
  BUF_X1 U31321 ( .A(n32141), .Z(n41016) );
  BUF_X1 U31322 ( .A(n32231), .Z(n40632) );
  BUF_X1 U31323 ( .A(n32140), .Z(n41022) );
  BUF_X1 U31324 ( .A(n32230), .Z(n40638) );
  BUF_X1 U31325 ( .A(n32139), .Z(n41028) );
  BUF_X1 U31326 ( .A(n32229), .Z(n40644) );
  BUF_X1 U31327 ( .A(n32138), .Z(n41034) );
  BUF_X1 U31328 ( .A(n32228), .Z(n40650) );
  BUF_X1 U31329 ( .A(n32137), .Z(n41040) );
  BUF_X1 U31330 ( .A(n32227), .Z(n40656) );
  BUF_X1 U31331 ( .A(n32136), .Z(n41046) );
  BUF_X1 U31332 ( .A(n32226), .Z(n40662) );
  BUF_X1 U31333 ( .A(n32135), .Z(n41052) );
  BUF_X1 U31334 ( .A(n32225), .Z(n40668) );
  BUF_X1 U31335 ( .A(n32134), .Z(n41058) );
  BUF_X1 U31336 ( .A(n32224), .Z(n40674) );
  BUF_X1 U31337 ( .A(n32133), .Z(n41064) );
  BUF_X1 U31338 ( .A(n32223), .Z(n40680) );
  BUF_X1 U31339 ( .A(n32132), .Z(n41070) );
  BUF_X1 U31340 ( .A(n32222), .Z(n40686) );
  BUF_X1 U31341 ( .A(n32131), .Z(n41076) );
  BUF_X1 U31342 ( .A(n32221), .Z(n40692) );
  BUF_X1 U31343 ( .A(n32130), .Z(n41082) );
  BUF_X1 U31344 ( .A(n32220), .Z(n40698) );
  BUF_X1 U31345 ( .A(n32129), .Z(n41088) );
  BUF_X1 U31346 ( .A(n32219), .Z(n40704) );
  BUF_X1 U31347 ( .A(n32128), .Z(n41094) );
  BUF_X1 U31348 ( .A(n32218), .Z(n40710) );
  BUF_X1 U31349 ( .A(n32127), .Z(n41100) );
  BUF_X1 U31350 ( .A(n32217), .Z(n40716) );
  BUF_X1 U31351 ( .A(n32126), .Z(n41106) );
  BUF_X1 U31352 ( .A(n32216), .Z(n40722) );
  BUF_X1 U31353 ( .A(n32125), .Z(n41112) );
  BUF_X1 U31354 ( .A(n32215), .Z(n40728) );
  BUF_X1 U31355 ( .A(n32147), .Z(n40981) );
  BUF_X1 U31356 ( .A(n32237), .Z(n40597) );
  BUF_X1 U31357 ( .A(n32146), .Z(n40987) );
  BUF_X1 U31358 ( .A(n32236), .Z(n40603) );
  BUF_X1 U31359 ( .A(n32145), .Z(n40993) );
  BUF_X1 U31360 ( .A(n32235), .Z(n40609) );
  BUF_X1 U31361 ( .A(n32144), .Z(n40999) );
  BUF_X1 U31362 ( .A(n32234), .Z(n40615) );
  BUF_X1 U31363 ( .A(n32143), .Z(n41005) );
  BUF_X1 U31364 ( .A(n32233), .Z(n40621) );
  BUF_X1 U31365 ( .A(n32142), .Z(n41011) );
  BUF_X1 U31366 ( .A(n32232), .Z(n40627) );
  BUF_X1 U31367 ( .A(n32141), .Z(n41017) );
  BUF_X1 U31368 ( .A(n32231), .Z(n40633) );
  BUF_X1 U31369 ( .A(n32140), .Z(n41023) );
  BUF_X1 U31370 ( .A(n32230), .Z(n40639) );
  BUF_X1 U31371 ( .A(n32139), .Z(n41029) );
  BUF_X1 U31372 ( .A(n32229), .Z(n40645) );
  BUF_X1 U31373 ( .A(n32138), .Z(n41035) );
  BUF_X1 U31374 ( .A(n32228), .Z(n40651) );
  BUF_X1 U31375 ( .A(n32137), .Z(n41041) );
  BUF_X1 U31376 ( .A(n32227), .Z(n40657) );
  BUF_X1 U31377 ( .A(n32136), .Z(n41047) );
  BUF_X1 U31378 ( .A(n32226), .Z(n40663) );
  BUF_X1 U31379 ( .A(n32135), .Z(n41053) );
  BUF_X1 U31380 ( .A(n32225), .Z(n40669) );
  BUF_X1 U31381 ( .A(n32134), .Z(n41059) );
  BUF_X1 U31382 ( .A(n32224), .Z(n40675) );
  BUF_X1 U31383 ( .A(n32133), .Z(n41065) );
  BUF_X1 U31384 ( .A(n32223), .Z(n40681) );
  BUF_X1 U31385 ( .A(n32132), .Z(n41071) );
  BUF_X1 U31386 ( .A(n32222), .Z(n40687) );
  BUF_X1 U31387 ( .A(n32131), .Z(n41077) );
  BUF_X1 U31388 ( .A(n32221), .Z(n40693) );
  BUF_X1 U31389 ( .A(n32130), .Z(n41083) );
  BUF_X1 U31390 ( .A(n32220), .Z(n40699) );
  BUF_X1 U31391 ( .A(n32129), .Z(n41089) );
  BUF_X1 U31392 ( .A(n32219), .Z(n40705) );
  BUF_X1 U31393 ( .A(n32128), .Z(n41095) );
  BUF_X1 U31394 ( .A(n32218), .Z(n40711) );
  BUF_X1 U31395 ( .A(n32127), .Z(n41101) );
  BUF_X1 U31396 ( .A(n32217), .Z(n40717) );
  BUF_X1 U31397 ( .A(n32126), .Z(n41107) );
  BUF_X1 U31398 ( .A(n32216), .Z(n40723) );
  BUF_X1 U31399 ( .A(n32125), .Z(n41113) );
  BUF_X1 U31400 ( .A(n32215), .Z(n40729) );
  BUF_X1 U31401 ( .A(n32124), .Z(n41119) );
  BUF_X1 U31402 ( .A(n32214), .Z(n40735) );
  BUF_X1 U31403 ( .A(n32123), .Z(n41125) );
  BUF_X1 U31404 ( .A(n32213), .Z(n40741) );
  BUF_X1 U31405 ( .A(n32122), .Z(n41131) );
  BUF_X1 U31406 ( .A(n32212), .Z(n40747) );
  BUF_X1 U31407 ( .A(n32121), .Z(n41137) );
  BUF_X1 U31408 ( .A(n32211), .Z(n40753) );
  BUF_X1 U31409 ( .A(n32120), .Z(n41143) );
  BUF_X1 U31410 ( .A(n32210), .Z(n40759) );
  BUF_X1 U31411 ( .A(n32119), .Z(n41149) );
  BUF_X1 U31412 ( .A(n32209), .Z(n40765) );
  BUF_X1 U31413 ( .A(n32118), .Z(n41155) );
  BUF_X1 U31414 ( .A(n32208), .Z(n40771) );
  BUF_X1 U31415 ( .A(n32117), .Z(n41161) );
  BUF_X1 U31416 ( .A(n32207), .Z(n40777) );
  BUF_X1 U31417 ( .A(n32116), .Z(n41167) );
  BUF_X1 U31418 ( .A(n32206), .Z(n40783) );
  BUF_X1 U31419 ( .A(n32115), .Z(n41173) );
  BUF_X1 U31420 ( .A(n32205), .Z(n40789) );
  BUF_X1 U31421 ( .A(n32114), .Z(n41179) );
  BUF_X1 U31422 ( .A(n32204), .Z(n40795) );
  BUF_X1 U31423 ( .A(n32113), .Z(n41185) );
  BUF_X1 U31424 ( .A(n32203), .Z(n40801) );
  BUF_X1 U31425 ( .A(n32112), .Z(n41191) );
  BUF_X1 U31426 ( .A(n32202), .Z(n40807) );
  BUF_X1 U31427 ( .A(n32111), .Z(n41197) );
  BUF_X1 U31428 ( .A(n32201), .Z(n40813) );
  BUF_X1 U31429 ( .A(n32110), .Z(n41203) );
  BUF_X1 U31430 ( .A(n32200), .Z(n40819) );
  BUF_X1 U31431 ( .A(n32109), .Z(n41209) );
  BUF_X1 U31432 ( .A(n32199), .Z(n40825) );
  BUF_X1 U31433 ( .A(n32108), .Z(n41215) );
  BUF_X1 U31434 ( .A(n32198), .Z(n40831) );
  BUF_X1 U31435 ( .A(n32107), .Z(n41221) );
  BUF_X1 U31436 ( .A(n32197), .Z(n40837) );
  BUF_X1 U31437 ( .A(n32106), .Z(n41227) );
  BUF_X1 U31438 ( .A(n32196), .Z(n40843) );
  BUF_X1 U31439 ( .A(n32105), .Z(n41233) );
  BUF_X1 U31440 ( .A(n32195), .Z(n40849) );
  BUF_X1 U31441 ( .A(n32104), .Z(n41239) );
  BUF_X1 U31442 ( .A(n32194), .Z(n40855) );
  BUF_X1 U31443 ( .A(n32103), .Z(n41245) );
  BUF_X1 U31444 ( .A(n32193), .Z(n40861) );
  BUF_X1 U31445 ( .A(n32102), .Z(n41251) );
  BUF_X1 U31446 ( .A(n32192), .Z(n40867) );
  BUF_X1 U31447 ( .A(n32101), .Z(n41257) );
  BUF_X1 U31448 ( .A(n32191), .Z(n40873) );
  BUF_X1 U31449 ( .A(n32100), .Z(n41263) );
  BUF_X1 U31450 ( .A(n32190), .Z(n40879) );
  BUF_X1 U31451 ( .A(n32099), .Z(n41269) );
  BUF_X1 U31452 ( .A(n32189), .Z(n40885) );
  BUF_X1 U31453 ( .A(n32098), .Z(n41275) );
  BUF_X1 U31454 ( .A(n32188), .Z(n40891) );
  BUF_X1 U31455 ( .A(n32097), .Z(n41281) );
  BUF_X1 U31456 ( .A(n32187), .Z(n40897) );
  BUF_X1 U31457 ( .A(n32096), .Z(n41287) );
  BUF_X1 U31458 ( .A(n32186), .Z(n40903) );
  BUF_X1 U31459 ( .A(n32095), .Z(n41293) );
  BUF_X1 U31460 ( .A(n32185), .Z(n40909) );
  BUF_X1 U31461 ( .A(n32094), .Z(n41299) );
  BUF_X1 U31462 ( .A(n32184), .Z(n40915) );
  BUF_X1 U31463 ( .A(n32093), .Z(n41305) );
  BUF_X1 U31464 ( .A(n32183), .Z(n40921) );
  BUF_X1 U31465 ( .A(n32092), .Z(n41311) );
  BUF_X1 U31466 ( .A(n32182), .Z(n40927) );
  BUF_X1 U31467 ( .A(n32091), .Z(n41317) );
  BUF_X1 U31468 ( .A(n32181), .Z(n40933) );
  BUF_X1 U31469 ( .A(n32090), .Z(n41323) );
  BUF_X1 U31470 ( .A(n32180), .Z(n40939) );
  BUF_X1 U31471 ( .A(n32089), .Z(n41329) );
  BUF_X1 U31472 ( .A(n32179), .Z(n40945) );
  BUF_X1 U31473 ( .A(n32088), .Z(n41335) );
  BUF_X1 U31474 ( .A(n32178), .Z(n40951) );
  BUF_X1 U31475 ( .A(n32087), .Z(n41341) );
  BUF_X1 U31476 ( .A(n32177), .Z(n40957) );
  BUF_X1 U31477 ( .A(n32086), .Z(n41347) );
  BUF_X1 U31478 ( .A(n32176), .Z(n40963) );
  BUF_X1 U31479 ( .A(n32085), .Z(n41353) );
  BUF_X1 U31480 ( .A(n32175), .Z(n40969) );
  BUF_X1 U31481 ( .A(n32084), .Z(n41359) );
  BUF_X1 U31482 ( .A(n32174), .Z(n40975) );
  NAND2_X1 U31483 ( .A1(n32253), .A2(n33208), .ZN(n34696) );
  NAND2_X1 U31484 ( .A1(n32253), .A2(n33207), .ZN(n35970) );
  NAND2_X1 U31485 ( .A1(n32253), .A2(n33209), .ZN(n33423) );
  NOR3_X1 U31486 ( .A1(n32239), .A2(n23853), .A3(N813), .ZN(n33298) );
  NOR2_X1 U31487 ( .A1(n2695), .A2(n32162), .ZN(\U3/U193/Z_4 ) );
  AOI221_X1 U31488 ( .B1(n39287), .B2(n30006), .C1(n39281), .C2(n30070), .A(
        n36085), .ZN(n36084) );
  OAI222_X1 U31489 ( .A1(n31994), .A2(n39275), .B1(n32286), .B2(n39269), .C1(
        n31934), .C2(n39263), .ZN(n36085) );
  AOI221_X1 U31490 ( .B1(n39287), .B2(n30005), .C1(n39281), .C2(n30069), .A(
        n36066), .ZN(n36065) );
  OAI222_X1 U31491 ( .A1(n31993), .A2(n39275), .B1(n32053), .B2(n39269), .C1(
        n31933), .C2(n39263), .ZN(n36066) );
  AOI221_X1 U31492 ( .B1(n39287), .B2(n30004), .C1(n39281), .C2(n30068), .A(
        n36047), .ZN(n36046) );
  OAI222_X1 U31493 ( .A1(n31992), .A2(n39275), .B1(n32052), .B2(n39269), .C1(
        n31932), .C2(n39263), .ZN(n36047) );
  AOI221_X1 U31494 ( .B1(n39287), .B2(n30003), .C1(n39281), .C2(n30067), .A(
        n35990), .ZN(n35987) );
  OAI222_X1 U31495 ( .A1(n31991), .A2(n39275), .B1(n32051), .B2(n39269), .C1(
        n31931), .C2(n39263), .ZN(n35990) );
  OAI222_X1 U31496 ( .A1(n40954), .A2(n40430), .B1(n41338), .B2(n40423), .C1(
        n40421), .C2(n33199), .ZN(n9319) );
  OAI222_X1 U31497 ( .A1(n40966), .A2(n40430), .B1(n41350), .B2(n40423), .C1(
        n40421), .C2(n33197), .ZN(n9317) );
  OAI222_X1 U31498 ( .A1(n40972), .A2(n40430), .B1(n41356), .B2(n40423), .C1(
        n40421), .C2(n33196), .ZN(n9316) );
  OAI222_X1 U31499 ( .A1(n40978), .A2(n40430), .B1(n41362), .B2(n40423), .C1(
        n40421), .C2(n33195), .ZN(n9315) );
  OAI222_X1 U31500 ( .A1(n40954), .A2(n40410), .B1(n41338), .B2(n40403), .C1(
        n40401), .C2(n33139), .ZN(n9255) );
  OAI222_X1 U31501 ( .A1(n40966), .A2(n40410), .B1(n41350), .B2(n40403), .C1(
        n40401), .C2(n33137), .ZN(n9253) );
  OAI222_X1 U31502 ( .A1(n40972), .A2(n40410), .B1(n41356), .B2(n40403), .C1(
        n40401), .C2(n33136), .ZN(n9252) );
  OAI222_X1 U31503 ( .A1(n40978), .A2(n40410), .B1(n41362), .B2(n40403), .C1(
        n40401), .C2(n33135), .ZN(n9251) );
  OAI222_X1 U31504 ( .A1(n40953), .A2(n40210), .B1(n41337), .B2(n40203), .C1(
        n40201), .C2(n33103), .ZN(n8615) );
  OAI222_X1 U31505 ( .A1(n40965), .A2(n40210), .B1(n41349), .B2(n40203), .C1(
        n40201), .C2(n33101), .ZN(n8613) );
  OAI222_X1 U31506 ( .A1(n40971), .A2(n40210), .B1(n41355), .B2(n40203), .C1(
        n40201), .C2(n33100), .ZN(n8612) );
  OAI222_X1 U31507 ( .A1(n40977), .A2(n40210), .B1(n41361), .B2(n40203), .C1(
        n40201), .C2(n33099), .ZN(n8611) );
  OAI222_X1 U31508 ( .A1(n40953), .A2(n40230), .B1(n41337), .B2(n40223), .C1(
        n40221), .C2(n33091), .ZN(n8679) );
  OAI222_X1 U31509 ( .A1(n40965), .A2(n40230), .B1(n41349), .B2(n40223), .C1(
        n40221), .C2(n33089), .ZN(n8677) );
  OAI222_X1 U31510 ( .A1(n40971), .A2(n40230), .B1(n41355), .B2(n40223), .C1(
        n40221), .C2(n33088), .ZN(n8676) );
  OAI222_X1 U31511 ( .A1(n40977), .A2(n40230), .B1(n41361), .B2(n40223), .C1(
        n40221), .C2(n33087), .ZN(n8675) );
  OAI222_X1 U31512 ( .A1(n40954), .A2(n40310), .B1(n41338), .B2(n40303), .C1(
        n40301), .C2(n32719), .ZN(n8935) );
  OAI222_X1 U31513 ( .A1(n40966), .A2(n40310), .B1(n41350), .B2(n40303), .C1(
        n40301), .C2(n32717), .ZN(n8933) );
  OAI222_X1 U31514 ( .A1(n40972), .A2(n40310), .B1(n41356), .B2(n40303), .C1(
        n40301), .C2(n32716), .ZN(n8932) );
  OAI222_X1 U31515 ( .A1(n40978), .A2(n40310), .B1(n41362), .B2(n40303), .C1(
        n40301), .C2(n32715), .ZN(n8931) );
  OAI222_X1 U31516 ( .A1(n40954), .A2(n40330), .B1(n41338), .B2(n40323), .C1(
        n40321), .C2(n32707), .ZN(n8999) );
  OAI222_X1 U31517 ( .A1(n40966), .A2(n40330), .B1(n41350), .B2(n40323), .C1(
        n40321), .C2(n32705), .ZN(n8997) );
  OAI222_X1 U31518 ( .A1(n40972), .A2(n40330), .B1(n41356), .B2(n40323), .C1(
        n40321), .C2(n32704), .ZN(n8996) );
  OAI222_X1 U31519 ( .A1(n40978), .A2(n40330), .B1(n41362), .B2(n40323), .C1(
        n40321), .C2(n32703), .ZN(n8995) );
  OAI222_X1 U31520 ( .A1(n40955), .A2(n40530), .B1(n41339), .B2(n40523), .C1(
        n40521), .C2(n32444), .ZN(n9639) );
  OAI222_X1 U31521 ( .A1(n40967), .A2(n40530), .B1(n41351), .B2(n40523), .C1(
        n40521), .C2(n38791), .ZN(n9637) );
  OAI222_X1 U31522 ( .A1(n40973), .A2(n40530), .B1(n41357), .B2(n40523), .C1(
        n40521), .C2(n38792), .ZN(n9636) );
  OAI222_X1 U31523 ( .A1(n40979), .A2(n40530), .B1(n41363), .B2(n40523), .C1(
        n40521), .C2(n38793), .ZN(n9635) );
  OAI222_X1 U31524 ( .A1(n40954), .A2(n40510), .B1(n41338), .B2(n40503), .C1(
        n40501), .C2(n32384), .ZN(n9575) );
  OAI222_X1 U31525 ( .A1(n40966), .A2(n40510), .B1(n41350), .B2(n40503), .C1(
        n40501), .C2(n38924), .ZN(n9573) );
  OAI222_X1 U31526 ( .A1(n40972), .A2(n40510), .B1(n41356), .B2(n40503), .C1(
        n40501), .C2(n38925), .ZN(n9572) );
  OAI222_X1 U31527 ( .A1(n40978), .A2(n40510), .B1(n41362), .B2(n40503), .C1(
        n40501), .C2(n38926), .ZN(n9571) );
  OAI222_X1 U31528 ( .A1(n40952), .A2(n39835), .B1(n41336), .B2(n39828), .C1(
        n39826), .C2(n32695), .ZN(n7399) );
  OAI222_X1 U31529 ( .A1(n40964), .A2(n39835), .B1(n41348), .B2(n39828), .C1(
        n39826), .C2(n32693), .ZN(n7397) );
  OAI222_X1 U31530 ( .A1(n40970), .A2(n39835), .B1(n41354), .B2(n39828), .C1(
        n39826), .C2(n32692), .ZN(n7396) );
  OAI222_X1 U31531 ( .A1(n40976), .A2(n39835), .B1(n41360), .B2(n39828), .C1(
        n39826), .C2(n32691), .ZN(n7395) );
  NOR3_X1 U31532 ( .A1(n33297), .A2(n23853), .A3(n32081), .ZN(n33332) );
  AOI221_X1 U31533 ( .B1(n39282), .B2(n30055), .C1(n39276), .C2(n30119), .A(
        n37016), .ZN(n37015) );
  OAI222_X1 U31534 ( .A1(n32043), .A2(n39270), .B1(n32067), .B2(n39264), .C1(
        n31983), .C2(n39258), .ZN(n37016) );
  AOI221_X1 U31535 ( .B1(n39283), .B2(n30054), .C1(n39277), .C2(n30118), .A(
        n36997), .ZN(n36996) );
  OAI222_X1 U31536 ( .A1(n32042), .A2(n39271), .B1(n32066), .B2(n39265), .C1(
        n31982), .C2(n39259), .ZN(n36997) );
  AOI221_X1 U31537 ( .B1(n39283), .B2(n30053), .C1(n39277), .C2(n30117), .A(
        n36978), .ZN(n36977) );
  OAI222_X1 U31538 ( .A1(n32041), .A2(n39271), .B1(n32065), .B2(n39265), .C1(
        n31981), .C2(n39259), .ZN(n36978) );
  AOI221_X1 U31539 ( .B1(n39283), .B2(n30052), .C1(n39277), .C2(n30116), .A(
        n36959), .ZN(n36958) );
  OAI222_X1 U31540 ( .A1(n32040), .A2(n39271), .B1(n32064), .B2(n39265), .C1(
        n31980), .C2(n39259), .ZN(n36959) );
  AOI221_X1 U31541 ( .B1(n39283), .B2(n30051), .C1(n39277), .C2(n30115), .A(
        n36940), .ZN(n36939) );
  OAI222_X1 U31542 ( .A1(n32039), .A2(n39271), .B1(n32063), .B2(n39265), .C1(
        n31979), .C2(n39259), .ZN(n36940) );
  AOI221_X1 U31543 ( .B1(n39283), .B2(n30050), .C1(n39277), .C2(n30114), .A(
        n36921), .ZN(n36920) );
  OAI222_X1 U31544 ( .A1(n32038), .A2(n39271), .B1(n32062), .B2(n39265), .C1(
        n31978), .C2(n39259), .ZN(n36921) );
  AOI221_X1 U31545 ( .B1(n39283), .B2(n30049), .C1(n39277), .C2(n30113), .A(
        n36902), .ZN(n36901) );
  OAI222_X1 U31546 ( .A1(n32037), .A2(n39271), .B1(n32061), .B2(n39265), .C1(
        n31977), .C2(n39259), .ZN(n36902) );
  AOI221_X1 U31547 ( .B1(n39283), .B2(n30048), .C1(n39277), .C2(n30112), .A(
        n36883), .ZN(n36882) );
  OAI222_X1 U31548 ( .A1(n32036), .A2(n39271), .B1(n32060), .B2(n39265), .C1(
        n31976), .C2(n39259), .ZN(n36883) );
  AOI221_X1 U31549 ( .B1(n39283), .B2(n30047), .C1(n39277), .C2(n30111), .A(
        n36864), .ZN(n36863) );
  OAI222_X1 U31550 ( .A1(n32035), .A2(n39271), .B1(n32059), .B2(n39265), .C1(
        n31975), .C2(n39259), .ZN(n36864) );
  AOI221_X1 U31551 ( .B1(n39283), .B2(n30046), .C1(n39277), .C2(n30110), .A(
        n36845), .ZN(n36844) );
  OAI222_X1 U31552 ( .A1(n32034), .A2(n39271), .B1(n32058), .B2(n39265), .C1(
        n31974), .C2(n39259), .ZN(n36845) );
  AOI221_X1 U31553 ( .B1(n39283), .B2(n30045), .C1(n39277), .C2(n30109), .A(
        n36826), .ZN(n36825) );
  OAI222_X1 U31554 ( .A1(n32033), .A2(n39271), .B1(n32057), .B2(n39265), .C1(
        n31973), .C2(n39259), .ZN(n36826) );
  AOI221_X1 U31555 ( .B1(n39283), .B2(n30044), .C1(n39277), .C2(n30108), .A(
        n36807), .ZN(n36806) );
  OAI222_X1 U31556 ( .A1(n32032), .A2(n39271), .B1(n32056), .B2(n39265), .C1(
        n31972), .C2(n39259), .ZN(n36807) );
  AOI221_X1 U31557 ( .B1(n39283), .B2(n30043), .C1(n39277), .C2(n30107), .A(
        n36788), .ZN(n36787) );
  OAI222_X1 U31558 ( .A1(n32031), .A2(n39271), .B1(n32055), .B2(n39265), .C1(
        n31971), .C2(n39259), .ZN(n36788) );
  AOI221_X1 U31559 ( .B1(n39284), .B2(n30042), .C1(n39278), .C2(n30106), .A(
        n36769), .ZN(n36768) );
  OAI222_X1 U31560 ( .A1(n32030), .A2(n39272), .B1(n32321), .B2(n39266), .C1(
        n31970), .C2(n39260), .ZN(n36769) );
  AOI221_X1 U31561 ( .B1(n39284), .B2(n30041), .C1(n39278), .C2(n30105), .A(
        n36750), .ZN(n36749) );
  OAI222_X1 U31562 ( .A1(n32029), .A2(n39272), .B1(n32320), .B2(n39266), .C1(
        n31969), .C2(n39260), .ZN(n36750) );
  AOI221_X1 U31563 ( .B1(n39284), .B2(n30040), .C1(n39278), .C2(n30104), .A(
        n36731), .ZN(n36730) );
  OAI222_X1 U31564 ( .A1(n32028), .A2(n39272), .B1(n32319), .B2(n39266), .C1(
        n31968), .C2(n39260), .ZN(n36731) );
  AOI221_X1 U31565 ( .B1(n39284), .B2(n30039), .C1(n39278), .C2(n30103), .A(
        n36712), .ZN(n36711) );
  OAI222_X1 U31566 ( .A1(n32027), .A2(n39272), .B1(n32318), .B2(n39266), .C1(
        n31967), .C2(n39260), .ZN(n36712) );
  AOI221_X1 U31567 ( .B1(n39284), .B2(n30038), .C1(n39278), .C2(n30102), .A(
        n36693), .ZN(n36692) );
  OAI222_X1 U31568 ( .A1(n32026), .A2(n39272), .B1(n32317), .B2(n39266), .C1(
        n31966), .C2(n39260), .ZN(n36693) );
  AOI221_X1 U31569 ( .B1(n39284), .B2(n30037), .C1(n39278), .C2(n30101), .A(
        n36674), .ZN(n36673) );
  OAI222_X1 U31570 ( .A1(n32025), .A2(n39272), .B1(n32316), .B2(n39266), .C1(
        n31965), .C2(n39260), .ZN(n36674) );
  AOI221_X1 U31571 ( .B1(n39284), .B2(n30036), .C1(n39278), .C2(n30100), .A(
        n36655), .ZN(n36654) );
  OAI222_X1 U31572 ( .A1(n32024), .A2(n39272), .B1(n32315), .B2(n39266), .C1(
        n31964), .C2(n39260), .ZN(n36655) );
  AOI221_X1 U31573 ( .B1(n39284), .B2(n30035), .C1(n39278), .C2(n30099), .A(
        n36636), .ZN(n36635) );
  OAI222_X1 U31574 ( .A1(n32023), .A2(n39272), .B1(n32314), .B2(n39266), .C1(
        n31963), .C2(n39260), .ZN(n36636) );
  AOI221_X1 U31575 ( .B1(n39284), .B2(n30034), .C1(n39278), .C2(n30098), .A(
        n36617), .ZN(n36616) );
  OAI222_X1 U31576 ( .A1(n32022), .A2(n39272), .B1(n32313), .B2(n39266), .C1(
        n31962), .C2(n39260), .ZN(n36617) );
  AOI221_X1 U31577 ( .B1(n39284), .B2(n30033), .C1(n39278), .C2(n30097), .A(
        n36598), .ZN(n36597) );
  OAI222_X1 U31578 ( .A1(n32021), .A2(n39272), .B1(n32312), .B2(n39266), .C1(
        n31961), .C2(n39260), .ZN(n36598) );
  AOI221_X1 U31579 ( .B1(n39284), .B2(n30032), .C1(n39278), .C2(n30096), .A(
        n36579), .ZN(n36578) );
  OAI222_X1 U31580 ( .A1(n32020), .A2(n39272), .B1(n32311), .B2(n39266), .C1(
        n31960), .C2(n39260), .ZN(n36579) );
  AOI221_X1 U31581 ( .B1(n39284), .B2(n30031), .C1(n39278), .C2(n30095), .A(
        n36560), .ZN(n36559) );
  OAI222_X1 U31582 ( .A1(n32019), .A2(n39272), .B1(n32310), .B2(n39266), .C1(
        n31959), .C2(n39260), .ZN(n36560) );
  AOI221_X1 U31583 ( .B1(n39285), .B2(n30030), .C1(n39279), .C2(n30094), .A(
        n36541), .ZN(n36540) );
  OAI222_X1 U31584 ( .A1(n32018), .A2(n39273), .B1(n32309), .B2(n39267), .C1(
        n31958), .C2(n39261), .ZN(n36541) );
  AOI221_X1 U31585 ( .B1(n39285), .B2(n30029), .C1(n39279), .C2(n30093), .A(
        n36522), .ZN(n36521) );
  OAI222_X1 U31586 ( .A1(n32017), .A2(n39273), .B1(n32308), .B2(n39267), .C1(
        n31957), .C2(n39261), .ZN(n36522) );
  AOI221_X1 U31587 ( .B1(n39285), .B2(n30028), .C1(n39279), .C2(n30092), .A(
        n36503), .ZN(n36502) );
  OAI222_X1 U31588 ( .A1(n32016), .A2(n39273), .B1(n32307), .B2(n39267), .C1(
        n31956), .C2(n39261), .ZN(n36503) );
  AOI221_X1 U31589 ( .B1(n39285), .B2(n30027), .C1(n39279), .C2(n30091), .A(
        n36484), .ZN(n36483) );
  OAI222_X1 U31590 ( .A1(n32015), .A2(n39273), .B1(n32306), .B2(n39267), .C1(
        n31955), .C2(n39261), .ZN(n36484) );
  AOI221_X1 U31591 ( .B1(n39285), .B2(n30026), .C1(n39279), .C2(n30090), .A(
        n36465), .ZN(n36464) );
  OAI222_X1 U31592 ( .A1(n32014), .A2(n39273), .B1(n32305), .B2(n39267), .C1(
        n31954), .C2(n39261), .ZN(n36465) );
  AOI221_X1 U31593 ( .B1(n39285), .B2(n30025), .C1(n39279), .C2(n30089), .A(
        n36446), .ZN(n36445) );
  OAI222_X1 U31594 ( .A1(n32013), .A2(n39273), .B1(n32304), .B2(n39267), .C1(
        n31953), .C2(n39261), .ZN(n36446) );
  AOI221_X1 U31595 ( .B1(n39285), .B2(n30024), .C1(n39279), .C2(n30088), .A(
        n36427), .ZN(n36426) );
  OAI222_X1 U31596 ( .A1(n32012), .A2(n39273), .B1(n32303), .B2(n39267), .C1(
        n31952), .C2(n39261), .ZN(n36427) );
  AOI221_X1 U31597 ( .B1(n39285), .B2(n30023), .C1(n39279), .C2(n30087), .A(
        n36408), .ZN(n36407) );
  OAI222_X1 U31598 ( .A1(n32011), .A2(n39273), .B1(n32302), .B2(n39267), .C1(
        n31951), .C2(n39261), .ZN(n36408) );
  AOI221_X1 U31599 ( .B1(n39285), .B2(n30022), .C1(n39279), .C2(n30086), .A(
        n36389), .ZN(n36388) );
  OAI222_X1 U31600 ( .A1(n32010), .A2(n39273), .B1(n32301), .B2(n39267), .C1(
        n31950), .C2(n39261), .ZN(n36389) );
  AOI221_X1 U31601 ( .B1(n39285), .B2(n30021), .C1(n39279), .C2(n30085), .A(
        n36370), .ZN(n36369) );
  OAI222_X1 U31602 ( .A1(n32009), .A2(n39273), .B1(n32300), .B2(n39267), .C1(
        n31949), .C2(n39261), .ZN(n36370) );
  AOI221_X1 U31603 ( .B1(n39285), .B2(n30020), .C1(n39279), .C2(n30084), .A(
        n36351), .ZN(n36350) );
  OAI222_X1 U31604 ( .A1(n32008), .A2(n39273), .B1(n32299), .B2(n39267), .C1(
        n31948), .C2(n39261), .ZN(n36351) );
  AOI221_X1 U31605 ( .B1(n39285), .B2(n30019), .C1(n39279), .C2(n30083), .A(
        n36332), .ZN(n36331) );
  OAI222_X1 U31606 ( .A1(n32007), .A2(n39273), .B1(n32298), .B2(n39267), .C1(
        n31947), .C2(n39261), .ZN(n36332) );
  AOI221_X1 U31607 ( .B1(n39286), .B2(n30018), .C1(n39280), .C2(n30082), .A(
        n36313), .ZN(n36312) );
  OAI222_X1 U31608 ( .A1(n32006), .A2(n39274), .B1(n32297), .B2(n39268), .C1(
        n31946), .C2(n39262), .ZN(n36313) );
  AOI221_X1 U31609 ( .B1(n39286), .B2(n30017), .C1(n39280), .C2(n30081), .A(
        n36294), .ZN(n36293) );
  OAI222_X1 U31610 ( .A1(n32005), .A2(n39274), .B1(n32296), .B2(n39268), .C1(
        n31945), .C2(n39262), .ZN(n36294) );
  AOI221_X1 U31611 ( .B1(n39286), .B2(n30016), .C1(n39280), .C2(n30080), .A(
        n36275), .ZN(n36274) );
  OAI222_X1 U31612 ( .A1(n32004), .A2(n39274), .B1(n32295), .B2(n39268), .C1(
        n31944), .C2(n39262), .ZN(n36275) );
  AOI221_X1 U31613 ( .B1(n39286), .B2(n30015), .C1(n39280), .C2(n30079), .A(
        n36256), .ZN(n36255) );
  OAI222_X1 U31614 ( .A1(n32003), .A2(n39274), .B1(n32294), .B2(n39268), .C1(
        n31943), .C2(n39262), .ZN(n36256) );
  AOI221_X1 U31615 ( .B1(n39286), .B2(n30014), .C1(n39280), .C2(n30078), .A(
        n36237), .ZN(n36236) );
  OAI222_X1 U31616 ( .A1(n32002), .A2(n39274), .B1(n32293), .B2(n39268), .C1(
        n31942), .C2(n39262), .ZN(n36237) );
  AOI221_X1 U31617 ( .B1(n39286), .B2(n30013), .C1(n39280), .C2(n30077), .A(
        n36218), .ZN(n36217) );
  OAI222_X1 U31618 ( .A1(n32001), .A2(n39274), .B1(n32292), .B2(n39268), .C1(
        n31941), .C2(n39262), .ZN(n36218) );
  AOI221_X1 U31619 ( .B1(n39162), .B2(n31119), .C1(n39156), .C2(n28849), .A(
        n37214), .ZN(n37213) );
  OAI222_X1 U31620 ( .A1(n31301), .A2(n39150), .B1(n31365), .B2(n39144), .C1(
        n31237), .C2(n39138), .ZN(n37214) );
  AOI221_X1 U31621 ( .B1(n39282), .B2(n30065), .C1(n39276), .C2(n30129), .A(
        n37206), .ZN(n37205) );
  OAI222_X1 U31622 ( .A1(n32280), .A2(n39270), .B1(n32264), .B2(n39264), .C1(
        n32284), .C2(n39258), .ZN(n37206) );
  AOI221_X1 U31623 ( .B1(n39162), .B2(n31118), .C1(n39156), .C2(n28848), .A(
        n37195), .ZN(n37194) );
  OAI222_X1 U31624 ( .A1(n31300), .A2(n39150), .B1(n31364), .B2(n39144), .C1(
        n31236), .C2(n39138), .ZN(n37195) );
  AOI221_X1 U31625 ( .B1(n39282), .B2(n30064), .C1(n39276), .C2(n30128), .A(
        n37187), .ZN(n37186) );
  OAI222_X1 U31626 ( .A1(n32279), .A2(n39270), .B1(n32263), .B2(n39264), .C1(
        n32283), .C2(n39258), .ZN(n37187) );
  AOI221_X1 U31627 ( .B1(n39162), .B2(n31117), .C1(n39156), .C2(n28847), .A(
        n37176), .ZN(n37175) );
  OAI222_X1 U31628 ( .A1(n31299), .A2(n39150), .B1(n31363), .B2(n39144), .C1(
        n31235), .C2(n39138), .ZN(n37176) );
  AOI221_X1 U31629 ( .B1(n39282), .B2(n30063), .C1(n39276), .C2(n30127), .A(
        n37168), .ZN(n37167) );
  OAI222_X1 U31630 ( .A1(n32278), .A2(n39270), .B1(n32262), .B2(n39264), .C1(
        n32282), .C2(n39258), .ZN(n37168) );
  AOI221_X1 U31631 ( .B1(n39162), .B2(n31116), .C1(n39156), .C2(n28846), .A(
        n37157), .ZN(n37156) );
  OAI222_X1 U31632 ( .A1(n31298), .A2(n39150), .B1(n31362), .B2(n39144), .C1(
        n31234), .C2(n39138), .ZN(n37157) );
  AOI221_X1 U31633 ( .B1(n39282), .B2(n30062), .C1(n39276), .C2(n30126), .A(
        n37149), .ZN(n37148) );
  OAI222_X1 U31634 ( .A1(n32050), .A2(n39270), .B1(n32074), .B2(n39264), .C1(
        n31990), .C2(n39258), .ZN(n37149) );
  AOI221_X1 U31635 ( .B1(n39162), .B2(n31115), .C1(n39156), .C2(n28845), .A(
        n37138), .ZN(n37137) );
  OAI222_X1 U31636 ( .A1(n31297), .A2(n39150), .B1(n31361), .B2(n39144), .C1(
        n31233), .C2(n39138), .ZN(n37138) );
  AOI221_X1 U31637 ( .B1(n39282), .B2(n30061), .C1(n39276), .C2(n30125), .A(
        n37130), .ZN(n37129) );
  OAI222_X1 U31638 ( .A1(n32049), .A2(n39270), .B1(n32073), .B2(n39264), .C1(
        n31989), .C2(n39258), .ZN(n37130) );
  AOI221_X1 U31639 ( .B1(n39162), .B2(n31120), .C1(n39156), .C2(n28850), .A(
        n37245), .ZN(n37244) );
  OAI222_X1 U31640 ( .A1(n31302), .A2(n39150), .B1(n31366), .B2(n39144), .C1(
        n31238), .C2(n39138), .ZN(n37245) );
  AOI221_X1 U31641 ( .B1(n39282), .B2(n30066), .C1(n39276), .C2(n30130), .A(
        n37225), .ZN(n37224) );
  OAI222_X1 U31642 ( .A1(n32281), .A2(n39270), .B1(n32265), .B2(n39264), .C1(
        n32285), .C2(n39258), .ZN(n37225) );
  AOI221_X1 U31643 ( .B1(n39162), .B2(n31114), .C1(n39156), .C2(n28844), .A(
        n37119), .ZN(n37118) );
  OAI222_X1 U31644 ( .A1(n31296), .A2(n39150), .B1(n31360), .B2(n39144), .C1(
        n31232), .C2(n39138), .ZN(n37119) );
  AOI221_X1 U31645 ( .B1(n39282), .B2(n30060), .C1(n39276), .C2(n30124), .A(
        n37111), .ZN(n37110) );
  OAI222_X1 U31646 ( .A1(n32048), .A2(n39270), .B1(n32072), .B2(n39264), .C1(
        n31988), .C2(n39258), .ZN(n37111) );
  AOI221_X1 U31647 ( .B1(n39162), .B2(n31113), .C1(n39156), .C2(n28843), .A(
        n37100), .ZN(n37099) );
  OAI222_X1 U31648 ( .A1(n31295), .A2(n39150), .B1(n31359), .B2(n39144), .C1(
        n31231), .C2(n39138), .ZN(n37100) );
  AOI221_X1 U31649 ( .B1(n39282), .B2(n30059), .C1(n39276), .C2(n30123), .A(
        n37092), .ZN(n37091) );
  OAI222_X1 U31650 ( .A1(n32047), .A2(n39270), .B1(n32071), .B2(n39264), .C1(
        n31987), .C2(n39258), .ZN(n37092) );
  AOI221_X1 U31651 ( .B1(n39162), .B2(n31112), .C1(n39156), .C2(n28842), .A(
        n37081), .ZN(n37080) );
  OAI222_X1 U31652 ( .A1(n31294), .A2(n39150), .B1(n31358), .B2(n39144), .C1(
        n31230), .C2(n39138), .ZN(n37081) );
  AOI221_X1 U31653 ( .B1(n39282), .B2(n30058), .C1(n39276), .C2(n30122), .A(
        n37073), .ZN(n37072) );
  OAI222_X1 U31654 ( .A1(n32046), .A2(n39270), .B1(n32070), .B2(n39264), .C1(
        n31986), .C2(n39258), .ZN(n37073) );
  AOI221_X1 U31655 ( .B1(n39162), .B2(n31111), .C1(n39156), .C2(n28841), .A(
        n37062), .ZN(n37061) );
  OAI222_X1 U31656 ( .A1(n31293), .A2(n39150), .B1(n31357), .B2(n39144), .C1(
        n31229), .C2(n39138), .ZN(n37062) );
  AOI221_X1 U31657 ( .B1(n39282), .B2(n30057), .C1(n39276), .C2(n30121), .A(
        n37054), .ZN(n37053) );
  OAI222_X1 U31658 ( .A1(n32045), .A2(n39270), .B1(n32069), .B2(n39264), .C1(
        n31985), .C2(n39258), .ZN(n37054) );
  AOI221_X1 U31659 ( .B1(n39282), .B2(n30056), .C1(n39276), .C2(n30120), .A(
        n37035), .ZN(n37034) );
  OAI222_X1 U31660 ( .A1(n32044), .A2(n39270), .B1(n32068), .B2(n39264), .C1(
        n31984), .C2(n39258), .ZN(n37035) );
  AOI221_X1 U31661 ( .B1(n39286), .B2(n30012), .C1(n39280), .C2(n30076), .A(
        n36199), .ZN(n36198) );
  OAI222_X1 U31662 ( .A1(n32000), .A2(n39274), .B1(n32291), .B2(n39268), .C1(
        n31940), .C2(n39262), .ZN(n36199) );
  AOI221_X1 U31663 ( .B1(n39286), .B2(n30011), .C1(n39280), .C2(n30075), .A(
        n36180), .ZN(n36179) );
  OAI222_X1 U31664 ( .A1(n31999), .A2(n39274), .B1(n32290), .B2(n39268), .C1(
        n31939), .C2(n39262), .ZN(n36180) );
  AOI221_X1 U31665 ( .B1(n39286), .B2(n30010), .C1(n39280), .C2(n30074), .A(
        n36161), .ZN(n36160) );
  OAI222_X1 U31666 ( .A1(n31998), .A2(n39274), .B1(n32289), .B2(n39268), .C1(
        n31938), .C2(n39262), .ZN(n36161) );
  AOI221_X1 U31667 ( .B1(n39286), .B2(n30009), .C1(n39280), .C2(n30073), .A(
        n36142), .ZN(n36141) );
  OAI222_X1 U31668 ( .A1(n31997), .A2(n39274), .B1(n32288), .B2(n39268), .C1(
        n31937), .C2(n39262), .ZN(n36142) );
  AOI221_X1 U31669 ( .B1(n39286), .B2(n30008), .C1(n39280), .C2(n30072), .A(
        n36123), .ZN(n36122) );
  OAI222_X1 U31670 ( .A1(n31996), .A2(n39274), .B1(n32287), .B2(n39268), .C1(
        n31936), .C2(n39262), .ZN(n36123) );
  AOI221_X1 U31671 ( .B1(n39286), .B2(n30007), .C1(n39280), .C2(n30071), .A(
        n36104), .ZN(n36103) );
  OAI222_X1 U31672 ( .A1(n31995), .A2(n39274), .B1(n32054), .B2(n39268), .C1(
        n31935), .C2(n39262), .ZN(n36104) );
  AOI221_X1 U31673 ( .B1(n39669), .B2(n31120), .C1(n39663), .C2(n28850), .A(
        n33463), .ZN(n33460) );
  OAI222_X1 U31674 ( .A1(n31302), .A2(n39657), .B1(n31366), .B2(n39651), .C1(
        n31238), .C2(n39645), .ZN(n33463) );
  AOI221_X1 U31675 ( .B1(n39789), .B2(n30066), .C1(n39783), .C2(n30130), .A(
        n33435), .ZN(n33432) );
  OAI222_X1 U31676 ( .A1(n32281), .A2(n39777), .B1(n32265), .B2(n39771), .C1(
        n32285), .C2(n39765), .ZN(n33435) );
  AOI221_X1 U31677 ( .B1(n39417), .B2(n31120), .C1(n39411), .C2(n28850), .A(
        n34737), .ZN(n34734) );
  OAI222_X1 U31678 ( .A1(n31302), .A2(n39405), .B1(n31366), .B2(n39399), .C1(
        n31238), .C2(n39393), .ZN(n34737) );
  AOI221_X1 U31679 ( .B1(n39537), .B2(n30066), .C1(n39531), .C2(n30130), .A(
        n34709), .ZN(n34706) );
  OAI222_X1 U31680 ( .A1(n32281), .A2(n39525), .B1(n32265), .B2(n39519), .C1(
        n32285), .C2(n39513), .ZN(n34709) );
  AOI221_X1 U31681 ( .B1(n39669), .B2(n31119), .C1(n39663), .C2(n28849), .A(
        n33500), .ZN(n33499) );
  OAI222_X1 U31682 ( .A1(n31301), .A2(n39657), .B1(n31365), .B2(n39651), .C1(
        n31237), .C2(n39645), .ZN(n33500) );
  AOI221_X1 U31683 ( .B1(n39789), .B2(n30065), .C1(n39783), .C2(n30129), .A(
        n33492), .ZN(n33491) );
  OAI222_X1 U31684 ( .A1(n32280), .A2(n39777), .B1(n32264), .B2(n39771), .C1(
        n32284), .C2(n39765), .ZN(n33492) );
  AOI221_X1 U31685 ( .B1(n39417), .B2(n31119), .C1(n39411), .C2(n28849), .A(
        n34774), .ZN(n34773) );
  OAI222_X1 U31686 ( .A1(n31301), .A2(n39405), .B1(n31365), .B2(n39399), .C1(
        n31237), .C2(n39393), .ZN(n34774) );
  AOI221_X1 U31687 ( .B1(n39537), .B2(n30065), .C1(n39531), .C2(n30129), .A(
        n34766), .ZN(n34765) );
  OAI222_X1 U31688 ( .A1(n32280), .A2(n39525), .B1(n32264), .B2(n39519), .C1(
        n32284), .C2(n39513), .ZN(n34766) );
  AOI221_X1 U31689 ( .B1(n39669), .B2(n31118), .C1(n39663), .C2(n28848), .A(
        n33519), .ZN(n33518) );
  OAI222_X1 U31690 ( .A1(n31300), .A2(n39657), .B1(n31364), .B2(n39651), .C1(
        n31236), .C2(n39645), .ZN(n33519) );
  AOI221_X1 U31691 ( .B1(n39789), .B2(n30064), .C1(n39783), .C2(n30128), .A(
        n33511), .ZN(n33510) );
  OAI222_X1 U31692 ( .A1(n32279), .A2(n39777), .B1(n32263), .B2(n39771), .C1(
        n32283), .C2(n39765), .ZN(n33511) );
  AOI221_X1 U31693 ( .B1(n39417), .B2(n31118), .C1(n39411), .C2(n28848), .A(
        n34793), .ZN(n34792) );
  OAI222_X1 U31694 ( .A1(n31300), .A2(n39405), .B1(n31364), .B2(n39399), .C1(
        n31236), .C2(n39393), .ZN(n34793) );
  AOI221_X1 U31695 ( .B1(n39537), .B2(n30064), .C1(n39531), .C2(n30128), .A(
        n34785), .ZN(n34784) );
  OAI222_X1 U31696 ( .A1(n32279), .A2(n39525), .B1(n32263), .B2(n39519), .C1(
        n32283), .C2(n39513), .ZN(n34785) );
  AOI221_X1 U31697 ( .B1(n39669), .B2(n31117), .C1(n39663), .C2(n28847), .A(
        n33538), .ZN(n33537) );
  OAI222_X1 U31698 ( .A1(n31299), .A2(n39657), .B1(n31363), .B2(n39651), .C1(
        n31235), .C2(n39645), .ZN(n33538) );
  AOI221_X1 U31699 ( .B1(n39789), .B2(n30063), .C1(n39783), .C2(n30127), .A(
        n33530), .ZN(n33529) );
  OAI222_X1 U31700 ( .A1(n32278), .A2(n39777), .B1(n32262), .B2(n39771), .C1(
        n32282), .C2(n39765), .ZN(n33530) );
  AOI221_X1 U31701 ( .B1(n39417), .B2(n31117), .C1(n39411), .C2(n28847), .A(
        n34812), .ZN(n34811) );
  OAI222_X1 U31702 ( .A1(n31299), .A2(n39405), .B1(n31363), .B2(n39399), .C1(
        n31235), .C2(n39393), .ZN(n34812) );
  AOI221_X1 U31703 ( .B1(n39537), .B2(n30063), .C1(n39531), .C2(n30127), .A(
        n34804), .ZN(n34803) );
  OAI222_X1 U31704 ( .A1(n32278), .A2(n39525), .B1(n32262), .B2(n39519), .C1(
        n32282), .C2(n39513), .ZN(n34804) );
  AOI221_X1 U31705 ( .B1(n39668), .B2(n31116), .C1(n39662), .C2(n28846), .A(
        n33557), .ZN(n33556) );
  OAI222_X1 U31706 ( .A1(n31298), .A2(n39656), .B1(n31362), .B2(n39650), .C1(
        n31234), .C2(n39644), .ZN(n33557) );
  AOI221_X1 U31707 ( .B1(n39788), .B2(n30062), .C1(n39782), .C2(n30126), .A(
        n33549), .ZN(n33548) );
  OAI222_X1 U31708 ( .A1(n32050), .A2(n39776), .B1(n32074), .B2(n39770), .C1(
        n31990), .C2(n39764), .ZN(n33549) );
  AOI221_X1 U31709 ( .B1(n39416), .B2(n31116), .C1(n39410), .C2(n28846), .A(
        n34831), .ZN(n34830) );
  OAI222_X1 U31710 ( .A1(n31298), .A2(n39404), .B1(n31362), .B2(n39398), .C1(
        n31234), .C2(n39392), .ZN(n34831) );
  AOI221_X1 U31711 ( .B1(n39536), .B2(n30062), .C1(n39530), .C2(n30126), .A(
        n34823), .ZN(n34822) );
  OAI222_X1 U31712 ( .A1(n32050), .A2(n39524), .B1(n32074), .B2(n39518), .C1(
        n31990), .C2(n39512), .ZN(n34823) );
  AOI221_X1 U31713 ( .B1(n39668), .B2(n31115), .C1(n39662), .C2(n28845), .A(
        n33576), .ZN(n33575) );
  OAI222_X1 U31714 ( .A1(n31297), .A2(n39656), .B1(n31361), .B2(n39650), .C1(
        n31233), .C2(n39644), .ZN(n33576) );
  AOI221_X1 U31715 ( .B1(n39788), .B2(n30061), .C1(n39782), .C2(n30125), .A(
        n33568), .ZN(n33567) );
  OAI222_X1 U31716 ( .A1(n32049), .A2(n39776), .B1(n32073), .B2(n39770), .C1(
        n31989), .C2(n39764), .ZN(n33568) );
  AOI221_X1 U31717 ( .B1(n39416), .B2(n31115), .C1(n39410), .C2(n28845), .A(
        n34850), .ZN(n34849) );
  OAI222_X1 U31718 ( .A1(n31297), .A2(n39404), .B1(n31361), .B2(n39398), .C1(
        n31233), .C2(n39392), .ZN(n34850) );
  AOI221_X1 U31719 ( .B1(n39536), .B2(n30061), .C1(n39530), .C2(n30125), .A(
        n34842), .ZN(n34841) );
  OAI222_X1 U31720 ( .A1(n32049), .A2(n39524), .B1(n32073), .B2(n39518), .C1(
        n31989), .C2(n39512), .ZN(n34842) );
  AOI221_X1 U31721 ( .B1(n39668), .B2(n31114), .C1(n39662), .C2(n28844), .A(
        n33595), .ZN(n33594) );
  OAI222_X1 U31722 ( .A1(n31296), .A2(n39656), .B1(n31360), .B2(n39650), .C1(
        n31232), .C2(n39644), .ZN(n33595) );
  AOI221_X1 U31723 ( .B1(n39788), .B2(n30060), .C1(n39782), .C2(n30124), .A(
        n33587), .ZN(n33586) );
  OAI222_X1 U31724 ( .A1(n32048), .A2(n39776), .B1(n32072), .B2(n39770), .C1(
        n31988), .C2(n39764), .ZN(n33587) );
  AOI221_X1 U31725 ( .B1(n39416), .B2(n31114), .C1(n39410), .C2(n28844), .A(
        n34869), .ZN(n34868) );
  OAI222_X1 U31726 ( .A1(n31296), .A2(n39404), .B1(n31360), .B2(n39398), .C1(
        n31232), .C2(n39392), .ZN(n34869) );
  AOI221_X1 U31727 ( .B1(n39536), .B2(n30060), .C1(n39530), .C2(n30124), .A(
        n34861), .ZN(n34860) );
  OAI222_X1 U31728 ( .A1(n32048), .A2(n39524), .B1(n32072), .B2(n39518), .C1(
        n31988), .C2(n39512), .ZN(n34861) );
  AOI221_X1 U31729 ( .B1(n39668), .B2(n31113), .C1(n39662), .C2(n28843), .A(
        n33614), .ZN(n33613) );
  OAI222_X1 U31730 ( .A1(n31295), .A2(n39656), .B1(n31359), .B2(n39650), .C1(
        n31231), .C2(n39644), .ZN(n33614) );
  AOI221_X1 U31731 ( .B1(n39788), .B2(n30059), .C1(n39782), .C2(n30123), .A(
        n33606), .ZN(n33605) );
  OAI222_X1 U31732 ( .A1(n32047), .A2(n39776), .B1(n32071), .B2(n39770), .C1(
        n31987), .C2(n39764), .ZN(n33606) );
  AOI221_X1 U31733 ( .B1(n39416), .B2(n31113), .C1(n39410), .C2(n28843), .A(
        n34888), .ZN(n34887) );
  OAI222_X1 U31734 ( .A1(n31295), .A2(n39404), .B1(n31359), .B2(n39398), .C1(
        n31231), .C2(n39392), .ZN(n34888) );
  AOI221_X1 U31735 ( .B1(n39536), .B2(n30059), .C1(n39530), .C2(n30123), .A(
        n34880), .ZN(n34879) );
  OAI222_X1 U31736 ( .A1(n32047), .A2(n39524), .B1(n32071), .B2(n39518), .C1(
        n31987), .C2(n39512), .ZN(n34880) );
  AOI221_X1 U31737 ( .B1(n39668), .B2(n31112), .C1(n39662), .C2(n28842), .A(
        n33633), .ZN(n33632) );
  OAI222_X1 U31738 ( .A1(n31294), .A2(n39656), .B1(n31358), .B2(n39650), .C1(
        n31230), .C2(n39644), .ZN(n33633) );
  AOI221_X1 U31739 ( .B1(n39788), .B2(n30058), .C1(n39782), .C2(n30122), .A(
        n33625), .ZN(n33624) );
  OAI222_X1 U31740 ( .A1(n32046), .A2(n39776), .B1(n32070), .B2(n39770), .C1(
        n31986), .C2(n39764), .ZN(n33625) );
  AOI221_X1 U31741 ( .B1(n39416), .B2(n31112), .C1(n39410), .C2(n28842), .A(
        n34907), .ZN(n34906) );
  OAI222_X1 U31742 ( .A1(n31294), .A2(n39404), .B1(n31358), .B2(n39398), .C1(
        n31230), .C2(n39392), .ZN(n34907) );
  AOI221_X1 U31743 ( .B1(n39536), .B2(n30058), .C1(n39530), .C2(n30122), .A(
        n34899), .ZN(n34898) );
  OAI222_X1 U31744 ( .A1(n32046), .A2(n39524), .B1(n32070), .B2(n39518), .C1(
        n31986), .C2(n39512), .ZN(n34899) );
  AOI221_X1 U31745 ( .B1(n39668), .B2(n31111), .C1(n39662), .C2(n28841), .A(
        n33652), .ZN(n33651) );
  OAI222_X1 U31746 ( .A1(n31293), .A2(n39656), .B1(n31357), .B2(n39650), .C1(
        n31229), .C2(n39644), .ZN(n33652) );
  AOI221_X1 U31747 ( .B1(n39788), .B2(n30057), .C1(n39782), .C2(n30121), .A(
        n33644), .ZN(n33643) );
  OAI222_X1 U31748 ( .A1(n32045), .A2(n39776), .B1(n32069), .B2(n39770), .C1(
        n31985), .C2(n39764), .ZN(n33644) );
  AOI221_X1 U31749 ( .B1(n39416), .B2(n31111), .C1(n39410), .C2(n28841), .A(
        n34926), .ZN(n34925) );
  OAI222_X1 U31750 ( .A1(n31293), .A2(n39404), .B1(n31357), .B2(n39398), .C1(
        n31229), .C2(n39392), .ZN(n34926) );
  AOI221_X1 U31751 ( .B1(n39536), .B2(n30057), .C1(n39530), .C2(n30121), .A(
        n34918), .ZN(n34917) );
  OAI222_X1 U31752 ( .A1(n32045), .A2(n39524), .B1(n32069), .B2(n39518), .C1(
        n31985), .C2(n39512), .ZN(n34918) );
  AOI221_X1 U31753 ( .B1(n39788), .B2(n30056), .C1(n39782), .C2(n30120), .A(
        n33663), .ZN(n33662) );
  OAI222_X1 U31754 ( .A1(n32044), .A2(n39776), .B1(n32068), .B2(n39770), .C1(
        n31984), .C2(n39764), .ZN(n33663) );
  AOI221_X1 U31755 ( .B1(n39536), .B2(n30056), .C1(n39530), .C2(n30120), .A(
        n34937), .ZN(n34936) );
  OAI222_X1 U31756 ( .A1(n32044), .A2(n39524), .B1(n32068), .B2(n39518), .C1(
        n31984), .C2(n39512), .ZN(n34937) );
  AOI221_X1 U31757 ( .B1(n39788), .B2(n30055), .C1(n39782), .C2(n30119), .A(
        n33682), .ZN(n33681) );
  OAI222_X1 U31758 ( .A1(n32043), .A2(n39776), .B1(n32067), .B2(n39770), .C1(
        n31983), .C2(n39764), .ZN(n33682) );
  AOI221_X1 U31759 ( .B1(n39536), .B2(n30055), .C1(n39530), .C2(n30119), .A(
        n34956), .ZN(n34955) );
  OAI222_X1 U31760 ( .A1(n32043), .A2(n39524), .B1(n32067), .B2(n39518), .C1(
        n31983), .C2(n39512), .ZN(n34956) );
  AOI221_X1 U31761 ( .B1(n39788), .B2(n30054), .C1(n39782), .C2(n30118), .A(
        n33701), .ZN(n33700) );
  OAI222_X1 U31762 ( .A1(n32042), .A2(n39776), .B1(n32066), .B2(n39770), .C1(
        n31982), .C2(n39764), .ZN(n33701) );
  AOI221_X1 U31763 ( .B1(n39536), .B2(n30054), .C1(n39530), .C2(n30118), .A(
        n34975), .ZN(n34974) );
  OAI222_X1 U31764 ( .A1(n32042), .A2(n39524), .B1(n32066), .B2(n39518), .C1(
        n31982), .C2(n39512), .ZN(n34975) );
  AOI221_X1 U31765 ( .B1(n39788), .B2(n30053), .C1(n39782), .C2(n30117), .A(
        n33720), .ZN(n33719) );
  OAI222_X1 U31766 ( .A1(n32041), .A2(n39776), .B1(n32065), .B2(n39770), .C1(
        n31981), .C2(n39764), .ZN(n33720) );
  AOI221_X1 U31767 ( .B1(n39536), .B2(n30053), .C1(n39530), .C2(n30117), .A(
        n34994), .ZN(n34993) );
  OAI222_X1 U31768 ( .A1(n32041), .A2(n39524), .B1(n32065), .B2(n39518), .C1(
        n31981), .C2(n39512), .ZN(n34994) );
  AOI221_X1 U31769 ( .B1(n39788), .B2(n30052), .C1(n39782), .C2(n30116), .A(
        n33739), .ZN(n33738) );
  OAI222_X1 U31770 ( .A1(n32040), .A2(n39776), .B1(n32064), .B2(n39770), .C1(
        n31980), .C2(n39764), .ZN(n33739) );
  AOI221_X1 U31771 ( .B1(n39536), .B2(n30052), .C1(n39530), .C2(n30116), .A(
        n35013), .ZN(n35012) );
  OAI222_X1 U31772 ( .A1(n32040), .A2(n39524), .B1(n32064), .B2(n39518), .C1(
        n31980), .C2(n39512), .ZN(n35013) );
  AOI221_X1 U31773 ( .B1(n39788), .B2(n30051), .C1(n39782), .C2(n30115), .A(
        n33758), .ZN(n33757) );
  OAI222_X1 U31774 ( .A1(n32039), .A2(n39776), .B1(n32063), .B2(n39770), .C1(
        n31979), .C2(n39764), .ZN(n33758) );
  AOI221_X1 U31775 ( .B1(n39536), .B2(n30051), .C1(n39530), .C2(n30115), .A(
        n35032), .ZN(n35031) );
  OAI222_X1 U31776 ( .A1(n32039), .A2(n39524), .B1(n32063), .B2(n39518), .C1(
        n31979), .C2(n39512), .ZN(n35032) );
  AOI221_X1 U31777 ( .B1(n39787), .B2(n30050), .C1(n39781), .C2(n30114), .A(
        n33777), .ZN(n33776) );
  OAI222_X1 U31778 ( .A1(n32038), .A2(n39775), .B1(n32062), .B2(n39769), .C1(
        n31978), .C2(n39763), .ZN(n33777) );
  AOI221_X1 U31779 ( .B1(n39535), .B2(n30050), .C1(n39529), .C2(n30114), .A(
        n35051), .ZN(n35050) );
  OAI222_X1 U31780 ( .A1(n32038), .A2(n39523), .B1(n32062), .B2(n39517), .C1(
        n31978), .C2(n39511), .ZN(n35051) );
  AOI221_X1 U31781 ( .B1(n39787), .B2(n30049), .C1(n39781), .C2(n30113), .A(
        n33796), .ZN(n33795) );
  OAI222_X1 U31782 ( .A1(n32037), .A2(n39775), .B1(n32061), .B2(n39769), .C1(
        n31977), .C2(n39763), .ZN(n33796) );
  AOI221_X1 U31783 ( .B1(n39535), .B2(n30049), .C1(n39529), .C2(n30113), .A(
        n35070), .ZN(n35069) );
  OAI222_X1 U31784 ( .A1(n32037), .A2(n39523), .B1(n32061), .B2(n39517), .C1(
        n31977), .C2(n39511), .ZN(n35070) );
  AOI221_X1 U31785 ( .B1(n39787), .B2(n30048), .C1(n39781), .C2(n30112), .A(
        n33815), .ZN(n33814) );
  OAI222_X1 U31786 ( .A1(n32036), .A2(n39775), .B1(n32060), .B2(n39769), .C1(
        n31976), .C2(n39763), .ZN(n33815) );
  AOI221_X1 U31787 ( .B1(n39535), .B2(n30048), .C1(n39529), .C2(n30112), .A(
        n35089), .ZN(n35088) );
  OAI222_X1 U31788 ( .A1(n32036), .A2(n39523), .B1(n32060), .B2(n39517), .C1(
        n31976), .C2(n39511), .ZN(n35089) );
  AOI221_X1 U31789 ( .B1(n39787), .B2(n30047), .C1(n39781), .C2(n30111), .A(
        n33834), .ZN(n33833) );
  OAI222_X1 U31790 ( .A1(n32035), .A2(n39775), .B1(n32059), .B2(n39769), .C1(
        n31975), .C2(n39763), .ZN(n33834) );
  AOI221_X1 U31791 ( .B1(n39535), .B2(n30047), .C1(n39529), .C2(n30111), .A(
        n35108), .ZN(n35107) );
  OAI222_X1 U31792 ( .A1(n32035), .A2(n39523), .B1(n32059), .B2(n39517), .C1(
        n31975), .C2(n39511), .ZN(n35108) );
  AOI221_X1 U31793 ( .B1(n39787), .B2(n30046), .C1(n39781), .C2(n30110), .A(
        n33853), .ZN(n33852) );
  OAI222_X1 U31794 ( .A1(n32034), .A2(n39775), .B1(n32058), .B2(n39769), .C1(
        n31974), .C2(n39763), .ZN(n33853) );
  AOI221_X1 U31795 ( .B1(n39535), .B2(n30046), .C1(n39529), .C2(n30110), .A(
        n35127), .ZN(n35126) );
  OAI222_X1 U31796 ( .A1(n32034), .A2(n39523), .B1(n32058), .B2(n39517), .C1(
        n31974), .C2(n39511), .ZN(n35127) );
  AOI221_X1 U31797 ( .B1(n39787), .B2(n30045), .C1(n39781), .C2(n30109), .A(
        n33872), .ZN(n33871) );
  OAI222_X1 U31798 ( .A1(n32033), .A2(n39775), .B1(n32057), .B2(n39769), .C1(
        n31973), .C2(n39763), .ZN(n33872) );
  AOI221_X1 U31799 ( .B1(n39535), .B2(n30045), .C1(n39529), .C2(n30109), .A(
        n35146), .ZN(n35145) );
  OAI222_X1 U31800 ( .A1(n32033), .A2(n39523), .B1(n32057), .B2(n39517), .C1(
        n31973), .C2(n39511), .ZN(n35146) );
  AOI221_X1 U31801 ( .B1(n39787), .B2(n30044), .C1(n39781), .C2(n30108), .A(
        n33891), .ZN(n33890) );
  OAI222_X1 U31802 ( .A1(n32032), .A2(n39775), .B1(n32056), .B2(n39769), .C1(
        n31972), .C2(n39763), .ZN(n33891) );
  AOI221_X1 U31803 ( .B1(n39535), .B2(n30044), .C1(n39529), .C2(n30108), .A(
        n35165), .ZN(n35164) );
  OAI222_X1 U31804 ( .A1(n32032), .A2(n39523), .B1(n32056), .B2(n39517), .C1(
        n31972), .C2(n39511), .ZN(n35165) );
  AOI221_X1 U31805 ( .B1(n39787), .B2(n30043), .C1(n39781), .C2(n30107), .A(
        n33910), .ZN(n33909) );
  OAI222_X1 U31806 ( .A1(n32031), .A2(n39775), .B1(n32055), .B2(n39769), .C1(
        n31971), .C2(n39763), .ZN(n33910) );
  AOI221_X1 U31807 ( .B1(n39535), .B2(n30043), .C1(n39529), .C2(n30107), .A(
        n35184), .ZN(n35183) );
  OAI222_X1 U31808 ( .A1(n32031), .A2(n39523), .B1(n32055), .B2(n39517), .C1(
        n31971), .C2(n39511), .ZN(n35184) );
  AOI221_X1 U31809 ( .B1(n39787), .B2(n30042), .C1(n39781), .C2(n30106), .A(
        n33929), .ZN(n33928) );
  OAI222_X1 U31810 ( .A1(n32030), .A2(n39775), .B1(n32321), .B2(n39769), .C1(
        n31970), .C2(n39763), .ZN(n33929) );
  AOI221_X1 U31811 ( .B1(n39535), .B2(n30042), .C1(n39529), .C2(n30106), .A(
        n35203), .ZN(n35202) );
  OAI222_X1 U31812 ( .A1(n32030), .A2(n39523), .B1(n32321), .B2(n39517), .C1(
        n31970), .C2(n39511), .ZN(n35203) );
  AOI221_X1 U31813 ( .B1(n39787), .B2(n30041), .C1(n39781), .C2(n30105), .A(
        n33948), .ZN(n33947) );
  OAI222_X1 U31814 ( .A1(n32029), .A2(n39775), .B1(n32320), .B2(n39769), .C1(
        n31969), .C2(n39763), .ZN(n33948) );
  AOI221_X1 U31815 ( .B1(n39535), .B2(n30041), .C1(n39529), .C2(n30105), .A(
        n35222), .ZN(n35221) );
  OAI222_X1 U31816 ( .A1(n32029), .A2(n39523), .B1(n32320), .B2(n39517), .C1(
        n31969), .C2(n39511), .ZN(n35222) );
  AOI221_X1 U31817 ( .B1(n39787), .B2(n30040), .C1(n39781), .C2(n30104), .A(
        n33967), .ZN(n33966) );
  OAI222_X1 U31818 ( .A1(n32028), .A2(n39775), .B1(n32319), .B2(n39769), .C1(
        n31968), .C2(n39763), .ZN(n33967) );
  AOI221_X1 U31819 ( .B1(n39535), .B2(n30040), .C1(n39529), .C2(n30104), .A(
        n35241), .ZN(n35240) );
  OAI222_X1 U31820 ( .A1(n32028), .A2(n39523), .B1(n32319), .B2(n39517), .C1(
        n31968), .C2(n39511), .ZN(n35241) );
  AOI221_X1 U31821 ( .B1(n39787), .B2(n30039), .C1(n39781), .C2(n30103), .A(
        n33986), .ZN(n33985) );
  OAI222_X1 U31822 ( .A1(n32027), .A2(n39775), .B1(n32318), .B2(n39769), .C1(
        n31967), .C2(n39763), .ZN(n33986) );
  AOI221_X1 U31823 ( .B1(n39535), .B2(n30039), .C1(n39529), .C2(n30103), .A(
        n35260), .ZN(n35259) );
  OAI222_X1 U31824 ( .A1(n32027), .A2(n39523), .B1(n32318), .B2(n39517), .C1(
        n31967), .C2(n39511), .ZN(n35260) );
  AOI221_X1 U31825 ( .B1(n39786), .B2(n30038), .C1(n39780), .C2(n30102), .A(
        n34005), .ZN(n34004) );
  OAI222_X1 U31826 ( .A1(n32026), .A2(n39774), .B1(n32317), .B2(n39768), .C1(
        n31966), .C2(n39762), .ZN(n34005) );
  AOI221_X1 U31827 ( .B1(n39534), .B2(n30038), .C1(n39528), .C2(n30102), .A(
        n35279), .ZN(n35278) );
  OAI222_X1 U31828 ( .A1(n32026), .A2(n39522), .B1(n32317), .B2(n39516), .C1(
        n31966), .C2(n39510), .ZN(n35279) );
  AOI221_X1 U31829 ( .B1(n39786), .B2(n30037), .C1(n39780), .C2(n30101), .A(
        n34024), .ZN(n34023) );
  OAI222_X1 U31830 ( .A1(n32025), .A2(n39774), .B1(n32316), .B2(n39768), .C1(
        n31965), .C2(n39762), .ZN(n34024) );
  AOI221_X1 U31831 ( .B1(n39534), .B2(n30037), .C1(n39528), .C2(n30101), .A(
        n35298), .ZN(n35297) );
  OAI222_X1 U31832 ( .A1(n32025), .A2(n39522), .B1(n32316), .B2(n39516), .C1(
        n31965), .C2(n39510), .ZN(n35298) );
  AOI221_X1 U31833 ( .B1(n39786), .B2(n30036), .C1(n39780), .C2(n30100), .A(
        n34043), .ZN(n34042) );
  OAI222_X1 U31834 ( .A1(n32024), .A2(n39774), .B1(n32315), .B2(n39768), .C1(
        n31964), .C2(n39762), .ZN(n34043) );
  AOI221_X1 U31835 ( .B1(n39534), .B2(n30036), .C1(n39528), .C2(n30100), .A(
        n35317), .ZN(n35316) );
  OAI222_X1 U31836 ( .A1(n32024), .A2(n39522), .B1(n32315), .B2(n39516), .C1(
        n31964), .C2(n39510), .ZN(n35317) );
  AOI221_X1 U31837 ( .B1(n39786), .B2(n30035), .C1(n39780), .C2(n30099), .A(
        n34062), .ZN(n34061) );
  OAI222_X1 U31838 ( .A1(n32023), .A2(n39774), .B1(n32314), .B2(n39768), .C1(
        n31963), .C2(n39762), .ZN(n34062) );
  AOI221_X1 U31839 ( .B1(n39534), .B2(n30035), .C1(n39528), .C2(n30099), .A(
        n35336), .ZN(n35335) );
  OAI222_X1 U31840 ( .A1(n32023), .A2(n39522), .B1(n32314), .B2(n39516), .C1(
        n31963), .C2(n39510), .ZN(n35336) );
  AOI221_X1 U31841 ( .B1(n39786), .B2(n30034), .C1(n39780), .C2(n30098), .A(
        n34081), .ZN(n34080) );
  OAI222_X1 U31842 ( .A1(n32022), .A2(n39774), .B1(n32313), .B2(n39768), .C1(
        n31962), .C2(n39762), .ZN(n34081) );
  AOI221_X1 U31843 ( .B1(n39534), .B2(n30034), .C1(n39528), .C2(n30098), .A(
        n35355), .ZN(n35354) );
  OAI222_X1 U31844 ( .A1(n32022), .A2(n39522), .B1(n32313), .B2(n39516), .C1(
        n31962), .C2(n39510), .ZN(n35355) );
  AOI221_X1 U31845 ( .B1(n39786), .B2(n30033), .C1(n39780), .C2(n30097), .A(
        n34100), .ZN(n34099) );
  OAI222_X1 U31846 ( .A1(n32021), .A2(n39774), .B1(n32312), .B2(n39768), .C1(
        n31961), .C2(n39762), .ZN(n34100) );
  AOI221_X1 U31847 ( .B1(n39534), .B2(n30033), .C1(n39528), .C2(n30097), .A(
        n35374), .ZN(n35373) );
  OAI222_X1 U31848 ( .A1(n32021), .A2(n39522), .B1(n32312), .B2(n39516), .C1(
        n31961), .C2(n39510), .ZN(n35374) );
  AOI221_X1 U31849 ( .B1(n39786), .B2(n30032), .C1(n39780), .C2(n30096), .A(
        n34119), .ZN(n34118) );
  OAI222_X1 U31850 ( .A1(n32020), .A2(n39774), .B1(n32311), .B2(n39768), .C1(
        n31960), .C2(n39762), .ZN(n34119) );
  AOI221_X1 U31851 ( .B1(n39534), .B2(n30032), .C1(n39528), .C2(n30096), .A(
        n35393), .ZN(n35392) );
  OAI222_X1 U31852 ( .A1(n32020), .A2(n39522), .B1(n32311), .B2(n39516), .C1(
        n31960), .C2(n39510), .ZN(n35393) );
  AOI221_X1 U31853 ( .B1(n39786), .B2(n30031), .C1(n39780), .C2(n30095), .A(
        n34138), .ZN(n34137) );
  OAI222_X1 U31854 ( .A1(n32019), .A2(n39774), .B1(n32310), .B2(n39768), .C1(
        n31959), .C2(n39762), .ZN(n34138) );
  AOI221_X1 U31855 ( .B1(n39534), .B2(n30031), .C1(n39528), .C2(n30095), .A(
        n35412), .ZN(n35411) );
  OAI222_X1 U31856 ( .A1(n32019), .A2(n39522), .B1(n32310), .B2(n39516), .C1(
        n31959), .C2(n39510), .ZN(n35412) );
  AOI221_X1 U31857 ( .B1(n39786), .B2(n30030), .C1(n39780), .C2(n30094), .A(
        n34157), .ZN(n34156) );
  OAI222_X1 U31858 ( .A1(n32018), .A2(n39774), .B1(n32309), .B2(n39768), .C1(
        n31958), .C2(n39762), .ZN(n34157) );
  AOI221_X1 U31859 ( .B1(n39534), .B2(n30030), .C1(n39528), .C2(n30094), .A(
        n35431), .ZN(n35430) );
  OAI222_X1 U31860 ( .A1(n32018), .A2(n39522), .B1(n32309), .B2(n39516), .C1(
        n31958), .C2(n39510), .ZN(n35431) );
  AOI221_X1 U31861 ( .B1(n39786), .B2(n30029), .C1(n39780), .C2(n30093), .A(
        n34176), .ZN(n34175) );
  OAI222_X1 U31862 ( .A1(n32017), .A2(n39774), .B1(n32308), .B2(n39768), .C1(
        n31957), .C2(n39762), .ZN(n34176) );
  AOI221_X1 U31863 ( .B1(n39534), .B2(n30029), .C1(n39528), .C2(n30093), .A(
        n35450), .ZN(n35449) );
  OAI222_X1 U31864 ( .A1(n32017), .A2(n39522), .B1(n32308), .B2(n39516), .C1(
        n31957), .C2(n39510), .ZN(n35450) );
  AOI221_X1 U31865 ( .B1(n39786), .B2(n30028), .C1(n39780), .C2(n30092), .A(
        n34195), .ZN(n34194) );
  OAI222_X1 U31866 ( .A1(n32016), .A2(n39774), .B1(n32307), .B2(n39768), .C1(
        n31956), .C2(n39762), .ZN(n34195) );
  AOI221_X1 U31867 ( .B1(n39534), .B2(n30028), .C1(n39528), .C2(n30092), .A(
        n35469), .ZN(n35468) );
  OAI222_X1 U31868 ( .A1(n32016), .A2(n39522), .B1(n32307), .B2(n39516), .C1(
        n31956), .C2(n39510), .ZN(n35469) );
  AOI221_X1 U31869 ( .B1(n39786), .B2(n30027), .C1(n39780), .C2(n30091), .A(
        n34214), .ZN(n34213) );
  OAI222_X1 U31870 ( .A1(n32015), .A2(n39774), .B1(n32306), .B2(n39768), .C1(
        n31955), .C2(n39762), .ZN(n34214) );
  AOI221_X1 U31871 ( .B1(n39534), .B2(n30027), .C1(n39528), .C2(n30091), .A(
        n35488), .ZN(n35487) );
  OAI222_X1 U31872 ( .A1(n32015), .A2(n39522), .B1(n32306), .B2(n39516), .C1(
        n31955), .C2(n39510), .ZN(n35488) );
  AOI221_X1 U31873 ( .B1(n39785), .B2(n30026), .C1(n39779), .C2(n30090), .A(
        n34233), .ZN(n34232) );
  OAI222_X1 U31874 ( .A1(n32014), .A2(n39773), .B1(n32305), .B2(n39767), .C1(
        n31954), .C2(n39761), .ZN(n34233) );
  AOI221_X1 U31875 ( .B1(n39533), .B2(n30026), .C1(n39527), .C2(n30090), .A(
        n35507), .ZN(n35506) );
  OAI222_X1 U31876 ( .A1(n32014), .A2(n39521), .B1(n32305), .B2(n39515), .C1(
        n31954), .C2(n39509), .ZN(n35507) );
  AOI221_X1 U31877 ( .B1(n39785), .B2(n30025), .C1(n39779), .C2(n30089), .A(
        n34252), .ZN(n34251) );
  OAI222_X1 U31878 ( .A1(n32013), .A2(n39773), .B1(n32304), .B2(n39767), .C1(
        n31953), .C2(n39761), .ZN(n34252) );
  AOI221_X1 U31879 ( .B1(n39533), .B2(n30025), .C1(n39527), .C2(n30089), .A(
        n35526), .ZN(n35525) );
  OAI222_X1 U31880 ( .A1(n32013), .A2(n39521), .B1(n32304), .B2(n39515), .C1(
        n31953), .C2(n39509), .ZN(n35526) );
  AOI221_X1 U31881 ( .B1(n39785), .B2(n30024), .C1(n39779), .C2(n30088), .A(
        n34271), .ZN(n34270) );
  OAI222_X1 U31882 ( .A1(n32012), .A2(n39773), .B1(n32303), .B2(n39767), .C1(
        n31952), .C2(n39761), .ZN(n34271) );
  AOI221_X1 U31883 ( .B1(n39533), .B2(n30024), .C1(n39527), .C2(n30088), .A(
        n35545), .ZN(n35544) );
  OAI222_X1 U31884 ( .A1(n32012), .A2(n39521), .B1(n32303), .B2(n39515), .C1(
        n31952), .C2(n39509), .ZN(n35545) );
  AOI221_X1 U31885 ( .B1(n39785), .B2(n30023), .C1(n39779), .C2(n30087), .A(
        n34290), .ZN(n34289) );
  OAI222_X1 U31886 ( .A1(n32011), .A2(n39773), .B1(n32302), .B2(n39767), .C1(
        n31951), .C2(n39761), .ZN(n34290) );
  AOI221_X1 U31887 ( .B1(n39533), .B2(n30023), .C1(n39527), .C2(n30087), .A(
        n35564), .ZN(n35563) );
  OAI222_X1 U31888 ( .A1(n32011), .A2(n39521), .B1(n32302), .B2(n39515), .C1(
        n31951), .C2(n39509), .ZN(n35564) );
  AOI221_X1 U31889 ( .B1(n39785), .B2(n30022), .C1(n39779), .C2(n30086), .A(
        n34309), .ZN(n34308) );
  OAI222_X1 U31890 ( .A1(n32010), .A2(n39773), .B1(n32301), .B2(n39767), .C1(
        n31950), .C2(n39761), .ZN(n34309) );
  AOI221_X1 U31891 ( .B1(n39533), .B2(n30022), .C1(n39527), .C2(n30086), .A(
        n35583), .ZN(n35582) );
  OAI222_X1 U31892 ( .A1(n32010), .A2(n39521), .B1(n32301), .B2(n39515), .C1(
        n31950), .C2(n39509), .ZN(n35583) );
  AOI221_X1 U31893 ( .B1(n39785), .B2(n30021), .C1(n39779), .C2(n30085), .A(
        n34328), .ZN(n34327) );
  OAI222_X1 U31894 ( .A1(n32009), .A2(n39773), .B1(n32300), .B2(n39767), .C1(
        n31949), .C2(n39761), .ZN(n34328) );
  AOI221_X1 U31895 ( .B1(n39533), .B2(n30021), .C1(n39527), .C2(n30085), .A(
        n35602), .ZN(n35601) );
  OAI222_X1 U31896 ( .A1(n32009), .A2(n39521), .B1(n32300), .B2(n39515), .C1(
        n31949), .C2(n39509), .ZN(n35602) );
  AOI221_X1 U31897 ( .B1(n39785), .B2(n30020), .C1(n39779), .C2(n30084), .A(
        n34347), .ZN(n34346) );
  OAI222_X1 U31898 ( .A1(n32008), .A2(n39773), .B1(n32299), .B2(n39767), .C1(
        n31948), .C2(n39761), .ZN(n34347) );
  AOI221_X1 U31899 ( .B1(n39533), .B2(n30020), .C1(n39527), .C2(n30084), .A(
        n35621), .ZN(n35620) );
  OAI222_X1 U31900 ( .A1(n32008), .A2(n39521), .B1(n32299), .B2(n39515), .C1(
        n31948), .C2(n39509), .ZN(n35621) );
  AOI221_X1 U31901 ( .B1(n39785), .B2(n30019), .C1(n39779), .C2(n30083), .A(
        n34366), .ZN(n34365) );
  OAI222_X1 U31902 ( .A1(n32007), .A2(n39773), .B1(n32298), .B2(n39767), .C1(
        n31947), .C2(n39761), .ZN(n34366) );
  AOI221_X1 U31903 ( .B1(n39533), .B2(n30019), .C1(n39527), .C2(n30083), .A(
        n35640), .ZN(n35639) );
  OAI222_X1 U31904 ( .A1(n32007), .A2(n39521), .B1(n32298), .B2(n39515), .C1(
        n31947), .C2(n39509), .ZN(n35640) );
  AOI221_X1 U31905 ( .B1(n39785), .B2(n30018), .C1(n39779), .C2(n30082), .A(
        n34385), .ZN(n34384) );
  OAI222_X1 U31906 ( .A1(n32006), .A2(n39773), .B1(n32297), .B2(n39767), .C1(
        n31946), .C2(n39761), .ZN(n34385) );
  AOI221_X1 U31907 ( .B1(n39533), .B2(n30018), .C1(n39527), .C2(n30082), .A(
        n35659), .ZN(n35658) );
  OAI222_X1 U31908 ( .A1(n32006), .A2(n39521), .B1(n32297), .B2(n39515), .C1(
        n31946), .C2(n39509), .ZN(n35659) );
  AOI221_X1 U31909 ( .B1(n39785), .B2(n30017), .C1(n39779), .C2(n30081), .A(
        n34404), .ZN(n34403) );
  OAI222_X1 U31910 ( .A1(n32005), .A2(n39773), .B1(n32296), .B2(n39767), .C1(
        n31945), .C2(n39761), .ZN(n34404) );
  AOI221_X1 U31911 ( .B1(n39533), .B2(n30017), .C1(n39527), .C2(n30081), .A(
        n35678), .ZN(n35677) );
  OAI222_X1 U31912 ( .A1(n32005), .A2(n39521), .B1(n32296), .B2(n39515), .C1(
        n31945), .C2(n39509), .ZN(n35678) );
  AOI221_X1 U31913 ( .B1(n39785), .B2(n30016), .C1(n39779), .C2(n30080), .A(
        n34423), .ZN(n34422) );
  OAI222_X1 U31914 ( .A1(n32004), .A2(n39773), .B1(n32295), .B2(n39767), .C1(
        n31944), .C2(n39761), .ZN(n34423) );
  AOI221_X1 U31915 ( .B1(n39533), .B2(n30016), .C1(n39527), .C2(n30080), .A(
        n35697), .ZN(n35696) );
  OAI222_X1 U31916 ( .A1(n32004), .A2(n39521), .B1(n32295), .B2(n39515), .C1(
        n31944), .C2(n39509), .ZN(n35697) );
  AOI221_X1 U31917 ( .B1(n39785), .B2(n30015), .C1(n39779), .C2(n30079), .A(
        n34442), .ZN(n34441) );
  OAI222_X1 U31918 ( .A1(n32003), .A2(n39773), .B1(n32294), .B2(n39767), .C1(
        n31943), .C2(n39761), .ZN(n34442) );
  AOI221_X1 U31919 ( .B1(n39533), .B2(n30015), .C1(n39527), .C2(n30079), .A(
        n35716), .ZN(n35715) );
  OAI222_X1 U31920 ( .A1(n32003), .A2(n39521), .B1(n32294), .B2(n39515), .C1(
        n31943), .C2(n39509), .ZN(n35716) );
  AOI221_X1 U31921 ( .B1(n39784), .B2(n30014), .C1(n39778), .C2(n30078), .A(
        n34461), .ZN(n34460) );
  OAI222_X1 U31922 ( .A1(n32002), .A2(n39772), .B1(n32293), .B2(n39766), .C1(
        n31942), .C2(n39760), .ZN(n34461) );
  AOI221_X1 U31923 ( .B1(n39532), .B2(n30014), .C1(n39526), .C2(n30078), .A(
        n35735), .ZN(n35734) );
  OAI222_X1 U31924 ( .A1(n32002), .A2(n39520), .B1(n32293), .B2(n39514), .C1(
        n31942), .C2(n39508), .ZN(n35735) );
  AOI221_X1 U31925 ( .B1(n39784), .B2(n30013), .C1(n39778), .C2(n30077), .A(
        n34480), .ZN(n34479) );
  OAI222_X1 U31926 ( .A1(n32001), .A2(n39772), .B1(n32292), .B2(n39766), .C1(
        n31941), .C2(n39760), .ZN(n34480) );
  AOI221_X1 U31927 ( .B1(n39532), .B2(n30013), .C1(n39526), .C2(n30077), .A(
        n35754), .ZN(n35753) );
  OAI222_X1 U31928 ( .A1(n32001), .A2(n39520), .B1(n32292), .B2(n39514), .C1(
        n31941), .C2(n39508), .ZN(n35754) );
  AOI221_X1 U31929 ( .B1(n39784), .B2(n30012), .C1(n39778), .C2(n30076), .A(
        n34499), .ZN(n34498) );
  OAI222_X1 U31930 ( .A1(n32000), .A2(n39772), .B1(n32291), .B2(n39766), .C1(
        n31940), .C2(n39760), .ZN(n34499) );
  AOI221_X1 U31931 ( .B1(n39532), .B2(n30012), .C1(n39526), .C2(n30076), .A(
        n35773), .ZN(n35772) );
  OAI222_X1 U31932 ( .A1(n32000), .A2(n39520), .B1(n32291), .B2(n39514), .C1(
        n31940), .C2(n39508), .ZN(n35773) );
  AOI221_X1 U31933 ( .B1(n39784), .B2(n30011), .C1(n39778), .C2(n30075), .A(
        n34518), .ZN(n34517) );
  OAI222_X1 U31934 ( .A1(n31999), .A2(n39772), .B1(n32290), .B2(n39766), .C1(
        n31939), .C2(n39760), .ZN(n34518) );
  AOI221_X1 U31935 ( .B1(n39532), .B2(n30011), .C1(n39526), .C2(n30075), .A(
        n35792), .ZN(n35791) );
  OAI222_X1 U31936 ( .A1(n31999), .A2(n39520), .B1(n32290), .B2(n39514), .C1(
        n31939), .C2(n39508), .ZN(n35792) );
  AOI221_X1 U31937 ( .B1(n39784), .B2(n30010), .C1(n39778), .C2(n30074), .A(
        n34537), .ZN(n34536) );
  OAI222_X1 U31938 ( .A1(n31998), .A2(n39772), .B1(n32289), .B2(n39766), .C1(
        n31938), .C2(n39760), .ZN(n34537) );
  AOI221_X1 U31939 ( .B1(n39532), .B2(n30010), .C1(n39526), .C2(n30074), .A(
        n35811), .ZN(n35810) );
  OAI222_X1 U31940 ( .A1(n31998), .A2(n39520), .B1(n32289), .B2(n39514), .C1(
        n31938), .C2(n39508), .ZN(n35811) );
  AOI221_X1 U31941 ( .B1(n39784), .B2(n30009), .C1(n39778), .C2(n30073), .A(
        n34556), .ZN(n34555) );
  OAI222_X1 U31942 ( .A1(n31997), .A2(n39772), .B1(n32288), .B2(n39766), .C1(
        n31937), .C2(n39760), .ZN(n34556) );
  AOI221_X1 U31943 ( .B1(n39532), .B2(n30009), .C1(n39526), .C2(n30073), .A(
        n35830), .ZN(n35829) );
  OAI222_X1 U31944 ( .A1(n31997), .A2(n39520), .B1(n32288), .B2(n39514), .C1(
        n31937), .C2(n39508), .ZN(n35830) );
  AOI221_X1 U31945 ( .B1(n39784), .B2(n30008), .C1(n39778), .C2(n30072), .A(
        n34575), .ZN(n34574) );
  OAI222_X1 U31946 ( .A1(n31996), .A2(n39772), .B1(n32287), .B2(n39766), .C1(
        n31936), .C2(n39760), .ZN(n34575) );
  AOI221_X1 U31947 ( .B1(n39532), .B2(n30008), .C1(n39526), .C2(n30072), .A(
        n35849), .ZN(n35848) );
  OAI222_X1 U31948 ( .A1(n31996), .A2(n39520), .B1(n32287), .B2(n39514), .C1(
        n31936), .C2(n39508), .ZN(n35849) );
  AOI221_X1 U31949 ( .B1(n39784), .B2(n30007), .C1(n39778), .C2(n30071), .A(
        n34594), .ZN(n34593) );
  OAI222_X1 U31950 ( .A1(n31995), .A2(n39772), .B1(n32054), .B2(n39766), .C1(
        n31935), .C2(n39760), .ZN(n34594) );
  AOI221_X1 U31951 ( .B1(n39532), .B2(n30007), .C1(n39526), .C2(n30071), .A(
        n35868), .ZN(n35867) );
  OAI222_X1 U31952 ( .A1(n31995), .A2(n39520), .B1(n32054), .B2(n39514), .C1(
        n31935), .C2(n39508), .ZN(n35868) );
  AOI221_X1 U31953 ( .B1(n39784), .B2(n30006), .C1(n39778), .C2(n30070), .A(
        n34613), .ZN(n34612) );
  OAI222_X1 U31954 ( .A1(n31994), .A2(n39772), .B1(n32286), .B2(n39766), .C1(
        n31934), .C2(n39760), .ZN(n34613) );
  AOI221_X1 U31955 ( .B1(n39532), .B2(n30006), .C1(n39526), .C2(n30070), .A(
        n35887), .ZN(n35886) );
  OAI222_X1 U31956 ( .A1(n31994), .A2(n39520), .B1(n32286), .B2(n39514), .C1(
        n31934), .C2(n39508), .ZN(n35887) );
  AOI221_X1 U31957 ( .B1(n39784), .B2(n30005), .C1(n39778), .C2(n30069), .A(
        n34632), .ZN(n34631) );
  OAI222_X1 U31958 ( .A1(n31993), .A2(n39772), .B1(n32053), .B2(n39766), .C1(
        n31933), .C2(n39760), .ZN(n34632) );
  AOI221_X1 U31959 ( .B1(n39532), .B2(n30005), .C1(n39526), .C2(n30069), .A(
        n35906), .ZN(n35905) );
  OAI222_X1 U31960 ( .A1(n31993), .A2(n39520), .B1(n32053), .B2(n39514), .C1(
        n31933), .C2(n39508), .ZN(n35906) );
  AOI221_X1 U31961 ( .B1(n39784), .B2(n30004), .C1(n39778), .C2(n30068), .A(
        n34651), .ZN(n34650) );
  OAI222_X1 U31962 ( .A1(n31992), .A2(n39772), .B1(n32052), .B2(n39766), .C1(
        n31932), .C2(n39760), .ZN(n34651) );
  AOI221_X1 U31963 ( .B1(n39532), .B2(n30004), .C1(n39526), .C2(n30068), .A(
        n35925), .ZN(n35924) );
  OAI222_X1 U31964 ( .A1(n31992), .A2(n39520), .B1(n32052), .B2(n39514), .C1(
        n31932), .C2(n39508), .ZN(n35925) );
  AOI221_X1 U31965 ( .B1(n39784), .B2(n30003), .C1(n39778), .C2(n30067), .A(
        n34670), .ZN(n34669) );
  OAI222_X1 U31966 ( .A1(n31991), .A2(n39772), .B1(n32051), .B2(n39766), .C1(
        n31931), .C2(n39760), .ZN(n34670) );
  AOI221_X1 U31967 ( .B1(n39532), .B2(n30003), .C1(n39526), .C2(n30067), .A(
        n35944), .ZN(n35943) );
  OAI222_X1 U31968 ( .A1(n31991), .A2(n39520), .B1(n32051), .B2(n39514), .C1(
        n31931), .C2(n39508), .ZN(n35944) );
  AOI221_X1 U31969 ( .B1(n39252), .B2(n29735), .C1(n39246), .C2(n29799), .A(
        n37017), .ZN(n37014) );
  OAI222_X1 U31970 ( .A1(n31863), .A2(n39240), .B1(n31923), .B2(n39234), .C1(
        n31803), .C2(n39228), .ZN(n37017) );
  AOI221_X1 U31971 ( .B1(n39253), .B2(n29734), .C1(n39247), .C2(n29798), .A(
        n36998), .ZN(n36995) );
  OAI222_X1 U31972 ( .A1(n31862), .A2(n39241), .B1(n31922), .B2(n39235), .C1(
        n31802), .C2(n39229), .ZN(n36998) );
  AOI221_X1 U31973 ( .B1(n39253), .B2(n29733), .C1(n39247), .C2(n29797), .A(
        n36979), .ZN(n36976) );
  OAI222_X1 U31974 ( .A1(n31861), .A2(n39241), .B1(n31921), .B2(n39235), .C1(
        n31801), .C2(n39229), .ZN(n36979) );
  AOI221_X1 U31975 ( .B1(n39253), .B2(n29732), .C1(n39247), .C2(n29796), .A(
        n36960), .ZN(n36957) );
  OAI222_X1 U31976 ( .A1(n31860), .A2(n39241), .B1(n31920), .B2(n39235), .C1(
        n31800), .C2(n39229), .ZN(n36960) );
  AOI221_X1 U31977 ( .B1(n39253), .B2(n29731), .C1(n39247), .C2(n29795), .A(
        n36941), .ZN(n36938) );
  OAI222_X1 U31978 ( .A1(n31859), .A2(n39241), .B1(n31919), .B2(n39235), .C1(
        n31799), .C2(n39229), .ZN(n36941) );
  AOI221_X1 U31979 ( .B1(n39253), .B2(n29730), .C1(n39247), .C2(n29794), .A(
        n36922), .ZN(n36919) );
  OAI222_X1 U31980 ( .A1(n31858), .A2(n39241), .B1(n31918), .B2(n39235), .C1(
        n31798), .C2(n39229), .ZN(n36922) );
  AOI221_X1 U31981 ( .B1(n39253), .B2(n29729), .C1(n39247), .C2(n29793), .A(
        n36903), .ZN(n36900) );
  OAI222_X1 U31982 ( .A1(n31857), .A2(n39241), .B1(n31917), .B2(n39235), .C1(
        n31797), .C2(n39229), .ZN(n36903) );
  AOI221_X1 U31983 ( .B1(n39253), .B2(n29728), .C1(n39247), .C2(n29792), .A(
        n36884), .ZN(n36881) );
  OAI222_X1 U31984 ( .A1(n31856), .A2(n39241), .B1(n31916), .B2(n39235), .C1(
        n31796), .C2(n39229), .ZN(n36884) );
  AOI221_X1 U31985 ( .B1(n39253), .B2(n29727), .C1(n39247), .C2(n29791), .A(
        n36865), .ZN(n36862) );
  OAI222_X1 U31986 ( .A1(n31855), .A2(n39241), .B1(n31915), .B2(n39235), .C1(
        n31795), .C2(n39229), .ZN(n36865) );
  AOI221_X1 U31987 ( .B1(n39253), .B2(n29726), .C1(n39247), .C2(n29790), .A(
        n36846), .ZN(n36843) );
  OAI222_X1 U31988 ( .A1(n31854), .A2(n39241), .B1(n31914), .B2(n39235), .C1(
        n31794), .C2(n39229), .ZN(n36846) );
  AOI221_X1 U31989 ( .B1(n39253), .B2(n29725), .C1(n39247), .C2(n29789), .A(
        n36827), .ZN(n36824) );
  OAI222_X1 U31990 ( .A1(n31853), .A2(n39241), .B1(n31913), .B2(n39235), .C1(
        n31793), .C2(n39229), .ZN(n36827) );
  AOI221_X1 U31991 ( .B1(n39253), .B2(n29724), .C1(n39247), .C2(n29788), .A(
        n36808), .ZN(n36805) );
  OAI222_X1 U31992 ( .A1(n31852), .A2(n39241), .B1(n31912), .B2(n39235), .C1(
        n31792), .C2(n39229), .ZN(n36808) );
  AOI221_X1 U31993 ( .B1(n39253), .B2(n29723), .C1(n39247), .C2(n29787), .A(
        n36789), .ZN(n36786) );
  OAI222_X1 U31994 ( .A1(n31851), .A2(n39241), .B1(n31911), .B2(n39235), .C1(
        n31791), .C2(n39229), .ZN(n36789) );
  AOI221_X1 U31995 ( .B1(n39254), .B2(n29722), .C1(n39248), .C2(n29786), .A(
        n36770), .ZN(n36767) );
  OAI222_X1 U31996 ( .A1(n31850), .A2(n39242), .B1(n31910), .B2(n39236), .C1(
        n31790), .C2(n39230), .ZN(n36770) );
  AOI221_X1 U31997 ( .B1(n39254), .B2(n29721), .C1(n39248), .C2(n29785), .A(
        n36751), .ZN(n36748) );
  OAI222_X1 U31998 ( .A1(n31849), .A2(n39242), .B1(n31909), .B2(n39236), .C1(
        n31789), .C2(n39230), .ZN(n36751) );
  AOI221_X1 U31999 ( .B1(n39254), .B2(n29720), .C1(n39248), .C2(n29784), .A(
        n36732), .ZN(n36729) );
  OAI222_X1 U32000 ( .A1(n31848), .A2(n39242), .B1(n31908), .B2(n39236), .C1(
        n31788), .C2(n39230), .ZN(n36732) );
  AOI221_X1 U32001 ( .B1(n39254), .B2(n29719), .C1(n39248), .C2(n29783), .A(
        n36713), .ZN(n36710) );
  OAI222_X1 U32002 ( .A1(n31847), .A2(n39242), .B1(n31907), .B2(n39236), .C1(
        n31787), .C2(n39230), .ZN(n36713) );
  AOI221_X1 U32003 ( .B1(n39254), .B2(n29718), .C1(n39248), .C2(n29782), .A(
        n36694), .ZN(n36691) );
  OAI222_X1 U32004 ( .A1(n31846), .A2(n39242), .B1(n31906), .B2(n39236), .C1(
        n31786), .C2(n39230), .ZN(n36694) );
  AOI221_X1 U32005 ( .B1(n39254), .B2(n29717), .C1(n39248), .C2(n29781), .A(
        n36675), .ZN(n36672) );
  OAI222_X1 U32006 ( .A1(n31845), .A2(n39242), .B1(n31905), .B2(n39236), .C1(
        n31785), .C2(n39230), .ZN(n36675) );
  AOI221_X1 U32007 ( .B1(n39254), .B2(n29716), .C1(n39248), .C2(n29780), .A(
        n36656), .ZN(n36653) );
  OAI222_X1 U32008 ( .A1(n31844), .A2(n39242), .B1(n31904), .B2(n39236), .C1(
        n31784), .C2(n39230), .ZN(n36656) );
  AOI221_X1 U32009 ( .B1(n39254), .B2(n29715), .C1(n39248), .C2(n29779), .A(
        n36637), .ZN(n36634) );
  OAI222_X1 U32010 ( .A1(n31843), .A2(n39242), .B1(n31903), .B2(n39236), .C1(
        n31783), .C2(n39230), .ZN(n36637) );
  AOI221_X1 U32011 ( .B1(n39254), .B2(n29714), .C1(n39248), .C2(n29778), .A(
        n36618), .ZN(n36615) );
  OAI222_X1 U32012 ( .A1(n31842), .A2(n39242), .B1(n31902), .B2(n39236), .C1(
        n31782), .C2(n39230), .ZN(n36618) );
  AOI221_X1 U32013 ( .B1(n39254), .B2(n29713), .C1(n39248), .C2(n29777), .A(
        n36599), .ZN(n36596) );
  OAI222_X1 U32014 ( .A1(n31841), .A2(n39242), .B1(n31901), .B2(n39236), .C1(
        n31781), .C2(n39230), .ZN(n36599) );
  AOI221_X1 U32015 ( .B1(n39254), .B2(n29712), .C1(n39248), .C2(n29776), .A(
        n36580), .ZN(n36577) );
  OAI222_X1 U32016 ( .A1(n31840), .A2(n39242), .B1(n31900), .B2(n39236), .C1(
        n31780), .C2(n39230), .ZN(n36580) );
  AOI221_X1 U32017 ( .B1(n39254), .B2(n29711), .C1(n39248), .C2(n29775), .A(
        n36561), .ZN(n36558) );
  OAI222_X1 U32018 ( .A1(n31839), .A2(n39242), .B1(n31899), .B2(n39236), .C1(
        n31779), .C2(n39230), .ZN(n36561) );
  AOI221_X1 U32019 ( .B1(n39255), .B2(n29710), .C1(n39249), .C2(n29774), .A(
        n36542), .ZN(n36539) );
  OAI222_X1 U32020 ( .A1(n31838), .A2(n39243), .B1(n31898), .B2(n39237), .C1(
        n31778), .C2(n39231), .ZN(n36542) );
  AOI221_X1 U32021 ( .B1(n39255), .B2(n29709), .C1(n39249), .C2(n29773), .A(
        n36523), .ZN(n36520) );
  OAI222_X1 U32022 ( .A1(n31837), .A2(n39243), .B1(n31897), .B2(n39237), .C1(
        n31777), .C2(n39231), .ZN(n36523) );
  AOI221_X1 U32023 ( .B1(n39255), .B2(n29708), .C1(n39249), .C2(n29772), .A(
        n36504), .ZN(n36501) );
  OAI222_X1 U32024 ( .A1(n31836), .A2(n39243), .B1(n31896), .B2(n39237), .C1(
        n31776), .C2(n39231), .ZN(n36504) );
  AOI221_X1 U32025 ( .B1(n39255), .B2(n29707), .C1(n39249), .C2(n29771), .A(
        n36485), .ZN(n36482) );
  OAI222_X1 U32026 ( .A1(n31835), .A2(n39243), .B1(n31895), .B2(n39237), .C1(
        n31775), .C2(n39231), .ZN(n36485) );
  AOI221_X1 U32027 ( .B1(n39255), .B2(n29706), .C1(n39249), .C2(n29770), .A(
        n36466), .ZN(n36463) );
  OAI222_X1 U32028 ( .A1(n31834), .A2(n39243), .B1(n31894), .B2(n39237), .C1(
        n31774), .C2(n39231), .ZN(n36466) );
  AOI221_X1 U32029 ( .B1(n39255), .B2(n29705), .C1(n39249), .C2(n29769), .A(
        n36447), .ZN(n36444) );
  OAI222_X1 U32030 ( .A1(n31833), .A2(n39243), .B1(n31893), .B2(n39237), .C1(
        n31773), .C2(n39231), .ZN(n36447) );
  AOI221_X1 U32031 ( .B1(n39255), .B2(n29704), .C1(n39249), .C2(n29768), .A(
        n36428), .ZN(n36425) );
  OAI222_X1 U32032 ( .A1(n31832), .A2(n39243), .B1(n31892), .B2(n39237), .C1(
        n31772), .C2(n39231), .ZN(n36428) );
  AOI221_X1 U32033 ( .B1(n39255), .B2(n29703), .C1(n39249), .C2(n29767), .A(
        n36409), .ZN(n36406) );
  OAI222_X1 U32034 ( .A1(n31831), .A2(n39243), .B1(n31891), .B2(n39237), .C1(
        n31771), .C2(n39231), .ZN(n36409) );
  AOI221_X1 U32035 ( .B1(n39255), .B2(n29702), .C1(n39249), .C2(n29766), .A(
        n36390), .ZN(n36387) );
  OAI222_X1 U32036 ( .A1(n31830), .A2(n39243), .B1(n31890), .B2(n39237), .C1(
        n31770), .C2(n39231), .ZN(n36390) );
  AOI221_X1 U32037 ( .B1(n39255), .B2(n29701), .C1(n39249), .C2(n29765), .A(
        n36371), .ZN(n36368) );
  OAI222_X1 U32038 ( .A1(n31829), .A2(n39243), .B1(n31889), .B2(n39237), .C1(
        n31769), .C2(n39231), .ZN(n36371) );
  AOI221_X1 U32039 ( .B1(n39255), .B2(n29700), .C1(n39249), .C2(n29764), .A(
        n36352), .ZN(n36349) );
  OAI222_X1 U32040 ( .A1(n31828), .A2(n39243), .B1(n31888), .B2(n39237), .C1(
        n31768), .C2(n39231), .ZN(n36352) );
  AOI221_X1 U32041 ( .B1(n39255), .B2(n29699), .C1(n39249), .C2(n29763), .A(
        n36333), .ZN(n36330) );
  OAI222_X1 U32042 ( .A1(n31827), .A2(n39243), .B1(n31887), .B2(n39237), .C1(
        n31767), .C2(n39231), .ZN(n36333) );
  AOI221_X1 U32043 ( .B1(n39256), .B2(n29698), .C1(n39250), .C2(n29762), .A(
        n36314), .ZN(n36311) );
  OAI222_X1 U32044 ( .A1(n31826), .A2(n39244), .B1(n31886), .B2(n39238), .C1(
        n31766), .C2(n39232), .ZN(n36314) );
  AOI221_X1 U32045 ( .B1(n39256), .B2(n29697), .C1(n39250), .C2(n29761), .A(
        n36295), .ZN(n36292) );
  OAI222_X1 U32046 ( .A1(n31825), .A2(n39244), .B1(n31885), .B2(n39238), .C1(
        n31765), .C2(n39232), .ZN(n36295) );
  AOI221_X1 U32047 ( .B1(n39256), .B2(n29696), .C1(n39250), .C2(n29760), .A(
        n36276), .ZN(n36273) );
  OAI222_X1 U32048 ( .A1(n31824), .A2(n39244), .B1(n31884), .B2(n39238), .C1(
        n31764), .C2(n39232), .ZN(n36276) );
  AOI221_X1 U32049 ( .B1(n39256), .B2(n29695), .C1(n39250), .C2(n29759), .A(
        n36257), .ZN(n36254) );
  OAI222_X1 U32050 ( .A1(n31823), .A2(n39244), .B1(n31883), .B2(n39238), .C1(
        n31763), .C2(n39232), .ZN(n36257) );
  AOI221_X1 U32051 ( .B1(n39256), .B2(n29694), .C1(n39250), .C2(n29758), .A(
        n36238), .ZN(n36235) );
  OAI222_X1 U32052 ( .A1(n31822), .A2(n39244), .B1(n31882), .B2(n39238), .C1(
        n31762), .C2(n39232), .ZN(n36238) );
  AOI221_X1 U32053 ( .B1(n39256), .B2(n29693), .C1(n39250), .C2(n29757), .A(
        n36219), .ZN(n36216) );
  OAI222_X1 U32054 ( .A1(n31821), .A2(n39244), .B1(n31881), .B2(n39238), .C1(
        n31761), .C2(n39232), .ZN(n36219) );
  AOI221_X1 U32055 ( .B1(n39252), .B2(n29745), .C1(n39246), .C2(n29809), .A(
        n37207), .ZN(n37204) );
  OAI222_X1 U32056 ( .A1(n32268), .A2(n39240), .B1(n32272), .B2(n39234), .C1(
        n32276), .C2(n39228), .ZN(n37207) );
  AOI221_X1 U32057 ( .B1(n39252), .B2(n29744), .C1(n39246), .C2(n29808), .A(
        n37188), .ZN(n37185) );
  OAI222_X1 U32058 ( .A1(n32267), .A2(n39240), .B1(n32271), .B2(n39234), .C1(
        n32275), .C2(n39228), .ZN(n37188) );
  AOI221_X1 U32059 ( .B1(n39252), .B2(n29743), .C1(n39246), .C2(n29807), .A(
        n37169), .ZN(n37166) );
  OAI222_X1 U32060 ( .A1(n32266), .A2(n39240), .B1(n32270), .B2(n39234), .C1(
        n32274), .C2(n39228), .ZN(n37169) );
  AOI221_X1 U32061 ( .B1(n39252), .B2(n29742), .C1(n39246), .C2(n29806), .A(
        n37150), .ZN(n37147) );
  OAI222_X1 U32062 ( .A1(n31870), .A2(n39240), .B1(n31930), .B2(n39234), .C1(
        n31810), .C2(n39228), .ZN(n37150) );
  AOI221_X1 U32063 ( .B1(n39252), .B2(n29741), .C1(n39246), .C2(n29805), .A(
        n37131), .ZN(n37128) );
  OAI222_X1 U32064 ( .A1(n31869), .A2(n39240), .B1(n31929), .B2(n39234), .C1(
        n31809), .C2(n39228), .ZN(n37131) );
  AOI221_X1 U32065 ( .B1(n39257), .B2(n29686), .C1(n39251), .C2(n29750), .A(
        n36086), .ZN(n36083) );
  OAI222_X1 U32066 ( .A1(n31814), .A2(n39245), .B1(n31874), .B2(n39239), .C1(
        n31754), .C2(n39233), .ZN(n36086) );
  AOI221_X1 U32067 ( .B1(n39257), .B2(n29685), .C1(n39251), .C2(n29749), .A(
        n36067), .ZN(n36064) );
  OAI222_X1 U32068 ( .A1(n31813), .A2(n39245), .B1(n31873), .B2(n39239), .C1(
        n31753), .C2(n39233), .ZN(n36067) );
  AOI221_X1 U32069 ( .B1(n39257), .B2(n29684), .C1(n39251), .C2(n29748), .A(
        n36048), .ZN(n36045) );
  OAI222_X1 U32070 ( .A1(n31812), .A2(n39245), .B1(n31872), .B2(n39239), .C1(
        n31752), .C2(n39233), .ZN(n36048) );
  AOI221_X1 U32071 ( .B1(n39257), .B2(n29683), .C1(n39251), .C2(n29747), .A(
        n35996), .ZN(n35986) );
  OAI222_X1 U32072 ( .A1(n31811), .A2(n39245), .B1(n31871), .B2(n39239), .C1(
        n31751), .C2(n39233), .ZN(n35996) );
  AOI221_X1 U32073 ( .B1(n39252), .B2(n29746), .C1(n39246), .C2(n29810), .A(
        n37232), .ZN(n37223) );
  OAI222_X1 U32074 ( .A1(n32269), .A2(n39240), .B1(n32273), .B2(n39234), .C1(
        n32277), .C2(n39228), .ZN(n37232) );
  AOI221_X1 U32075 ( .B1(n39252), .B2(n29740), .C1(n39246), .C2(n29804), .A(
        n37112), .ZN(n37109) );
  OAI222_X1 U32076 ( .A1(n31868), .A2(n39240), .B1(n31928), .B2(n39234), .C1(
        n31808), .C2(n39228), .ZN(n37112) );
  AOI221_X1 U32077 ( .B1(n39252), .B2(n29739), .C1(n39246), .C2(n29803), .A(
        n37093), .ZN(n37090) );
  OAI222_X1 U32078 ( .A1(n31867), .A2(n39240), .B1(n31927), .B2(n39234), .C1(
        n31807), .C2(n39228), .ZN(n37093) );
  AOI221_X1 U32079 ( .B1(n39252), .B2(n29738), .C1(n39246), .C2(n29802), .A(
        n37074), .ZN(n37071) );
  OAI222_X1 U32080 ( .A1(n31866), .A2(n39240), .B1(n31926), .B2(n39234), .C1(
        n31806), .C2(n39228), .ZN(n37074) );
  AOI221_X1 U32081 ( .B1(n39252), .B2(n29737), .C1(n39246), .C2(n29801), .A(
        n37055), .ZN(n37052) );
  OAI222_X1 U32082 ( .A1(n31865), .A2(n39240), .B1(n31925), .B2(n39234), .C1(
        n31805), .C2(n39228), .ZN(n37055) );
  AOI221_X1 U32083 ( .B1(n39252), .B2(n29736), .C1(n39246), .C2(n29800), .A(
        n37036), .ZN(n37033) );
  OAI222_X1 U32084 ( .A1(n31864), .A2(n39240), .B1(n31924), .B2(n39234), .C1(
        n31804), .C2(n39228), .ZN(n37036) );
  AOI221_X1 U32085 ( .B1(n39256), .B2(n29692), .C1(n39250), .C2(n29756), .A(
        n36200), .ZN(n36197) );
  OAI222_X1 U32086 ( .A1(n31820), .A2(n39244), .B1(n31880), .B2(n39238), .C1(
        n31760), .C2(n39232), .ZN(n36200) );
  AOI221_X1 U32087 ( .B1(n39256), .B2(n29691), .C1(n39250), .C2(n29755), .A(
        n36181), .ZN(n36178) );
  OAI222_X1 U32088 ( .A1(n31819), .A2(n39244), .B1(n31879), .B2(n39238), .C1(
        n31759), .C2(n39232), .ZN(n36181) );
  AOI221_X1 U32089 ( .B1(n39256), .B2(n29690), .C1(n39250), .C2(n29754), .A(
        n36162), .ZN(n36159) );
  OAI222_X1 U32090 ( .A1(n31818), .A2(n39244), .B1(n31878), .B2(n39238), .C1(
        n31758), .C2(n39232), .ZN(n36162) );
  AOI221_X1 U32091 ( .B1(n39256), .B2(n29689), .C1(n39250), .C2(n29753), .A(
        n36143), .ZN(n36140) );
  OAI222_X1 U32092 ( .A1(n31817), .A2(n39244), .B1(n31877), .B2(n39238), .C1(
        n31757), .C2(n39232), .ZN(n36143) );
  AOI221_X1 U32093 ( .B1(n39256), .B2(n29688), .C1(n39250), .C2(n29752), .A(
        n36124), .ZN(n36121) );
  OAI222_X1 U32094 ( .A1(n31816), .A2(n39244), .B1(n31876), .B2(n39238), .C1(
        n31756), .C2(n39232), .ZN(n36124) );
  AOI221_X1 U32095 ( .B1(n39256), .B2(n29687), .C1(n39250), .C2(n29751), .A(
        n36105), .ZN(n36102) );
  OAI222_X1 U32096 ( .A1(n31815), .A2(n39244), .B1(n31875), .B2(n39238), .C1(
        n31755), .C2(n39232), .ZN(n36105) );
  AOI221_X1 U32097 ( .B1(n39759), .B2(n29746), .C1(n39753), .C2(n29810), .A(
        n33441), .ZN(n33431) );
  OAI222_X1 U32098 ( .A1(n32269), .A2(n39747), .B1(n32273), .B2(n39741), .C1(
        n32277), .C2(n39735), .ZN(n33441) );
  AOI221_X1 U32099 ( .B1(n39507), .B2(n29746), .C1(n39501), .C2(n29810), .A(
        n34715), .ZN(n34705) );
  OAI222_X1 U32100 ( .A1(n32269), .A2(n39495), .B1(n32273), .B2(n39489), .C1(
        n32277), .C2(n39483), .ZN(n34715) );
  AOI221_X1 U32101 ( .B1(n39759), .B2(n29745), .C1(n39753), .C2(n29809), .A(
        n33493), .ZN(n33490) );
  OAI222_X1 U32102 ( .A1(n32268), .A2(n39747), .B1(n32272), .B2(n39741), .C1(
        n32276), .C2(n39735), .ZN(n33493) );
  AOI221_X1 U32103 ( .B1(n39507), .B2(n29745), .C1(n39501), .C2(n29809), .A(
        n34767), .ZN(n34764) );
  OAI222_X1 U32104 ( .A1(n32268), .A2(n39495), .B1(n32272), .B2(n39489), .C1(
        n32276), .C2(n39483), .ZN(n34767) );
  AOI221_X1 U32105 ( .B1(n39759), .B2(n29744), .C1(n39753), .C2(n29808), .A(
        n33512), .ZN(n33509) );
  OAI222_X1 U32106 ( .A1(n32267), .A2(n39747), .B1(n32271), .B2(n39741), .C1(
        n32275), .C2(n39735), .ZN(n33512) );
  AOI221_X1 U32107 ( .B1(n39507), .B2(n29744), .C1(n39501), .C2(n29808), .A(
        n34786), .ZN(n34783) );
  OAI222_X1 U32108 ( .A1(n32267), .A2(n39495), .B1(n32271), .B2(n39489), .C1(
        n32275), .C2(n39483), .ZN(n34786) );
  AOI221_X1 U32109 ( .B1(n39759), .B2(n29743), .C1(n39753), .C2(n29807), .A(
        n33531), .ZN(n33528) );
  OAI222_X1 U32110 ( .A1(n32266), .A2(n39747), .B1(n32270), .B2(n39741), .C1(
        n32274), .C2(n39735), .ZN(n33531) );
  AOI221_X1 U32111 ( .B1(n39507), .B2(n29743), .C1(n39501), .C2(n29807), .A(
        n34805), .ZN(n34802) );
  OAI222_X1 U32112 ( .A1(n32266), .A2(n39495), .B1(n32270), .B2(n39489), .C1(
        n32274), .C2(n39483), .ZN(n34805) );
  AOI221_X1 U32113 ( .B1(n39758), .B2(n29742), .C1(n39752), .C2(n29806), .A(
        n33550), .ZN(n33547) );
  OAI222_X1 U32114 ( .A1(n31870), .A2(n39746), .B1(n31930), .B2(n39740), .C1(
        n31810), .C2(n39734), .ZN(n33550) );
  AOI221_X1 U32115 ( .B1(n39506), .B2(n29742), .C1(n39500), .C2(n29806), .A(
        n34824), .ZN(n34821) );
  OAI222_X1 U32116 ( .A1(n31870), .A2(n39494), .B1(n31930), .B2(n39488), .C1(
        n31810), .C2(n39482), .ZN(n34824) );
  AOI221_X1 U32117 ( .B1(n39758), .B2(n29741), .C1(n39752), .C2(n29805), .A(
        n33569), .ZN(n33566) );
  OAI222_X1 U32118 ( .A1(n31869), .A2(n39746), .B1(n31929), .B2(n39740), .C1(
        n31809), .C2(n39734), .ZN(n33569) );
  AOI221_X1 U32119 ( .B1(n39506), .B2(n29741), .C1(n39500), .C2(n29805), .A(
        n34843), .ZN(n34840) );
  OAI222_X1 U32120 ( .A1(n31869), .A2(n39494), .B1(n31929), .B2(n39488), .C1(
        n31809), .C2(n39482), .ZN(n34843) );
  AOI221_X1 U32121 ( .B1(n39758), .B2(n29740), .C1(n39752), .C2(n29804), .A(
        n33588), .ZN(n33585) );
  OAI222_X1 U32122 ( .A1(n31868), .A2(n39746), .B1(n31928), .B2(n39740), .C1(
        n31808), .C2(n39734), .ZN(n33588) );
  AOI221_X1 U32123 ( .B1(n39506), .B2(n29740), .C1(n39500), .C2(n29804), .A(
        n34862), .ZN(n34859) );
  OAI222_X1 U32124 ( .A1(n31868), .A2(n39494), .B1(n31928), .B2(n39488), .C1(
        n31808), .C2(n39482), .ZN(n34862) );
  AOI221_X1 U32125 ( .B1(n39758), .B2(n29739), .C1(n39752), .C2(n29803), .A(
        n33607), .ZN(n33604) );
  OAI222_X1 U32126 ( .A1(n31867), .A2(n39746), .B1(n31927), .B2(n39740), .C1(
        n31807), .C2(n39734), .ZN(n33607) );
  AOI221_X1 U32127 ( .B1(n39506), .B2(n29739), .C1(n39500), .C2(n29803), .A(
        n34881), .ZN(n34878) );
  OAI222_X1 U32128 ( .A1(n31867), .A2(n39494), .B1(n31927), .B2(n39488), .C1(
        n31807), .C2(n39482), .ZN(n34881) );
  AOI221_X1 U32129 ( .B1(n39758), .B2(n29738), .C1(n39752), .C2(n29802), .A(
        n33626), .ZN(n33623) );
  OAI222_X1 U32130 ( .A1(n31866), .A2(n39746), .B1(n31926), .B2(n39740), .C1(
        n31806), .C2(n39734), .ZN(n33626) );
  AOI221_X1 U32131 ( .B1(n39506), .B2(n29738), .C1(n39500), .C2(n29802), .A(
        n34900), .ZN(n34897) );
  OAI222_X1 U32132 ( .A1(n31866), .A2(n39494), .B1(n31926), .B2(n39488), .C1(
        n31806), .C2(n39482), .ZN(n34900) );
  AOI221_X1 U32133 ( .B1(n39758), .B2(n29737), .C1(n39752), .C2(n29801), .A(
        n33645), .ZN(n33642) );
  OAI222_X1 U32134 ( .A1(n31865), .A2(n39746), .B1(n31925), .B2(n39740), .C1(
        n31805), .C2(n39734), .ZN(n33645) );
  AOI221_X1 U32135 ( .B1(n39506), .B2(n29737), .C1(n39500), .C2(n29801), .A(
        n34919), .ZN(n34916) );
  OAI222_X1 U32136 ( .A1(n31865), .A2(n39494), .B1(n31925), .B2(n39488), .C1(
        n31805), .C2(n39482), .ZN(n34919) );
  AOI221_X1 U32137 ( .B1(n39758), .B2(n29736), .C1(n39752), .C2(n29800), .A(
        n33664), .ZN(n33661) );
  OAI222_X1 U32138 ( .A1(n31864), .A2(n39746), .B1(n31924), .B2(n39740), .C1(
        n31804), .C2(n39734), .ZN(n33664) );
  AOI221_X1 U32139 ( .B1(n39506), .B2(n29736), .C1(n39500), .C2(n29800), .A(
        n34938), .ZN(n34935) );
  OAI222_X1 U32140 ( .A1(n31864), .A2(n39494), .B1(n31924), .B2(n39488), .C1(
        n31804), .C2(n39482), .ZN(n34938) );
  AOI221_X1 U32141 ( .B1(n39758), .B2(n29735), .C1(n39752), .C2(n29799), .A(
        n33683), .ZN(n33680) );
  OAI222_X1 U32142 ( .A1(n31863), .A2(n39746), .B1(n31923), .B2(n39740), .C1(
        n31803), .C2(n39734), .ZN(n33683) );
  AOI221_X1 U32143 ( .B1(n39506), .B2(n29735), .C1(n39500), .C2(n29799), .A(
        n34957), .ZN(n34954) );
  OAI222_X1 U32144 ( .A1(n31863), .A2(n39494), .B1(n31923), .B2(n39488), .C1(
        n31803), .C2(n39482), .ZN(n34957) );
  AOI221_X1 U32145 ( .B1(n39758), .B2(n29734), .C1(n39752), .C2(n29798), .A(
        n33702), .ZN(n33699) );
  OAI222_X1 U32146 ( .A1(n31862), .A2(n39746), .B1(n31922), .B2(n39740), .C1(
        n31802), .C2(n39734), .ZN(n33702) );
  AOI221_X1 U32147 ( .B1(n39506), .B2(n29734), .C1(n39500), .C2(n29798), .A(
        n34976), .ZN(n34973) );
  OAI222_X1 U32148 ( .A1(n31862), .A2(n39494), .B1(n31922), .B2(n39488), .C1(
        n31802), .C2(n39482), .ZN(n34976) );
  AOI221_X1 U32149 ( .B1(n39758), .B2(n29733), .C1(n39752), .C2(n29797), .A(
        n33721), .ZN(n33718) );
  OAI222_X1 U32150 ( .A1(n31861), .A2(n39746), .B1(n31921), .B2(n39740), .C1(
        n31801), .C2(n39734), .ZN(n33721) );
  AOI221_X1 U32151 ( .B1(n39506), .B2(n29733), .C1(n39500), .C2(n29797), .A(
        n34995), .ZN(n34992) );
  OAI222_X1 U32152 ( .A1(n31861), .A2(n39494), .B1(n31921), .B2(n39488), .C1(
        n31801), .C2(n39482), .ZN(n34995) );
  AOI221_X1 U32153 ( .B1(n39758), .B2(n29732), .C1(n39752), .C2(n29796), .A(
        n33740), .ZN(n33737) );
  OAI222_X1 U32154 ( .A1(n31860), .A2(n39746), .B1(n31920), .B2(n39740), .C1(
        n31800), .C2(n39734), .ZN(n33740) );
  AOI221_X1 U32155 ( .B1(n39506), .B2(n29732), .C1(n39500), .C2(n29796), .A(
        n35014), .ZN(n35011) );
  OAI222_X1 U32156 ( .A1(n31860), .A2(n39494), .B1(n31920), .B2(n39488), .C1(
        n31800), .C2(n39482), .ZN(n35014) );
  AOI221_X1 U32157 ( .B1(n39758), .B2(n29731), .C1(n39752), .C2(n29795), .A(
        n33759), .ZN(n33756) );
  OAI222_X1 U32158 ( .A1(n31859), .A2(n39746), .B1(n31919), .B2(n39740), .C1(
        n31799), .C2(n39734), .ZN(n33759) );
  AOI221_X1 U32159 ( .B1(n39506), .B2(n29731), .C1(n39500), .C2(n29795), .A(
        n35033), .ZN(n35030) );
  OAI222_X1 U32160 ( .A1(n31859), .A2(n39494), .B1(n31919), .B2(n39488), .C1(
        n31799), .C2(n39482), .ZN(n35033) );
  AOI221_X1 U32161 ( .B1(n39757), .B2(n29730), .C1(n39751), .C2(n29794), .A(
        n33778), .ZN(n33775) );
  OAI222_X1 U32162 ( .A1(n31858), .A2(n39745), .B1(n31918), .B2(n39739), .C1(
        n31798), .C2(n39733), .ZN(n33778) );
  AOI221_X1 U32163 ( .B1(n39505), .B2(n29730), .C1(n39499), .C2(n29794), .A(
        n35052), .ZN(n35049) );
  OAI222_X1 U32164 ( .A1(n31858), .A2(n39493), .B1(n31918), .B2(n39487), .C1(
        n31798), .C2(n39481), .ZN(n35052) );
  AOI221_X1 U32165 ( .B1(n39757), .B2(n29729), .C1(n39751), .C2(n29793), .A(
        n33797), .ZN(n33794) );
  OAI222_X1 U32166 ( .A1(n31857), .A2(n39745), .B1(n31917), .B2(n39739), .C1(
        n31797), .C2(n39733), .ZN(n33797) );
  AOI221_X1 U32167 ( .B1(n39505), .B2(n29729), .C1(n39499), .C2(n29793), .A(
        n35071), .ZN(n35068) );
  OAI222_X1 U32168 ( .A1(n31857), .A2(n39493), .B1(n31917), .B2(n39487), .C1(
        n31797), .C2(n39481), .ZN(n35071) );
  AOI221_X1 U32169 ( .B1(n39757), .B2(n29728), .C1(n39751), .C2(n29792), .A(
        n33816), .ZN(n33813) );
  OAI222_X1 U32170 ( .A1(n31856), .A2(n39745), .B1(n31916), .B2(n39739), .C1(
        n31796), .C2(n39733), .ZN(n33816) );
  AOI221_X1 U32171 ( .B1(n39505), .B2(n29728), .C1(n39499), .C2(n29792), .A(
        n35090), .ZN(n35087) );
  OAI222_X1 U32172 ( .A1(n31856), .A2(n39493), .B1(n31916), .B2(n39487), .C1(
        n31796), .C2(n39481), .ZN(n35090) );
  AOI221_X1 U32173 ( .B1(n39757), .B2(n29727), .C1(n39751), .C2(n29791), .A(
        n33835), .ZN(n33832) );
  OAI222_X1 U32174 ( .A1(n31855), .A2(n39745), .B1(n31915), .B2(n39739), .C1(
        n31795), .C2(n39733), .ZN(n33835) );
  AOI221_X1 U32175 ( .B1(n39505), .B2(n29727), .C1(n39499), .C2(n29791), .A(
        n35109), .ZN(n35106) );
  OAI222_X1 U32176 ( .A1(n31855), .A2(n39493), .B1(n31915), .B2(n39487), .C1(
        n31795), .C2(n39481), .ZN(n35109) );
  AOI221_X1 U32177 ( .B1(n39757), .B2(n29726), .C1(n39751), .C2(n29790), .A(
        n33854), .ZN(n33851) );
  OAI222_X1 U32178 ( .A1(n31854), .A2(n39745), .B1(n31914), .B2(n39739), .C1(
        n31794), .C2(n39733), .ZN(n33854) );
  AOI221_X1 U32179 ( .B1(n39505), .B2(n29726), .C1(n39499), .C2(n29790), .A(
        n35128), .ZN(n35125) );
  OAI222_X1 U32180 ( .A1(n31854), .A2(n39493), .B1(n31914), .B2(n39487), .C1(
        n31794), .C2(n39481), .ZN(n35128) );
  AOI221_X1 U32181 ( .B1(n39757), .B2(n29725), .C1(n39751), .C2(n29789), .A(
        n33873), .ZN(n33870) );
  OAI222_X1 U32182 ( .A1(n31853), .A2(n39745), .B1(n31913), .B2(n39739), .C1(
        n31793), .C2(n39733), .ZN(n33873) );
  AOI221_X1 U32183 ( .B1(n39505), .B2(n29725), .C1(n39499), .C2(n29789), .A(
        n35147), .ZN(n35144) );
  OAI222_X1 U32184 ( .A1(n31853), .A2(n39493), .B1(n31913), .B2(n39487), .C1(
        n31793), .C2(n39481), .ZN(n35147) );
  AOI221_X1 U32185 ( .B1(n39757), .B2(n29724), .C1(n39751), .C2(n29788), .A(
        n33892), .ZN(n33889) );
  OAI222_X1 U32186 ( .A1(n31852), .A2(n39745), .B1(n31912), .B2(n39739), .C1(
        n31792), .C2(n39733), .ZN(n33892) );
  AOI221_X1 U32187 ( .B1(n39505), .B2(n29724), .C1(n39499), .C2(n29788), .A(
        n35166), .ZN(n35163) );
  OAI222_X1 U32188 ( .A1(n31852), .A2(n39493), .B1(n31912), .B2(n39487), .C1(
        n31792), .C2(n39481), .ZN(n35166) );
  AOI221_X1 U32189 ( .B1(n39757), .B2(n29723), .C1(n39751), .C2(n29787), .A(
        n33911), .ZN(n33908) );
  OAI222_X1 U32190 ( .A1(n31851), .A2(n39745), .B1(n31911), .B2(n39739), .C1(
        n31791), .C2(n39733), .ZN(n33911) );
  AOI221_X1 U32191 ( .B1(n39505), .B2(n29723), .C1(n39499), .C2(n29787), .A(
        n35185), .ZN(n35182) );
  OAI222_X1 U32192 ( .A1(n31851), .A2(n39493), .B1(n31911), .B2(n39487), .C1(
        n31791), .C2(n39481), .ZN(n35185) );
  AOI221_X1 U32193 ( .B1(n39757), .B2(n29722), .C1(n39751), .C2(n29786), .A(
        n33930), .ZN(n33927) );
  OAI222_X1 U32194 ( .A1(n31850), .A2(n39745), .B1(n31910), .B2(n39739), .C1(
        n31790), .C2(n39733), .ZN(n33930) );
  AOI221_X1 U32195 ( .B1(n39505), .B2(n29722), .C1(n39499), .C2(n29786), .A(
        n35204), .ZN(n35201) );
  OAI222_X1 U32196 ( .A1(n31850), .A2(n39493), .B1(n31910), .B2(n39487), .C1(
        n31790), .C2(n39481), .ZN(n35204) );
  AOI221_X1 U32197 ( .B1(n39757), .B2(n29721), .C1(n39751), .C2(n29785), .A(
        n33949), .ZN(n33946) );
  OAI222_X1 U32198 ( .A1(n31849), .A2(n39745), .B1(n31909), .B2(n39739), .C1(
        n31789), .C2(n39733), .ZN(n33949) );
  AOI221_X1 U32199 ( .B1(n39505), .B2(n29721), .C1(n39499), .C2(n29785), .A(
        n35223), .ZN(n35220) );
  OAI222_X1 U32200 ( .A1(n31849), .A2(n39493), .B1(n31909), .B2(n39487), .C1(
        n31789), .C2(n39481), .ZN(n35223) );
  AOI221_X1 U32201 ( .B1(n39757), .B2(n29720), .C1(n39751), .C2(n29784), .A(
        n33968), .ZN(n33965) );
  OAI222_X1 U32202 ( .A1(n31848), .A2(n39745), .B1(n31908), .B2(n39739), .C1(
        n31788), .C2(n39733), .ZN(n33968) );
  AOI221_X1 U32203 ( .B1(n39505), .B2(n29720), .C1(n39499), .C2(n29784), .A(
        n35242), .ZN(n35239) );
  OAI222_X1 U32204 ( .A1(n31848), .A2(n39493), .B1(n31908), .B2(n39487), .C1(
        n31788), .C2(n39481), .ZN(n35242) );
  AOI221_X1 U32205 ( .B1(n39757), .B2(n29719), .C1(n39751), .C2(n29783), .A(
        n33987), .ZN(n33984) );
  OAI222_X1 U32206 ( .A1(n31847), .A2(n39745), .B1(n31907), .B2(n39739), .C1(
        n31787), .C2(n39733), .ZN(n33987) );
  AOI221_X1 U32207 ( .B1(n39505), .B2(n29719), .C1(n39499), .C2(n29783), .A(
        n35261), .ZN(n35258) );
  OAI222_X1 U32208 ( .A1(n31847), .A2(n39493), .B1(n31907), .B2(n39487), .C1(
        n31787), .C2(n39481), .ZN(n35261) );
  AOI221_X1 U32209 ( .B1(n39756), .B2(n29718), .C1(n39750), .C2(n29782), .A(
        n34006), .ZN(n34003) );
  OAI222_X1 U32210 ( .A1(n31846), .A2(n39744), .B1(n31906), .B2(n39738), .C1(
        n31786), .C2(n39732), .ZN(n34006) );
  AOI221_X1 U32211 ( .B1(n39504), .B2(n29718), .C1(n39498), .C2(n29782), .A(
        n35280), .ZN(n35277) );
  OAI222_X1 U32212 ( .A1(n31846), .A2(n39492), .B1(n31906), .B2(n39486), .C1(
        n31786), .C2(n39480), .ZN(n35280) );
  AOI221_X1 U32213 ( .B1(n39756), .B2(n29717), .C1(n39750), .C2(n29781), .A(
        n34025), .ZN(n34022) );
  OAI222_X1 U32214 ( .A1(n31845), .A2(n39744), .B1(n31905), .B2(n39738), .C1(
        n31785), .C2(n39732), .ZN(n34025) );
  AOI221_X1 U32215 ( .B1(n39504), .B2(n29717), .C1(n39498), .C2(n29781), .A(
        n35299), .ZN(n35296) );
  OAI222_X1 U32216 ( .A1(n31845), .A2(n39492), .B1(n31905), .B2(n39486), .C1(
        n31785), .C2(n39480), .ZN(n35299) );
  AOI221_X1 U32217 ( .B1(n39756), .B2(n29716), .C1(n39750), .C2(n29780), .A(
        n34044), .ZN(n34041) );
  OAI222_X1 U32218 ( .A1(n31844), .A2(n39744), .B1(n31904), .B2(n39738), .C1(
        n31784), .C2(n39732), .ZN(n34044) );
  AOI221_X1 U32219 ( .B1(n39504), .B2(n29716), .C1(n39498), .C2(n29780), .A(
        n35318), .ZN(n35315) );
  OAI222_X1 U32220 ( .A1(n31844), .A2(n39492), .B1(n31904), .B2(n39486), .C1(
        n31784), .C2(n39480), .ZN(n35318) );
  AOI221_X1 U32221 ( .B1(n39756), .B2(n29715), .C1(n39750), .C2(n29779), .A(
        n34063), .ZN(n34060) );
  OAI222_X1 U32222 ( .A1(n31843), .A2(n39744), .B1(n31903), .B2(n39738), .C1(
        n31783), .C2(n39732), .ZN(n34063) );
  AOI221_X1 U32223 ( .B1(n39504), .B2(n29715), .C1(n39498), .C2(n29779), .A(
        n35337), .ZN(n35334) );
  OAI222_X1 U32224 ( .A1(n31843), .A2(n39492), .B1(n31903), .B2(n39486), .C1(
        n31783), .C2(n39480), .ZN(n35337) );
  AOI221_X1 U32225 ( .B1(n39756), .B2(n29714), .C1(n39750), .C2(n29778), .A(
        n34082), .ZN(n34079) );
  OAI222_X1 U32226 ( .A1(n31842), .A2(n39744), .B1(n31902), .B2(n39738), .C1(
        n31782), .C2(n39732), .ZN(n34082) );
  AOI221_X1 U32227 ( .B1(n39504), .B2(n29714), .C1(n39498), .C2(n29778), .A(
        n35356), .ZN(n35353) );
  OAI222_X1 U32228 ( .A1(n31842), .A2(n39492), .B1(n31902), .B2(n39486), .C1(
        n31782), .C2(n39480), .ZN(n35356) );
  AOI221_X1 U32229 ( .B1(n39756), .B2(n29713), .C1(n39750), .C2(n29777), .A(
        n34101), .ZN(n34098) );
  OAI222_X1 U32230 ( .A1(n31841), .A2(n39744), .B1(n31901), .B2(n39738), .C1(
        n31781), .C2(n39732), .ZN(n34101) );
  AOI221_X1 U32231 ( .B1(n39504), .B2(n29713), .C1(n39498), .C2(n29777), .A(
        n35375), .ZN(n35372) );
  OAI222_X1 U32232 ( .A1(n31841), .A2(n39492), .B1(n31901), .B2(n39486), .C1(
        n31781), .C2(n39480), .ZN(n35375) );
  AOI221_X1 U32233 ( .B1(n39756), .B2(n29712), .C1(n39750), .C2(n29776), .A(
        n34120), .ZN(n34117) );
  OAI222_X1 U32234 ( .A1(n31840), .A2(n39744), .B1(n31900), .B2(n39738), .C1(
        n31780), .C2(n39732), .ZN(n34120) );
  AOI221_X1 U32235 ( .B1(n39504), .B2(n29712), .C1(n39498), .C2(n29776), .A(
        n35394), .ZN(n35391) );
  OAI222_X1 U32236 ( .A1(n31840), .A2(n39492), .B1(n31900), .B2(n39486), .C1(
        n31780), .C2(n39480), .ZN(n35394) );
  AOI221_X1 U32237 ( .B1(n39756), .B2(n29711), .C1(n39750), .C2(n29775), .A(
        n34139), .ZN(n34136) );
  OAI222_X1 U32238 ( .A1(n31839), .A2(n39744), .B1(n31899), .B2(n39738), .C1(
        n31779), .C2(n39732), .ZN(n34139) );
  AOI221_X1 U32239 ( .B1(n39504), .B2(n29711), .C1(n39498), .C2(n29775), .A(
        n35413), .ZN(n35410) );
  OAI222_X1 U32240 ( .A1(n31839), .A2(n39492), .B1(n31899), .B2(n39486), .C1(
        n31779), .C2(n39480), .ZN(n35413) );
  AOI221_X1 U32241 ( .B1(n39756), .B2(n29710), .C1(n39750), .C2(n29774), .A(
        n34158), .ZN(n34155) );
  OAI222_X1 U32242 ( .A1(n31838), .A2(n39744), .B1(n31898), .B2(n39738), .C1(
        n31778), .C2(n39732), .ZN(n34158) );
  AOI221_X1 U32243 ( .B1(n39504), .B2(n29710), .C1(n39498), .C2(n29774), .A(
        n35432), .ZN(n35429) );
  OAI222_X1 U32244 ( .A1(n31838), .A2(n39492), .B1(n31898), .B2(n39486), .C1(
        n31778), .C2(n39480), .ZN(n35432) );
  AOI221_X1 U32245 ( .B1(n39756), .B2(n29709), .C1(n39750), .C2(n29773), .A(
        n34177), .ZN(n34174) );
  OAI222_X1 U32246 ( .A1(n31837), .A2(n39744), .B1(n31897), .B2(n39738), .C1(
        n31777), .C2(n39732), .ZN(n34177) );
  AOI221_X1 U32247 ( .B1(n39504), .B2(n29709), .C1(n39498), .C2(n29773), .A(
        n35451), .ZN(n35448) );
  OAI222_X1 U32248 ( .A1(n31837), .A2(n39492), .B1(n31897), .B2(n39486), .C1(
        n31777), .C2(n39480), .ZN(n35451) );
  AOI221_X1 U32249 ( .B1(n39756), .B2(n29708), .C1(n39750), .C2(n29772), .A(
        n34196), .ZN(n34193) );
  OAI222_X1 U32250 ( .A1(n31836), .A2(n39744), .B1(n31896), .B2(n39738), .C1(
        n31776), .C2(n39732), .ZN(n34196) );
  AOI221_X1 U32251 ( .B1(n39504), .B2(n29708), .C1(n39498), .C2(n29772), .A(
        n35470), .ZN(n35467) );
  OAI222_X1 U32252 ( .A1(n31836), .A2(n39492), .B1(n31896), .B2(n39486), .C1(
        n31776), .C2(n39480), .ZN(n35470) );
  AOI221_X1 U32253 ( .B1(n39756), .B2(n29707), .C1(n39750), .C2(n29771), .A(
        n34215), .ZN(n34212) );
  OAI222_X1 U32254 ( .A1(n31835), .A2(n39744), .B1(n31895), .B2(n39738), .C1(
        n31775), .C2(n39732), .ZN(n34215) );
  AOI221_X1 U32255 ( .B1(n39504), .B2(n29707), .C1(n39498), .C2(n29771), .A(
        n35489), .ZN(n35486) );
  OAI222_X1 U32256 ( .A1(n31835), .A2(n39492), .B1(n31895), .B2(n39486), .C1(
        n31775), .C2(n39480), .ZN(n35489) );
  AOI221_X1 U32257 ( .B1(n39755), .B2(n29706), .C1(n39749), .C2(n29770), .A(
        n34234), .ZN(n34231) );
  OAI222_X1 U32258 ( .A1(n31834), .A2(n39743), .B1(n31894), .B2(n39737), .C1(
        n31774), .C2(n39731), .ZN(n34234) );
  AOI221_X1 U32259 ( .B1(n39503), .B2(n29706), .C1(n39497), .C2(n29770), .A(
        n35508), .ZN(n35505) );
  OAI222_X1 U32260 ( .A1(n31834), .A2(n39491), .B1(n31894), .B2(n39485), .C1(
        n31774), .C2(n39479), .ZN(n35508) );
  AOI221_X1 U32261 ( .B1(n39755), .B2(n29705), .C1(n39749), .C2(n29769), .A(
        n34253), .ZN(n34250) );
  OAI222_X1 U32262 ( .A1(n31833), .A2(n39743), .B1(n31893), .B2(n39737), .C1(
        n31773), .C2(n39731), .ZN(n34253) );
  AOI221_X1 U32263 ( .B1(n39503), .B2(n29705), .C1(n39497), .C2(n29769), .A(
        n35527), .ZN(n35524) );
  OAI222_X1 U32264 ( .A1(n31833), .A2(n39491), .B1(n31893), .B2(n39485), .C1(
        n31773), .C2(n39479), .ZN(n35527) );
  AOI221_X1 U32265 ( .B1(n39755), .B2(n29704), .C1(n39749), .C2(n29768), .A(
        n34272), .ZN(n34269) );
  OAI222_X1 U32266 ( .A1(n31832), .A2(n39743), .B1(n31892), .B2(n39737), .C1(
        n31772), .C2(n39731), .ZN(n34272) );
  AOI221_X1 U32267 ( .B1(n39503), .B2(n29704), .C1(n39497), .C2(n29768), .A(
        n35546), .ZN(n35543) );
  OAI222_X1 U32268 ( .A1(n31832), .A2(n39491), .B1(n31892), .B2(n39485), .C1(
        n31772), .C2(n39479), .ZN(n35546) );
  AOI221_X1 U32269 ( .B1(n39755), .B2(n29703), .C1(n39749), .C2(n29767), .A(
        n34291), .ZN(n34288) );
  OAI222_X1 U32270 ( .A1(n31831), .A2(n39743), .B1(n31891), .B2(n39737), .C1(
        n31771), .C2(n39731), .ZN(n34291) );
  AOI221_X1 U32271 ( .B1(n39503), .B2(n29703), .C1(n39497), .C2(n29767), .A(
        n35565), .ZN(n35562) );
  OAI222_X1 U32272 ( .A1(n31831), .A2(n39491), .B1(n31891), .B2(n39485), .C1(
        n31771), .C2(n39479), .ZN(n35565) );
  AOI221_X1 U32273 ( .B1(n39755), .B2(n29702), .C1(n39749), .C2(n29766), .A(
        n34310), .ZN(n34307) );
  OAI222_X1 U32274 ( .A1(n31830), .A2(n39743), .B1(n31890), .B2(n39737), .C1(
        n31770), .C2(n39731), .ZN(n34310) );
  AOI221_X1 U32275 ( .B1(n39503), .B2(n29702), .C1(n39497), .C2(n29766), .A(
        n35584), .ZN(n35581) );
  OAI222_X1 U32276 ( .A1(n31830), .A2(n39491), .B1(n31890), .B2(n39485), .C1(
        n31770), .C2(n39479), .ZN(n35584) );
  AOI221_X1 U32277 ( .B1(n39755), .B2(n29701), .C1(n39749), .C2(n29765), .A(
        n34329), .ZN(n34326) );
  OAI222_X1 U32278 ( .A1(n31829), .A2(n39743), .B1(n31889), .B2(n39737), .C1(
        n31769), .C2(n39731), .ZN(n34329) );
  AOI221_X1 U32279 ( .B1(n39503), .B2(n29701), .C1(n39497), .C2(n29765), .A(
        n35603), .ZN(n35600) );
  OAI222_X1 U32280 ( .A1(n31829), .A2(n39491), .B1(n31889), .B2(n39485), .C1(
        n31769), .C2(n39479), .ZN(n35603) );
  AOI221_X1 U32281 ( .B1(n39755), .B2(n29700), .C1(n39749), .C2(n29764), .A(
        n34348), .ZN(n34345) );
  OAI222_X1 U32282 ( .A1(n31828), .A2(n39743), .B1(n31888), .B2(n39737), .C1(
        n31768), .C2(n39731), .ZN(n34348) );
  AOI221_X1 U32283 ( .B1(n39503), .B2(n29700), .C1(n39497), .C2(n29764), .A(
        n35622), .ZN(n35619) );
  OAI222_X1 U32284 ( .A1(n31828), .A2(n39491), .B1(n31888), .B2(n39485), .C1(
        n31768), .C2(n39479), .ZN(n35622) );
  AOI221_X1 U32285 ( .B1(n39755), .B2(n29699), .C1(n39749), .C2(n29763), .A(
        n34367), .ZN(n34364) );
  OAI222_X1 U32286 ( .A1(n31827), .A2(n39743), .B1(n31887), .B2(n39737), .C1(
        n31767), .C2(n39731), .ZN(n34367) );
  AOI221_X1 U32287 ( .B1(n39503), .B2(n29699), .C1(n39497), .C2(n29763), .A(
        n35641), .ZN(n35638) );
  OAI222_X1 U32288 ( .A1(n31827), .A2(n39491), .B1(n31887), .B2(n39485), .C1(
        n31767), .C2(n39479), .ZN(n35641) );
  AOI221_X1 U32289 ( .B1(n39755), .B2(n29698), .C1(n39749), .C2(n29762), .A(
        n34386), .ZN(n34383) );
  OAI222_X1 U32290 ( .A1(n31826), .A2(n39743), .B1(n31886), .B2(n39737), .C1(
        n31766), .C2(n39731), .ZN(n34386) );
  AOI221_X1 U32291 ( .B1(n39503), .B2(n29698), .C1(n39497), .C2(n29762), .A(
        n35660), .ZN(n35657) );
  OAI222_X1 U32292 ( .A1(n31826), .A2(n39491), .B1(n31886), .B2(n39485), .C1(
        n31766), .C2(n39479), .ZN(n35660) );
  AOI221_X1 U32293 ( .B1(n39755), .B2(n29697), .C1(n39749), .C2(n29761), .A(
        n34405), .ZN(n34402) );
  OAI222_X1 U32294 ( .A1(n31825), .A2(n39743), .B1(n31885), .B2(n39737), .C1(
        n31765), .C2(n39731), .ZN(n34405) );
  AOI221_X1 U32295 ( .B1(n39503), .B2(n29697), .C1(n39497), .C2(n29761), .A(
        n35679), .ZN(n35676) );
  OAI222_X1 U32296 ( .A1(n31825), .A2(n39491), .B1(n31885), .B2(n39485), .C1(
        n31765), .C2(n39479), .ZN(n35679) );
  AOI221_X1 U32297 ( .B1(n39755), .B2(n29696), .C1(n39749), .C2(n29760), .A(
        n34424), .ZN(n34421) );
  OAI222_X1 U32298 ( .A1(n31824), .A2(n39743), .B1(n31884), .B2(n39737), .C1(
        n31764), .C2(n39731), .ZN(n34424) );
  AOI221_X1 U32299 ( .B1(n39503), .B2(n29696), .C1(n39497), .C2(n29760), .A(
        n35698), .ZN(n35695) );
  OAI222_X1 U32300 ( .A1(n31824), .A2(n39491), .B1(n31884), .B2(n39485), .C1(
        n31764), .C2(n39479), .ZN(n35698) );
  AOI221_X1 U32301 ( .B1(n39755), .B2(n29695), .C1(n39749), .C2(n29759), .A(
        n34443), .ZN(n34440) );
  OAI222_X1 U32302 ( .A1(n31823), .A2(n39743), .B1(n31883), .B2(n39737), .C1(
        n31763), .C2(n39731), .ZN(n34443) );
  AOI221_X1 U32303 ( .B1(n39503), .B2(n29695), .C1(n39497), .C2(n29759), .A(
        n35717), .ZN(n35714) );
  OAI222_X1 U32304 ( .A1(n31823), .A2(n39491), .B1(n31883), .B2(n39485), .C1(
        n31763), .C2(n39479), .ZN(n35717) );
  AOI221_X1 U32305 ( .B1(n39754), .B2(n29694), .C1(n39748), .C2(n29758), .A(
        n34462), .ZN(n34459) );
  OAI222_X1 U32306 ( .A1(n31822), .A2(n39742), .B1(n31882), .B2(n39736), .C1(
        n31762), .C2(n39730), .ZN(n34462) );
  AOI221_X1 U32307 ( .B1(n39502), .B2(n29694), .C1(n39496), .C2(n29758), .A(
        n35736), .ZN(n35733) );
  OAI222_X1 U32308 ( .A1(n31822), .A2(n39490), .B1(n31882), .B2(n39484), .C1(
        n31762), .C2(n39478), .ZN(n35736) );
  AOI221_X1 U32309 ( .B1(n39754), .B2(n29693), .C1(n39748), .C2(n29757), .A(
        n34481), .ZN(n34478) );
  OAI222_X1 U32310 ( .A1(n31821), .A2(n39742), .B1(n31881), .B2(n39736), .C1(
        n31761), .C2(n39730), .ZN(n34481) );
  AOI221_X1 U32311 ( .B1(n39502), .B2(n29693), .C1(n39496), .C2(n29757), .A(
        n35755), .ZN(n35752) );
  OAI222_X1 U32312 ( .A1(n31821), .A2(n39490), .B1(n31881), .B2(n39484), .C1(
        n31761), .C2(n39478), .ZN(n35755) );
  AOI221_X1 U32313 ( .B1(n39754), .B2(n29692), .C1(n39748), .C2(n29756), .A(
        n34500), .ZN(n34497) );
  OAI222_X1 U32314 ( .A1(n31820), .A2(n39742), .B1(n31880), .B2(n39736), .C1(
        n31760), .C2(n39730), .ZN(n34500) );
  AOI221_X1 U32315 ( .B1(n39502), .B2(n29692), .C1(n39496), .C2(n29756), .A(
        n35774), .ZN(n35771) );
  OAI222_X1 U32316 ( .A1(n31820), .A2(n39490), .B1(n31880), .B2(n39484), .C1(
        n31760), .C2(n39478), .ZN(n35774) );
  AOI221_X1 U32317 ( .B1(n39754), .B2(n29691), .C1(n39748), .C2(n29755), .A(
        n34519), .ZN(n34516) );
  OAI222_X1 U32318 ( .A1(n31819), .A2(n39742), .B1(n31879), .B2(n39736), .C1(
        n31759), .C2(n39730), .ZN(n34519) );
  AOI221_X1 U32319 ( .B1(n39502), .B2(n29691), .C1(n39496), .C2(n29755), .A(
        n35793), .ZN(n35790) );
  OAI222_X1 U32320 ( .A1(n31819), .A2(n39490), .B1(n31879), .B2(n39484), .C1(
        n31759), .C2(n39478), .ZN(n35793) );
  AOI221_X1 U32321 ( .B1(n39754), .B2(n29690), .C1(n39748), .C2(n29754), .A(
        n34538), .ZN(n34535) );
  OAI222_X1 U32322 ( .A1(n31818), .A2(n39742), .B1(n31878), .B2(n39736), .C1(
        n31758), .C2(n39730), .ZN(n34538) );
  AOI221_X1 U32323 ( .B1(n39502), .B2(n29690), .C1(n39496), .C2(n29754), .A(
        n35812), .ZN(n35809) );
  OAI222_X1 U32324 ( .A1(n31818), .A2(n39490), .B1(n31878), .B2(n39484), .C1(
        n31758), .C2(n39478), .ZN(n35812) );
  AOI221_X1 U32325 ( .B1(n39754), .B2(n29689), .C1(n39748), .C2(n29753), .A(
        n34557), .ZN(n34554) );
  OAI222_X1 U32326 ( .A1(n31817), .A2(n39742), .B1(n31877), .B2(n39736), .C1(
        n31757), .C2(n39730), .ZN(n34557) );
  AOI221_X1 U32327 ( .B1(n39502), .B2(n29689), .C1(n39496), .C2(n29753), .A(
        n35831), .ZN(n35828) );
  OAI222_X1 U32328 ( .A1(n31817), .A2(n39490), .B1(n31877), .B2(n39484), .C1(
        n31757), .C2(n39478), .ZN(n35831) );
  AOI221_X1 U32329 ( .B1(n39754), .B2(n29688), .C1(n39748), .C2(n29752), .A(
        n34576), .ZN(n34573) );
  OAI222_X1 U32330 ( .A1(n31816), .A2(n39742), .B1(n31876), .B2(n39736), .C1(
        n31756), .C2(n39730), .ZN(n34576) );
  AOI221_X1 U32331 ( .B1(n39502), .B2(n29688), .C1(n39496), .C2(n29752), .A(
        n35850), .ZN(n35847) );
  OAI222_X1 U32332 ( .A1(n31816), .A2(n39490), .B1(n31876), .B2(n39484), .C1(
        n31756), .C2(n39478), .ZN(n35850) );
  AOI221_X1 U32333 ( .B1(n39754), .B2(n29687), .C1(n39748), .C2(n29751), .A(
        n34595), .ZN(n34592) );
  OAI222_X1 U32334 ( .A1(n31815), .A2(n39742), .B1(n31875), .B2(n39736), .C1(
        n31755), .C2(n39730), .ZN(n34595) );
  AOI221_X1 U32335 ( .B1(n39502), .B2(n29687), .C1(n39496), .C2(n29751), .A(
        n35869), .ZN(n35866) );
  OAI222_X1 U32336 ( .A1(n31815), .A2(n39490), .B1(n31875), .B2(n39484), .C1(
        n31755), .C2(n39478), .ZN(n35869) );
  AOI221_X1 U32337 ( .B1(n39754), .B2(n29686), .C1(n39748), .C2(n29750), .A(
        n34614), .ZN(n34611) );
  OAI222_X1 U32338 ( .A1(n31814), .A2(n39742), .B1(n31874), .B2(n39736), .C1(
        n31754), .C2(n39730), .ZN(n34614) );
  AOI221_X1 U32339 ( .B1(n39502), .B2(n29686), .C1(n39496), .C2(n29750), .A(
        n35888), .ZN(n35885) );
  OAI222_X1 U32340 ( .A1(n31814), .A2(n39490), .B1(n31874), .B2(n39484), .C1(
        n31754), .C2(n39478), .ZN(n35888) );
  AOI221_X1 U32341 ( .B1(n39754), .B2(n29685), .C1(n39748), .C2(n29749), .A(
        n34633), .ZN(n34630) );
  OAI222_X1 U32342 ( .A1(n31813), .A2(n39742), .B1(n31873), .B2(n39736), .C1(
        n31753), .C2(n39730), .ZN(n34633) );
  AOI221_X1 U32343 ( .B1(n39502), .B2(n29685), .C1(n39496), .C2(n29749), .A(
        n35907), .ZN(n35904) );
  OAI222_X1 U32344 ( .A1(n31813), .A2(n39490), .B1(n31873), .B2(n39484), .C1(
        n31753), .C2(n39478), .ZN(n35907) );
  AOI221_X1 U32345 ( .B1(n39754), .B2(n29684), .C1(n39748), .C2(n29748), .A(
        n34652), .ZN(n34649) );
  OAI222_X1 U32346 ( .A1(n31812), .A2(n39742), .B1(n31872), .B2(n39736), .C1(
        n31752), .C2(n39730), .ZN(n34652) );
  AOI221_X1 U32347 ( .B1(n39502), .B2(n29684), .C1(n39496), .C2(n29748), .A(
        n35926), .ZN(n35923) );
  OAI222_X1 U32348 ( .A1(n31812), .A2(n39490), .B1(n31872), .B2(n39484), .C1(
        n31752), .C2(n39478), .ZN(n35926) );
  AOI221_X1 U32349 ( .B1(n39754), .B2(n29683), .C1(n39748), .C2(n29747), .A(
        n34677), .ZN(n34668) );
  OAI222_X1 U32350 ( .A1(n31811), .A2(n39742), .B1(n31871), .B2(n39736), .C1(
        n31751), .C2(n39730), .ZN(n34677) );
  AOI221_X1 U32351 ( .B1(n39502), .B2(n29683), .C1(n39496), .C2(n29747), .A(
        n35951), .ZN(n35942) );
  OAI222_X1 U32352 ( .A1(n31811), .A2(n39490), .B1(n31871), .B2(n39484), .C1(
        n31751), .C2(n39478), .ZN(n35951) );
  OAI222_X1 U32353 ( .A1(n40910), .A2(n39914), .B1(n41294), .B2(n39907), .C1(
        n390), .C2(n39901), .ZN(n7662) );
  OAI222_X1 U32354 ( .A1(n40916), .A2(n39914), .B1(n41300), .B2(n39907), .C1(
        n389), .C2(n39901), .ZN(n7661) );
  OAI222_X1 U32355 ( .A1(n40922), .A2(n39914), .B1(n41306), .B2(n39907), .C1(
        n388), .C2(n39901), .ZN(n7660) );
  OAI222_X1 U32356 ( .A1(n40928), .A2(n39914), .B1(n41312), .B2(n39907), .C1(
        n387), .C2(n39901), .ZN(n7659) );
  OAI222_X1 U32357 ( .A1(n40934), .A2(n39914), .B1(n41318), .B2(n39907), .C1(
        n386), .C2(n39901), .ZN(n7658) );
  OAI222_X1 U32358 ( .A1(n40940), .A2(n39914), .B1(n41324), .B2(n39907), .C1(
        n385), .C2(n39901), .ZN(n7657) );
  OAI222_X1 U32359 ( .A1(n40946), .A2(n39914), .B1(n41330), .B2(n39907), .C1(
        n384), .C2(n39901), .ZN(n7656) );
  OAI222_X1 U32360 ( .A1(n40952), .A2(n39914), .B1(n41336), .B2(n39907), .C1(
        n383), .C2(n39901), .ZN(n7655) );
  OAI222_X1 U32361 ( .A1(n40958), .A2(n39914), .B1(n41342), .B2(n39907), .C1(
        n382), .C2(n39901), .ZN(n7654) );
  OAI222_X1 U32362 ( .A1(n40964), .A2(n39914), .B1(n41348), .B2(n39907), .C1(
        n381), .C2(n39901), .ZN(n7653) );
  OAI222_X1 U32363 ( .A1(n40970), .A2(n39914), .B1(n41354), .B2(n39907), .C1(
        n380), .C2(n39901), .ZN(n7652) );
  OAI222_X1 U32364 ( .A1(n40976), .A2(n39914), .B1(n41360), .B2(n39907), .C1(
        n379), .C2(n39901), .ZN(n7651) );
  OAI222_X1 U32365 ( .A1(n40910), .A2(n39933), .B1(n41294), .B2(n39926), .C1(
        n454), .C2(n39920), .ZN(n7726) );
  OAI222_X1 U32366 ( .A1(n40916), .A2(n39933), .B1(n41300), .B2(n39926), .C1(
        n453), .C2(n39920), .ZN(n7725) );
  OAI222_X1 U32367 ( .A1(n40922), .A2(n39933), .B1(n41306), .B2(n39926), .C1(
        n452), .C2(n39920), .ZN(n7724) );
  OAI222_X1 U32368 ( .A1(n40928), .A2(n39933), .B1(n41312), .B2(n39926), .C1(
        n451), .C2(n39920), .ZN(n7723) );
  OAI222_X1 U32369 ( .A1(n40934), .A2(n39933), .B1(n41318), .B2(n39926), .C1(
        n450), .C2(n39920), .ZN(n7722) );
  OAI222_X1 U32370 ( .A1(n40940), .A2(n39933), .B1(n41324), .B2(n39926), .C1(
        n449), .C2(n39920), .ZN(n7721) );
  OAI222_X1 U32371 ( .A1(n40946), .A2(n39933), .B1(n41330), .B2(n39926), .C1(
        n448), .C2(n39920), .ZN(n7720) );
  OAI222_X1 U32372 ( .A1(n40952), .A2(n39933), .B1(n41336), .B2(n39926), .C1(
        n447), .C2(n39920), .ZN(n7719) );
  OAI222_X1 U32373 ( .A1(n40958), .A2(n39933), .B1(n41342), .B2(n39926), .C1(
        n446), .C2(n39920), .ZN(n7718) );
  OAI222_X1 U32374 ( .A1(n40964), .A2(n39933), .B1(n41348), .B2(n39926), .C1(
        n445), .C2(n39920), .ZN(n7717) );
  OAI222_X1 U32375 ( .A1(n40970), .A2(n39933), .B1(n41354), .B2(n39926), .C1(
        n444), .C2(n39920), .ZN(n7716) );
  OAI222_X1 U32376 ( .A1(n40976), .A2(n39933), .B1(n41360), .B2(n39926), .C1(
        n443), .C2(n39920), .ZN(n7715) );
  OAI222_X1 U32377 ( .A1(n40622), .A2(n39918), .B1(n41006), .B2(n39911), .C1(
        n438), .C2(n39905), .ZN(n7710) );
  OAI222_X1 U32378 ( .A1(n40628), .A2(n39918), .B1(n41012), .B2(n39911), .C1(
        n437), .C2(n39905), .ZN(n7709) );
  OAI222_X1 U32379 ( .A1(n40634), .A2(n39918), .B1(n41018), .B2(n39911), .C1(
        n436), .C2(n39905), .ZN(n7708) );
  OAI222_X1 U32380 ( .A1(n40640), .A2(n39918), .B1(n41024), .B2(n39911), .C1(
        n435), .C2(n39905), .ZN(n7707) );
  OAI222_X1 U32381 ( .A1(n40646), .A2(n39918), .B1(n41030), .B2(n39911), .C1(
        n434), .C2(n39905), .ZN(n7706) );
  OAI222_X1 U32382 ( .A1(n40652), .A2(n39918), .B1(n41036), .B2(n39911), .C1(
        n433), .C2(n39905), .ZN(n7705) );
  OAI222_X1 U32383 ( .A1(n40658), .A2(n39918), .B1(n41042), .B2(n39911), .C1(
        n432), .C2(n39905), .ZN(n7704) );
  OAI222_X1 U32384 ( .A1(n40664), .A2(n39918), .B1(n41048), .B2(n39911), .C1(
        n431), .C2(n39905), .ZN(n7703) );
  OAI222_X1 U32385 ( .A1(n40670), .A2(n39918), .B1(n41054), .B2(n39911), .C1(
        n430), .C2(n39905), .ZN(n7702) );
  OAI222_X1 U32386 ( .A1(n40676), .A2(n39918), .B1(n41060), .B2(n39911), .C1(
        n429), .C2(n39904), .ZN(n7701) );
  OAI222_X1 U32387 ( .A1(n40682), .A2(n39918), .B1(n41066), .B2(n39911), .C1(
        n428), .C2(n39904), .ZN(n7700) );
  OAI222_X1 U32388 ( .A1(n40688), .A2(n39918), .B1(n41072), .B2(n39911), .C1(
        n427), .C2(n39904), .ZN(n7699) );
  OAI222_X1 U32389 ( .A1(n40694), .A2(n39917), .B1(n41078), .B2(n39910), .C1(
        n426), .C2(n39904), .ZN(n7698) );
  OAI222_X1 U32390 ( .A1(n40700), .A2(n39917), .B1(n41084), .B2(n39910), .C1(
        n425), .C2(n39904), .ZN(n7697) );
  OAI222_X1 U32391 ( .A1(n40706), .A2(n39917), .B1(n41090), .B2(n39910), .C1(
        n424), .C2(n39904), .ZN(n7696) );
  OAI222_X1 U32392 ( .A1(n40712), .A2(n39917), .B1(n41096), .B2(n39910), .C1(
        n423), .C2(n39904), .ZN(n7695) );
  OAI222_X1 U32393 ( .A1(n40718), .A2(n39917), .B1(n41102), .B2(n39910), .C1(
        n422), .C2(n39904), .ZN(n7694) );
  OAI222_X1 U32394 ( .A1(n40724), .A2(n39917), .B1(n41108), .B2(n39910), .C1(
        n421), .C2(n39904), .ZN(n7693) );
  OAI222_X1 U32395 ( .A1(n40730), .A2(n39917), .B1(n41114), .B2(n39910), .C1(
        n420), .C2(n39904), .ZN(n7692) );
  OAI222_X1 U32396 ( .A1(n40736), .A2(n39917), .B1(n41120), .B2(n39910), .C1(
        n419), .C2(n39904), .ZN(n7691) );
  OAI222_X1 U32397 ( .A1(n40742), .A2(n39917), .B1(n41126), .B2(n39910), .C1(
        n418), .C2(n39904), .ZN(n7690) );
  OAI222_X1 U32398 ( .A1(n40748), .A2(n39917), .B1(n41132), .B2(n39910), .C1(
        n417), .C2(n39904), .ZN(n7689) );
  OAI222_X1 U32399 ( .A1(n40754), .A2(n39917), .B1(n41138), .B2(n39910), .C1(
        n416), .C2(n39903), .ZN(n7688) );
  OAI222_X1 U32400 ( .A1(n40760), .A2(n39917), .B1(n41144), .B2(n39910), .C1(
        n415), .C2(n39903), .ZN(n7687) );
  OAI222_X1 U32401 ( .A1(n40766), .A2(n39916), .B1(n41150), .B2(n39909), .C1(
        n414), .C2(n39903), .ZN(n7686) );
  OAI222_X1 U32402 ( .A1(n40772), .A2(n39916), .B1(n41156), .B2(n39909), .C1(
        n413), .C2(n39903), .ZN(n7685) );
  OAI222_X1 U32403 ( .A1(n40778), .A2(n39916), .B1(n41162), .B2(n39909), .C1(
        n412), .C2(n39903), .ZN(n7684) );
  OAI222_X1 U32404 ( .A1(n40784), .A2(n39916), .B1(n41168), .B2(n39909), .C1(
        n411), .C2(n39903), .ZN(n7683) );
  OAI222_X1 U32405 ( .A1(n40790), .A2(n39916), .B1(n41174), .B2(n39909), .C1(
        n410), .C2(n39903), .ZN(n7682) );
  OAI222_X1 U32406 ( .A1(n40796), .A2(n39916), .B1(n41180), .B2(n39909), .C1(
        n409), .C2(n39903), .ZN(n7681) );
  OAI222_X1 U32407 ( .A1(n40802), .A2(n39916), .B1(n41186), .B2(n39909), .C1(
        n408), .C2(n39903), .ZN(n7680) );
  OAI222_X1 U32408 ( .A1(n40808), .A2(n39916), .B1(n41192), .B2(n39909), .C1(
        n407), .C2(n39903), .ZN(n7679) );
  OAI222_X1 U32409 ( .A1(n40814), .A2(n39916), .B1(n41198), .B2(n39909), .C1(
        n406), .C2(n39903), .ZN(n7678) );
  OAI222_X1 U32410 ( .A1(n40820), .A2(n39916), .B1(n41204), .B2(n39909), .C1(
        n405), .C2(n39903), .ZN(n7677) );
  OAI222_X1 U32411 ( .A1(n40826), .A2(n39916), .B1(n41210), .B2(n39909), .C1(
        n404), .C2(n39903), .ZN(n7676) );
  OAI222_X1 U32412 ( .A1(n40832), .A2(n39916), .B1(n41216), .B2(n39909), .C1(
        n403), .C2(n39902), .ZN(n7675) );
  OAI222_X1 U32413 ( .A1(n40838), .A2(n39915), .B1(n41222), .B2(n39908), .C1(
        n402), .C2(n39902), .ZN(n7674) );
  OAI222_X1 U32414 ( .A1(n40844), .A2(n39915), .B1(n41228), .B2(n39908), .C1(
        n401), .C2(n39902), .ZN(n7673) );
  OAI222_X1 U32415 ( .A1(n40850), .A2(n39915), .B1(n41234), .B2(n39908), .C1(
        n400), .C2(n39902), .ZN(n7672) );
  OAI222_X1 U32416 ( .A1(n40856), .A2(n39915), .B1(n41240), .B2(n39908), .C1(
        n399), .C2(n39902), .ZN(n7671) );
  OAI222_X1 U32417 ( .A1(n40862), .A2(n39915), .B1(n41246), .B2(n39908), .C1(
        n398), .C2(n39902), .ZN(n7670) );
  OAI222_X1 U32418 ( .A1(n40868), .A2(n39915), .B1(n41252), .B2(n39908), .C1(
        n397), .C2(n39902), .ZN(n7669) );
  OAI222_X1 U32419 ( .A1(n40874), .A2(n39915), .B1(n41258), .B2(n39908), .C1(
        n396), .C2(n39902), .ZN(n7668) );
  OAI222_X1 U32420 ( .A1(n40880), .A2(n39915), .B1(n41264), .B2(n39908), .C1(
        n395), .C2(n39902), .ZN(n7667) );
  OAI222_X1 U32421 ( .A1(n40886), .A2(n39915), .B1(n41270), .B2(n39908), .C1(
        n394), .C2(n39902), .ZN(n7666) );
  OAI222_X1 U32422 ( .A1(n40892), .A2(n39915), .B1(n41276), .B2(n39908), .C1(
        n393), .C2(n39902), .ZN(n7665) );
  OAI222_X1 U32423 ( .A1(n40898), .A2(n39915), .B1(n41282), .B2(n39908), .C1(
        n392), .C2(n39902), .ZN(n7664) );
  OAI222_X1 U32424 ( .A1(n40904), .A2(n39915), .B1(n41288), .B2(n39908), .C1(
        n391), .C2(n39902), .ZN(n7663) );
  OAI222_X1 U32425 ( .A1(n40622), .A2(n39937), .B1(n41006), .B2(n39930), .C1(
        n502), .C2(n39924), .ZN(n7774) );
  OAI222_X1 U32426 ( .A1(n40628), .A2(n39937), .B1(n41012), .B2(n39930), .C1(
        n501), .C2(n39924), .ZN(n7773) );
  OAI222_X1 U32427 ( .A1(n40634), .A2(n39937), .B1(n41018), .B2(n39930), .C1(
        n500), .C2(n39924), .ZN(n7772) );
  OAI222_X1 U32428 ( .A1(n40640), .A2(n39937), .B1(n41024), .B2(n39930), .C1(
        n499), .C2(n39924), .ZN(n7771) );
  OAI222_X1 U32429 ( .A1(n40646), .A2(n39937), .B1(n41030), .B2(n39930), .C1(
        n498), .C2(n39924), .ZN(n7770) );
  OAI222_X1 U32430 ( .A1(n40652), .A2(n39937), .B1(n41036), .B2(n39930), .C1(
        n497), .C2(n39924), .ZN(n7769) );
  OAI222_X1 U32431 ( .A1(n40658), .A2(n39937), .B1(n41042), .B2(n39930), .C1(
        n496), .C2(n39924), .ZN(n7768) );
  OAI222_X1 U32432 ( .A1(n40664), .A2(n39937), .B1(n41048), .B2(n39930), .C1(
        n495), .C2(n39924), .ZN(n7767) );
  OAI222_X1 U32433 ( .A1(n40670), .A2(n39937), .B1(n41054), .B2(n39930), .C1(
        n494), .C2(n39924), .ZN(n7766) );
  OAI222_X1 U32434 ( .A1(n40676), .A2(n39937), .B1(n41060), .B2(n39930), .C1(
        n493), .C2(n39923), .ZN(n7765) );
  OAI222_X1 U32435 ( .A1(n40682), .A2(n39937), .B1(n41066), .B2(n39930), .C1(
        n492), .C2(n39923), .ZN(n7764) );
  OAI222_X1 U32436 ( .A1(n40688), .A2(n39937), .B1(n41072), .B2(n39930), .C1(
        n491), .C2(n39923), .ZN(n7763) );
  OAI222_X1 U32437 ( .A1(n40694), .A2(n39936), .B1(n41078), .B2(n39929), .C1(
        n490), .C2(n39923), .ZN(n7762) );
  OAI222_X1 U32438 ( .A1(n40700), .A2(n39936), .B1(n41084), .B2(n39929), .C1(
        n489), .C2(n39923), .ZN(n7761) );
  OAI222_X1 U32439 ( .A1(n40706), .A2(n39936), .B1(n41090), .B2(n39929), .C1(
        n488), .C2(n39923), .ZN(n7760) );
  OAI222_X1 U32440 ( .A1(n40712), .A2(n39936), .B1(n41096), .B2(n39929), .C1(
        n487), .C2(n39923), .ZN(n7759) );
  OAI222_X1 U32441 ( .A1(n40718), .A2(n39936), .B1(n41102), .B2(n39929), .C1(
        n486), .C2(n39923), .ZN(n7758) );
  OAI222_X1 U32442 ( .A1(n40724), .A2(n39936), .B1(n41108), .B2(n39929), .C1(
        n485), .C2(n39923), .ZN(n7757) );
  OAI222_X1 U32443 ( .A1(n40730), .A2(n39936), .B1(n41114), .B2(n39929), .C1(
        n484), .C2(n39923), .ZN(n7756) );
  OAI222_X1 U32444 ( .A1(n40736), .A2(n39936), .B1(n41120), .B2(n39929), .C1(
        n483), .C2(n39923), .ZN(n7755) );
  OAI222_X1 U32445 ( .A1(n40742), .A2(n39936), .B1(n41126), .B2(n39929), .C1(
        n482), .C2(n39923), .ZN(n7754) );
  OAI222_X1 U32446 ( .A1(n40748), .A2(n39936), .B1(n41132), .B2(n39929), .C1(
        n481), .C2(n39923), .ZN(n7753) );
  OAI222_X1 U32447 ( .A1(n40754), .A2(n39936), .B1(n41138), .B2(n39929), .C1(
        n480), .C2(n39922), .ZN(n7752) );
  OAI222_X1 U32448 ( .A1(n40760), .A2(n39936), .B1(n41144), .B2(n39929), .C1(
        n479), .C2(n39922), .ZN(n7751) );
  OAI222_X1 U32449 ( .A1(n40766), .A2(n39935), .B1(n41150), .B2(n39928), .C1(
        n478), .C2(n39922), .ZN(n7750) );
  OAI222_X1 U32450 ( .A1(n40772), .A2(n39935), .B1(n41156), .B2(n39928), .C1(
        n477), .C2(n39922), .ZN(n7749) );
  OAI222_X1 U32451 ( .A1(n40778), .A2(n39935), .B1(n41162), .B2(n39928), .C1(
        n476), .C2(n39922), .ZN(n7748) );
  OAI222_X1 U32452 ( .A1(n40784), .A2(n39935), .B1(n41168), .B2(n39928), .C1(
        n475), .C2(n39922), .ZN(n7747) );
  OAI222_X1 U32453 ( .A1(n40790), .A2(n39935), .B1(n41174), .B2(n39928), .C1(
        n474), .C2(n39922), .ZN(n7746) );
  OAI222_X1 U32454 ( .A1(n40796), .A2(n39935), .B1(n41180), .B2(n39928), .C1(
        n473), .C2(n39922), .ZN(n7745) );
  OAI222_X1 U32455 ( .A1(n40802), .A2(n39935), .B1(n41186), .B2(n39928), .C1(
        n472), .C2(n39922), .ZN(n7744) );
  OAI222_X1 U32456 ( .A1(n40808), .A2(n39935), .B1(n41192), .B2(n39928), .C1(
        n471), .C2(n39922), .ZN(n7743) );
  OAI222_X1 U32457 ( .A1(n40814), .A2(n39935), .B1(n41198), .B2(n39928), .C1(
        n470), .C2(n39922), .ZN(n7742) );
  OAI222_X1 U32458 ( .A1(n40820), .A2(n39935), .B1(n41204), .B2(n39928), .C1(
        n469), .C2(n39922), .ZN(n7741) );
  OAI222_X1 U32459 ( .A1(n40826), .A2(n39935), .B1(n41210), .B2(n39928), .C1(
        n468), .C2(n39922), .ZN(n7740) );
  OAI222_X1 U32460 ( .A1(n40832), .A2(n39935), .B1(n41216), .B2(n39928), .C1(
        n467), .C2(n39921), .ZN(n7739) );
  OAI222_X1 U32461 ( .A1(n40838), .A2(n39934), .B1(n41222), .B2(n39927), .C1(
        n466), .C2(n39921), .ZN(n7738) );
  OAI222_X1 U32462 ( .A1(n40844), .A2(n39934), .B1(n41228), .B2(n39927), .C1(
        n465), .C2(n39921), .ZN(n7737) );
  OAI222_X1 U32463 ( .A1(n40850), .A2(n39934), .B1(n41234), .B2(n39927), .C1(
        n464), .C2(n39921), .ZN(n7736) );
  OAI222_X1 U32464 ( .A1(n40856), .A2(n39934), .B1(n41240), .B2(n39927), .C1(
        n463), .C2(n39921), .ZN(n7735) );
  OAI222_X1 U32465 ( .A1(n40862), .A2(n39934), .B1(n41246), .B2(n39927), .C1(
        n462), .C2(n39921), .ZN(n7734) );
  OAI222_X1 U32466 ( .A1(n40868), .A2(n39934), .B1(n41252), .B2(n39927), .C1(
        n461), .C2(n39921), .ZN(n7733) );
  OAI222_X1 U32467 ( .A1(n40874), .A2(n39934), .B1(n41258), .B2(n39927), .C1(
        n460), .C2(n39921), .ZN(n7732) );
  OAI222_X1 U32468 ( .A1(n40880), .A2(n39934), .B1(n41264), .B2(n39927), .C1(
        n459), .C2(n39921), .ZN(n7731) );
  OAI222_X1 U32469 ( .A1(n40886), .A2(n39934), .B1(n41270), .B2(n39927), .C1(
        n458), .C2(n39921), .ZN(n7730) );
  OAI222_X1 U32470 ( .A1(n40892), .A2(n39934), .B1(n41276), .B2(n39927), .C1(
        n457), .C2(n39921), .ZN(n7729) );
  OAI222_X1 U32471 ( .A1(n40898), .A2(n39934), .B1(n41282), .B2(n39927), .C1(
        n456), .C2(n39921), .ZN(n7728) );
  OAI222_X1 U32472 ( .A1(n40904), .A2(n39934), .B1(n41288), .B2(n39927), .C1(
        n455), .C2(n39921), .ZN(n7727) );
  OAI222_X1 U32473 ( .A1(n40910), .A2(n40012), .B1(n41294), .B2(n40005), .C1(
        n710), .C2(n39999), .ZN(n7982) );
  OAI222_X1 U32474 ( .A1(n40916), .A2(n40012), .B1(n41300), .B2(n40005), .C1(
        n709), .C2(n39999), .ZN(n7981) );
  OAI222_X1 U32475 ( .A1(n40922), .A2(n40012), .B1(n41306), .B2(n40005), .C1(
        n708), .C2(n39999), .ZN(n7980) );
  OAI222_X1 U32476 ( .A1(n40928), .A2(n40012), .B1(n41312), .B2(n40005), .C1(
        n707), .C2(n39999), .ZN(n7979) );
  OAI222_X1 U32477 ( .A1(n40934), .A2(n40012), .B1(n41318), .B2(n40005), .C1(
        n706), .C2(n39999), .ZN(n7978) );
  OAI222_X1 U32478 ( .A1(n40940), .A2(n40012), .B1(n41324), .B2(n40005), .C1(
        n705), .C2(n39999), .ZN(n7977) );
  OAI222_X1 U32479 ( .A1(n40946), .A2(n40012), .B1(n41330), .B2(n40005), .C1(
        n704), .C2(n39999), .ZN(n7976) );
  OAI222_X1 U32480 ( .A1(n40952), .A2(n40012), .B1(n41336), .B2(n40005), .C1(
        n703), .C2(n39999), .ZN(n7975) );
  OAI222_X1 U32481 ( .A1(n40958), .A2(n40012), .B1(n41342), .B2(n40005), .C1(
        n702), .C2(n39999), .ZN(n7974) );
  OAI222_X1 U32482 ( .A1(n40964), .A2(n40012), .B1(n41348), .B2(n40005), .C1(
        n701), .C2(n39999), .ZN(n7973) );
  OAI222_X1 U32483 ( .A1(n40970), .A2(n40012), .B1(n41354), .B2(n40005), .C1(
        n700), .C2(n39999), .ZN(n7972) );
  OAI222_X1 U32484 ( .A1(n40976), .A2(n40012), .B1(n41360), .B2(n40005), .C1(
        n699), .C2(n39999), .ZN(n7971) );
  OAI222_X1 U32485 ( .A1(n40910), .A2(n40031), .B1(n41294), .B2(n40024), .C1(
        n774), .C2(n40018), .ZN(n8046) );
  OAI222_X1 U32486 ( .A1(n40916), .A2(n40031), .B1(n41300), .B2(n40024), .C1(
        n773), .C2(n40018), .ZN(n8045) );
  OAI222_X1 U32487 ( .A1(n40922), .A2(n40031), .B1(n41306), .B2(n40024), .C1(
        n772), .C2(n40018), .ZN(n8044) );
  OAI222_X1 U32488 ( .A1(n40928), .A2(n40031), .B1(n41312), .B2(n40024), .C1(
        n771), .C2(n40018), .ZN(n8043) );
  OAI222_X1 U32489 ( .A1(n40934), .A2(n40031), .B1(n41318), .B2(n40024), .C1(
        n770), .C2(n40018), .ZN(n8042) );
  OAI222_X1 U32490 ( .A1(n40940), .A2(n40031), .B1(n41324), .B2(n40024), .C1(
        n769), .C2(n40018), .ZN(n8041) );
  OAI222_X1 U32491 ( .A1(n40946), .A2(n40031), .B1(n41330), .B2(n40024), .C1(
        n768), .C2(n40018), .ZN(n8040) );
  OAI222_X1 U32492 ( .A1(n40952), .A2(n40031), .B1(n41336), .B2(n40024), .C1(
        n767), .C2(n40018), .ZN(n8039) );
  OAI222_X1 U32493 ( .A1(n40958), .A2(n40031), .B1(n41342), .B2(n40024), .C1(
        n766), .C2(n40018), .ZN(n8038) );
  OAI222_X1 U32494 ( .A1(n40964), .A2(n40031), .B1(n41348), .B2(n40024), .C1(
        n765), .C2(n40018), .ZN(n8037) );
  OAI222_X1 U32495 ( .A1(n40970), .A2(n40031), .B1(n41354), .B2(n40024), .C1(
        n764), .C2(n40018), .ZN(n8036) );
  OAI222_X1 U32496 ( .A1(n40976), .A2(n40031), .B1(n41360), .B2(n40024), .C1(
        n763), .C2(n40018), .ZN(n8035) );
  OAI222_X1 U32497 ( .A1(n40622), .A2(n40016), .B1(n41006), .B2(n40009), .C1(
        n758), .C2(n40003), .ZN(n8030) );
  OAI222_X1 U32498 ( .A1(n40628), .A2(n40016), .B1(n41012), .B2(n40009), .C1(
        n757), .C2(n40003), .ZN(n8029) );
  OAI222_X1 U32499 ( .A1(n40634), .A2(n40016), .B1(n41018), .B2(n40009), .C1(
        n756), .C2(n40003), .ZN(n8028) );
  OAI222_X1 U32500 ( .A1(n40640), .A2(n40016), .B1(n41024), .B2(n40009), .C1(
        n755), .C2(n40003), .ZN(n8027) );
  OAI222_X1 U32501 ( .A1(n40646), .A2(n40016), .B1(n41030), .B2(n40009), .C1(
        n754), .C2(n40003), .ZN(n8026) );
  OAI222_X1 U32502 ( .A1(n40652), .A2(n40016), .B1(n41036), .B2(n40009), .C1(
        n753), .C2(n40003), .ZN(n8025) );
  OAI222_X1 U32503 ( .A1(n40658), .A2(n40016), .B1(n41042), .B2(n40009), .C1(
        n752), .C2(n40003), .ZN(n8024) );
  OAI222_X1 U32504 ( .A1(n40664), .A2(n40016), .B1(n41048), .B2(n40009), .C1(
        n751), .C2(n40003), .ZN(n8023) );
  OAI222_X1 U32505 ( .A1(n40670), .A2(n40016), .B1(n41054), .B2(n40009), .C1(
        n750), .C2(n40003), .ZN(n8022) );
  OAI222_X1 U32506 ( .A1(n40676), .A2(n40016), .B1(n41060), .B2(n40009), .C1(
        n749), .C2(n40002), .ZN(n8021) );
  OAI222_X1 U32507 ( .A1(n40682), .A2(n40016), .B1(n41066), .B2(n40009), .C1(
        n748), .C2(n40002), .ZN(n8020) );
  OAI222_X1 U32508 ( .A1(n40688), .A2(n40016), .B1(n41072), .B2(n40009), .C1(
        n747), .C2(n40002), .ZN(n8019) );
  OAI222_X1 U32509 ( .A1(n40694), .A2(n40015), .B1(n41078), .B2(n40008), .C1(
        n746), .C2(n40002), .ZN(n8018) );
  OAI222_X1 U32510 ( .A1(n40700), .A2(n40015), .B1(n41084), .B2(n40008), .C1(
        n745), .C2(n40002), .ZN(n8017) );
  OAI222_X1 U32511 ( .A1(n40706), .A2(n40015), .B1(n41090), .B2(n40008), .C1(
        n744), .C2(n40002), .ZN(n8016) );
  OAI222_X1 U32512 ( .A1(n40712), .A2(n40015), .B1(n41096), .B2(n40008), .C1(
        n743), .C2(n40002), .ZN(n8015) );
  OAI222_X1 U32513 ( .A1(n40718), .A2(n40015), .B1(n41102), .B2(n40008), .C1(
        n742), .C2(n40002), .ZN(n8014) );
  OAI222_X1 U32514 ( .A1(n40724), .A2(n40015), .B1(n41108), .B2(n40008), .C1(
        n741), .C2(n40002), .ZN(n8013) );
  OAI222_X1 U32515 ( .A1(n40730), .A2(n40015), .B1(n41114), .B2(n40008), .C1(
        n740), .C2(n40002), .ZN(n8012) );
  OAI222_X1 U32516 ( .A1(n40736), .A2(n40015), .B1(n41120), .B2(n40008), .C1(
        n739), .C2(n40002), .ZN(n8011) );
  OAI222_X1 U32517 ( .A1(n40742), .A2(n40015), .B1(n41126), .B2(n40008), .C1(
        n738), .C2(n40002), .ZN(n8010) );
  OAI222_X1 U32518 ( .A1(n40748), .A2(n40015), .B1(n41132), .B2(n40008), .C1(
        n737), .C2(n40002), .ZN(n8009) );
  OAI222_X1 U32519 ( .A1(n40754), .A2(n40015), .B1(n41138), .B2(n40008), .C1(
        n736), .C2(n40001), .ZN(n8008) );
  OAI222_X1 U32520 ( .A1(n40760), .A2(n40015), .B1(n41144), .B2(n40008), .C1(
        n735), .C2(n40001), .ZN(n8007) );
  OAI222_X1 U32521 ( .A1(n40766), .A2(n40014), .B1(n41150), .B2(n40007), .C1(
        n734), .C2(n40001), .ZN(n8006) );
  OAI222_X1 U32522 ( .A1(n40772), .A2(n40014), .B1(n41156), .B2(n40007), .C1(
        n733), .C2(n40001), .ZN(n8005) );
  OAI222_X1 U32523 ( .A1(n40778), .A2(n40014), .B1(n41162), .B2(n40007), .C1(
        n732), .C2(n40001), .ZN(n8004) );
  OAI222_X1 U32524 ( .A1(n40784), .A2(n40014), .B1(n41168), .B2(n40007), .C1(
        n731), .C2(n40001), .ZN(n8003) );
  OAI222_X1 U32525 ( .A1(n40790), .A2(n40014), .B1(n41174), .B2(n40007), .C1(
        n730), .C2(n40001), .ZN(n8002) );
  OAI222_X1 U32526 ( .A1(n40796), .A2(n40014), .B1(n41180), .B2(n40007), .C1(
        n729), .C2(n40001), .ZN(n8001) );
  OAI222_X1 U32527 ( .A1(n40802), .A2(n40014), .B1(n41186), .B2(n40007), .C1(
        n728), .C2(n40001), .ZN(n8000) );
  OAI222_X1 U32528 ( .A1(n40808), .A2(n40014), .B1(n41192), .B2(n40007), .C1(
        n727), .C2(n40001), .ZN(n7999) );
  OAI222_X1 U32529 ( .A1(n40814), .A2(n40014), .B1(n41198), .B2(n40007), .C1(
        n726), .C2(n40001), .ZN(n7998) );
  OAI222_X1 U32530 ( .A1(n40820), .A2(n40014), .B1(n41204), .B2(n40007), .C1(
        n725), .C2(n40001), .ZN(n7997) );
  OAI222_X1 U32531 ( .A1(n40826), .A2(n40014), .B1(n41210), .B2(n40007), .C1(
        n724), .C2(n40001), .ZN(n7996) );
  OAI222_X1 U32532 ( .A1(n40832), .A2(n40014), .B1(n41216), .B2(n40007), .C1(
        n723), .C2(n40000), .ZN(n7995) );
  OAI222_X1 U32533 ( .A1(n40838), .A2(n40013), .B1(n41222), .B2(n40006), .C1(
        n722), .C2(n40000), .ZN(n7994) );
  OAI222_X1 U32534 ( .A1(n40844), .A2(n40013), .B1(n41228), .B2(n40006), .C1(
        n721), .C2(n40000), .ZN(n7993) );
  OAI222_X1 U32535 ( .A1(n40850), .A2(n40013), .B1(n41234), .B2(n40006), .C1(
        n720), .C2(n40000), .ZN(n7992) );
  OAI222_X1 U32536 ( .A1(n40856), .A2(n40013), .B1(n41240), .B2(n40006), .C1(
        n719), .C2(n40000), .ZN(n7991) );
  OAI222_X1 U32537 ( .A1(n40862), .A2(n40013), .B1(n41246), .B2(n40006), .C1(
        n718), .C2(n40000), .ZN(n7990) );
  OAI222_X1 U32538 ( .A1(n40868), .A2(n40013), .B1(n41252), .B2(n40006), .C1(
        n717), .C2(n40000), .ZN(n7989) );
  OAI222_X1 U32539 ( .A1(n40874), .A2(n40013), .B1(n41258), .B2(n40006), .C1(
        n716), .C2(n40000), .ZN(n7988) );
  OAI222_X1 U32540 ( .A1(n40880), .A2(n40013), .B1(n41264), .B2(n40006), .C1(
        n715), .C2(n40000), .ZN(n7987) );
  OAI222_X1 U32541 ( .A1(n40886), .A2(n40013), .B1(n41270), .B2(n40006), .C1(
        n714), .C2(n40000), .ZN(n7986) );
  OAI222_X1 U32542 ( .A1(n40892), .A2(n40013), .B1(n41276), .B2(n40006), .C1(
        n713), .C2(n40000), .ZN(n7985) );
  OAI222_X1 U32543 ( .A1(n40898), .A2(n40013), .B1(n41282), .B2(n40006), .C1(
        n712), .C2(n40000), .ZN(n7984) );
  OAI222_X1 U32544 ( .A1(n40904), .A2(n40013), .B1(n41288), .B2(n40006), .C1(
        n711), .C2(n40000), .ZN(n7983) );
  OAI222_X1 U32545 ( .A1(n40622), .A2(n40035), .B1(n41006), .B2(n40028), .C1(
        n822), .C2(n40022), .ZN(n8094) );
  OAI222_X1 U32546 ( .A1(n40628), .A2(n40035), .B1(n41012), .B2(n40028), .C1(
        n821), .C2(n40022), .ZN(n8093) );
  OAI222_X1 U32547 ( .A1(n40634), .A2(n40035), .B1(n41018), .B2(n40028), .C1(
        n820), .C2(n40022), .ZN(n8092) );
  OAI222_X1 U32548 ( .A1(n40640), .A2(n40035), .B1(n41024), .B2(n40028), .C1(
        n819), .C2(n40022), .ZN(n8091) );
  OAI222_X1 U32549 ( .A1(n40646), .A2(n40035), .B1(n41030), .B2(n40028), .C1(
        n818), .C2(n40022), .ZN(n8090) );
  OAI222_X1 U32550 ( .A1(n40652), .A2(n40035), .B1(n41036), .B2(n40028), .C1(
        n817), .C2(n40022), .ZN(n8089) );
  OAI222_X1 U32551 ( .A1(n40658), .A2(n40035), .B1(n41042), .B2(n40028), .C1(
        n816), .C2(n40022), .ZN(n8088) );
  OAI222_X1 U32552 ( .A1(n40664), .A2(n40035), .B1(n41048), .B2(n40028), .C1(
        n815), .C2(n40022), .ZN(n8087) );
  OAI222_X1 U32553 ( .A1(n40670), .A2(n40035), .B1(n41054), .B2(n40028), .C1(
        n814), .C2(n40022), .ZN(n8086) );
  OAI222_X1 U32554 ( .A1(n40676), .A2(n40035), .B1(n41060), .B2(n40028), .C1(
        n813), .C2(n40021), .ZN(n8085) );
  OAI222_X1 U32555 ( .A1(n40682), .A2(n40035), .B1(n41066), .B2(n40028), .C1(
        n812), .C2(n40021), .ZN(n8084) );
  OAI222_X1 U32556 ( .A1(n40688), .A2(n40035), .B1(n41072), .B2(n40028), .C1(
        n811), .C2(n40021), .ZN(n8083) );
  OAI222_X1 U32557 ( .A1(n40694), .A2(n40034), .B1(n41078), .B2(n40027), .C1(
        n810), .C2(n40021), .ZN(n8082) );
  OAI222_X1 U32558 ( .A1(n40700), .A2(n40034), .B1(n41084), .B2(n40027), .C1(
        n809), .C2(n40021), .ZN(n8081) );
  OAI222_X1 U32559 ( .A1(n40706), .A2(n40034), .B1(n41090), .B2(n40027), .C1(
        n808), .C2(n40021), .ZN(n8080) );
  OAI222_X1 U32560 ( .A1(n40712), .A2(n40034), .B1(n41096), .B2(n40027), .C1(
        n807), .C2(n40021), .ZN(n8079) );
  OAI222_X1 U32561 ( .A1(n40718), .A2(n40034), .B1(n41102), .B2(n40027), .C1(
        n806), .C2(n40021), .ZN(n8078) );
  OAI222_X1 U32562 ( .A1(n40724), .A2(n40034), .B1(n41108), .B2(n40027), .C1(
        n805), .C2(n40021), .ZN(n8077) );
  OAI222_X1 U32563 ( .A1(n40730), .A2(n40034), .B1(n41114), .B2(n40027), .C1(
        n804), .C2(n40021), .ZN(n8076) );
  OAI222_X1 U32564 ( .A1(n40736), .A2(n40034), .B1(n41120), .B2(n40027), .C1(
        n803), .C2(n40021), .ZN(n8075) );
  OAI222_X1 U32565 ( .A1(n40742), .A2(n40034), .B1(n41126), .B2(n40027), .C1(
        n802), .C2(n40021), .ZN(n8074) );
  OAI222_X1 U32566 ( .A1(n40748), .A2(n40034), .B1(n41132), .B2(n40027), .C1(
        n801), .C2(n40021), .ZN(n8073) );
  OAI222_X1 U32567 ( .A1(n40754), .A2(n40034), .B1(n41138), .B2(n40027), .C1(
        n800), .C2(n40020), .ZN(n8072) );
  OAI222_X1 U32568 ( .A1(n40760), .A2(n40034), .B1(n41144), .B2(n40027), .C1(
        n799), .C2(n40020), .ZN(n8071) );
  OAI222_X1 U32569 ( .A1(n40766), .A2(n40033), .B1(n41150), .B2(n40026), .C1(
        n798), .C2(n40020), .ZN(n8070) );
  OAI222_X1 U32570 ( .A1(n40772), .A2(n40033), .B1(n41156), .B2(n40026), .C1(
        n797), .C2(n40020), .ZN(n8069) );
  OAI222_X1 U32571 ( .A1(n40778), .A2(n40033), .B1(n41162), .B2(n40026), .C1(
        n796), .C2(n40020), .ZN(n8068) );
  OAI222_X1 U32572 ( .A1(n40784), .A2(n40033), .B1(n41168), .B2(n40026), .C1(
        n795), .C2(n40020), .ZN(n8067) );
  OAI222_X1 U32573 ( .A1(n40790), .A2(n40033), .B1(n41174), .B2(n40026), .C1(
        n794), .C2(n40020), .ZN(n8066) );
  OAI222_X1 U32574 ( .A1(n40796), .A2(n40033), .B1(n41180), .B2(n40026), .C1(
        n793), .C2(n40020), .ZN(n8065) );
  OAI222_X1 U32575 ( .A1(n40802), .A2(n40033), .B1(n41186), .B2(n40026), .C1(
        n792), .C2(n40020), .ZN(n8064) );
  OAI222_X1 U32576 ( .A1(n40808), .A2(n40033), .B1(n41192), .B2(n40026), .C1(
        n791), .C2(n40020), .ZN(n8063) );
  OAI222_X1 U32577 ( .A1(n40814), .A2(n40033), .B1(n41198), .B2(n40026), .C1(
        n790), .C2(n40020), .ZN(n8062) );
  OAI222_X1 U32578 ( .A1(n40820), .A2(n40033), .B1(n41204), .B2(n40026), .C1(
        n789), .C2(n40020), .ZN(n8061) );
  OAI222_X1 U32579 ( .A1(n40826), .A2(n40033), .B1(n41210), .B2(n40026), .C1(
        n788), .C2(n40020), .ZN(n8060) );
  OAI222_X1 U32580 ( .A1(n40832), .A2(n40033), .B1(n41216), .B2(n40026), .C1(
        n787), .C2(n40019), .ZN(n8059) );
  OAI222_X1 U32581 ( .A1(n40838), .A2(n40032), .B1(n41222), .B2(n40025), .C1(
        n786), .C2(n40019), .ZN(n8058) );
  OAI222_X1 U32582 ( .A1(n40844), .A2(n40032), .B1(n41228), .B2(n40025), .C1(
        n785), .C2(n40019), .ZN(n8057) );
  OAI222_X1 U32583 ( .A1(n40850), .A2(n40032), .B1(n41234), .B2(n40025), .C1(
        n784), .C2(n40019), .ZN(n8056) );
  OAI222_X1 U32584 ( .A1(n40856), .A2(n40032), .B1(n41240), .B2(n40025), .C1(
        n783), .C2(n40019), .ZN(n8055) );
  OAI222_X1 U32585 ( .A1(n40862), .A2(n40032), .B1(n41246), .B2(n40025), .C1(
        n782), .C2(n40019), .ZN(n8054) );
  OAI222_X1 U32586 ( .A1(n40868), .A2(n40032), .B1(n41252), .B2(n40025), .C1(
        n781), .C2(n40019), .ZN(n8053) );
  OAI222_X1 U32587 ( .A1(n40874), .A2(n40032), .B1(n41258), .B2(n40025), .C1(
        n780), .C2(n40019), .ZN(n8052) );
  OAI222_X1 U32588 ( .A1(n40880), .A2(n40032), .B1(n41264), .B2(n40025), .C1(
        n779), .C2(n40019), .ZN(n8051) );
  OAI222_X1 U32589 ( .A1(n40886), .A2(n40032), .B1(n41270), .B2(n40025), .C1(
        n778), .C2(n40019), .ZN(n8050) );
  OAI222_X1 U32590 ( .A1(n40892), .A2(n40032), .B1(n41276), .B2(n40025), .C1(
        n777), .C2(n40019), .ZN(n8049) );
  OAI222_X1 U32591 ( .A1(n40898), .A2(n40032), .B1(n41282), .B2(n40025), .C1(
        n776), .C2(n40019), .ZN(n8048) );
  OAI222_X1 U32592 ( .A1(n40904), .A2(n40032), .B1(n41288), .B2(n40025), .C1(
        n775), .C2(n40019), .ZN(n8047) );
  OAI222_X1 U32593 ( .A1(n40736), .A2(n39818), .B1(n41120), .B2(n39811), .C1(
        n99), .C2(n39805), .ZN(n7371) );
  OAI222_X1 U32594 ( .A1(n40742), .A2(n39818), .B1(n41126), .B2(n39811), .C1(
        n98), .C2(n39805), .ZN(n7370) );
  OAI222_X1 U32595 ( .A1(n40748), .A2(n39818), .B1(n41132), .B2(n39811), .C1(
        n97), .C2(n39805), .ZN(n7369) );
  OAI222_X1 U32596 ( .A1(n40754), .A2(n39818), .B1(n41138), .B2(n39811), .C1(
        n96), .C2(n39804), .ZN(n7368) );
  OAI222_X1 U32597 ( .A1(n40760), .A2(n39818), .B1(n41144), .B2(n39811), .C1(
        n95), .C2(n39804), .ZN(n7367) );
  OAI222_X1 U32598 ( .A1(n40766), .A2(n39817), .B1(n41150), .B2(n39810), .C1(
        n94), .C2(n39804), .ZN(n7366) );
  OAI222_X1 U32599 ( .A1(n40772), .A2(n39817), .B1(n41156), .B2(n39810), .C1(
        n93), .C2(n39804), .ZN(n7365) );
  OAI222_X1 U32600 ( .A1(n40778), .A2(n39817), .B1(n41162), .B2(n39810), .C1(
        n92), .C2(n39804), .ZN(n7364) );
  OAI222_X1 U32601 ( .A1(n40784), .A2(n39817), .B1(n41168), .B2(n39810), .C1(
        n91), .C2(n39804), .ZN(n7363) );
  OAI222_X1 U32602 ( .A1(n40790), .A2(n39817), .B1(n41174), .B2(n39810), .C1(
        n90), .C2(n39804), .ZN(n7362) );
  OAI222_X1 U32603 ( .A1(n40796), .A2(n39817), .B1(n41180), .B2(n39810), .C1(
        n89), .C2(n39804), .ZN(n7361) );
  OAI222_X1 U32604 ( .A1(n40802), .A2(n39817), .B1(n41186), .B2(n39810), .C1(
        n88), .C2(n39804), .ZN(n7360) );
  OAI222_X1 U32605 ( .A1(n40808), .A2(n39817), .B1(n41192), .B2(n39810), .C1(
        n87), .C2(n39804), .ZN(n7359) );
  OAI222_X1 U32606 ( .A1(n40814), .A2(n39817), .B1(n41198), .B2(n39810), .C1(
        n86), .C2(n39804), .ZN(n7358) );
  OAI222_X1 U32607 ( .A1(n40820), .A2(n39817), .B1(n41204), .B2(n39810), .C1(
        n85), .C2(n39804), .ZN(n7357) );
  OAI222_X1 U32608 ( .A1(n40826), .A2(n39817), .B1(n41210), .B2(n39810), .C1(
        n84), .C2(n39804), .ZN(n7356) );
  OAI222_X1 U32609 ( .A1(n40832), .A2(n39817), .B1(n41216), .B2(n39810), .C1(
        n83), .C2(n39803), .ZN(n7355) );
  OAI222_X1 U32610 ( .A1(n40838), .A2(n39816), .B1(n41222), .B2(n39809), .C1(
        n82), .C2(n39803), .ZN(n7354) );
  OAI222_X1 U32611 ( .A1(n40844), .A2(n39816), .B1(n41228), .B2(n39809), .C1(
        n81), .C2(n39803), .ZN(n7353) );
  OAI222_X1 U32612 ( .A1(n40850), .A2(n39816), .B1(n41234), .B2(n39809), .C1(
        n80), .C2(n39803), .ZN(n7352) );
  OAI222_X1 U32613 ( .A1(n40856), .A2(n39816), .B1(n41240), .B2(n39809), .C1(
        n79), .C2(n39803), .ZN(n7351) );
  OAI222_X1 U32614 ( .A1(n40862), .A2(n39816), .B1(n41246), .B2(n39809), .C1(
        n78), .C2(n39803), .ZN(n7350) );
  OAI222_X1 U32615 ( .A1(n40868), .A2(n39816), .B1(n41252), .B2(n39809), .C1(
        n77), .C2(n39803), .ZN(n7349) );
  OAI222_X1 U32616 ( .A1(n40874), .A2(n39816), .B1(n41258), .B2(n39809), .C1(
        n76), .C2(n39803), .ZN(n7348) );
  OAI222_X1 U32617 ( .A1(n40880), .A2(n39816), .B1(n41264), .B2(n39809), .C1(
        n75), .C2(n39803), .ZN(n7347) );
  OAI222_X1 U32618 ( .A1(n40886), .A2(n39816), .B1(n41270), .B2(n39809), .C1(
        n74), .C2(n39803), .ZN(n7346) );
  OAI222_X1 U32619 ( .A1(n40892), .A2(n39816), .B1(n41276), .B2(n39809), .C1(
        n73), .C2(n39803), .ZN(n7345) );
  OAI222_X1 U32620 ( .A1(n40898), .A2(n39816), .B1(n41282), .B2(n39809), .C1(
        n72), .C2(n39803), .ZN(n7344) );
  OAI222_X1 U32621 ( .A1(n40904), .A2(n39816), .B1(n41288), .B2(n39809), .C1(
        n71), .C2(n39803), .ZN(n7343) );
  OAI222_X1 U32622 ( .A1(n40910), .A2(n39815), .B1(n41294), .B2(n39808), .C1(
        n70), .C2(n39802), .ZN(n7342) );
  OAI222_X1 U32623 ( .A1(n40916), .A2(n39815), .B1(n41300), .B2(n39808), .C1(
        n69), .C2(n39802), .ZN(n7341) );
  OAI222_X1 U32624 ( .A1(n40922), .A2(n39815), .B1(n41306), .B2(n39808), .C1(
        n68), .C2(n39802), .ZN(n7340) );
  OAI222_X1 U32625 ( .A1(n40928), .A2(n39815), .B1(n41312), .B2(n39808), .C1(
        n67), .C2(n39802), .ZN(n7339) );
  OAI222_X1 U32626 ( .A1(n40934), .A2(n39815), .B1(n41318), .B2(n39808), .C1(
        n66), .C2(n39802), .ZN(n7338) );
  OAI222_X1 U32627 ( .A1(n40940), .A2(n39815), .B1(n41324), .B2(n39808), .C1(
        n65), .C2(n39802), .ZN(n7337) );
  OAI222_X1 U32628 ( .A1(n40946), .A2(n39815), .B1(n41330), .B2(n39808), .C1(
        n64), .C2(n39802), .ZN(n7336) );
  OAI222_X1 U32629 ( .A1(n40952), .A2(n39815), .B1(n41336), .B2(n39808), .C1(
        n63), .C2(n39802), .ZN(n7335) );
  OAI222_X1 U32630 ( .A1(n40970), .A2(n39815), .B1(n41354), .B2(n39808), .C1(
        n60), .C2(n39802), .ZN(n7332) );
  OAI222_X1 U32631 ( .A1(n40976), .A2(n39815), .B1(n41360), .B2(n39808), .C1(
        n59), .C2(n39802), .ZN(n7331) );
  OAI222_X1 U32632 ( .A1(n40958), .A2(n39815), .B1(n41342), .B2(n39808), .C1(
        n62), .C2(n39802), .ZN(n7334) );
  OAI222_X1 U32633 ( .A1(n40964), .A2(n39815), .B1(n41348), .B2(n39808), .C1(
        n61), .C2(n39802), .ZN(n7333) );
  OAI222_X1 U32634 ( .A1(n40598), .A2(n39919), .B1(n40982), .B2(n39912), .C1(
        n442), .C2(n39905), .ZN(n7714) );
  OAI222_X1 U32635 ( .A1(n40604), .A2(n39919), .B1(n40988), .B2(n39912), .C1(
        n441), .C2(n39905), .ZN(n7713) );
  OAI222_X1 U32636 ( .A1(n40610), .A2(n39919), .B1(n40994), .B2(n39912), .C1(
        n440), .C2(n39905), .ZN(n7712) );
  OAI222_X1 U32637 ( .A1(n40616), .A2(n39919), .B1(n41000), .B2(n39912), .C1(
        n439), .C2(n39905), .ZN(n7711) );
  OAI222_X1 U32638 ( .A1(n40598), .A2(n39938), .B1(n40982), .B2(n39931), .C1(
        n506), .C2(n39924), .ZN(n7778) );
  OAI222_X1 U32639 ( .A1(n40604), .A2(n39938), .B1(n40988), .B2(n39931), .C1(
        n505), .C2(n39924), .ZN(n7777) );
  OAI222_X1 U32640 ( .A1(n40610), .A2(n39938), .B1(n40994), .B2(n39931), .C1(
        n504), .C2(n39924), .ZN(n7776) );
  OAI222_X1 U32641 ( .A1(n40616), .A2(n39938), .B1(n41000), .B2(n39931), .C1(
        n503), .C2(n39924), .ZN(n7775) );
  OAI222_X1 U32642 ( .A1(n40598), .A2(n40017), .B1(n40982), .B2(n40010), .C1(
        n762), .C2(n40003), .ZN(n8034) );
  OAI222_X1 U32643 ( .A1(n40604), .A2(n40017), .B1(n40988), .B2(n40010), .C1(
        n761), .C2(n40003), .ZN(n8033) );
  OAI222_X1 U32644 ( .A1(n40610), .A2(n40017), .B1(n40994), .B2(n40010), .C1(
        n760), .C2(n40003), .ZN(n8032) );
  OAI222_X1 U32645 ( .A1(n40616), .A2(n40017), .B1(n41000), .B2(n40010), .C1(
        n759), .C2(n40003), .ZN(n8031) );
  OAI222_X1 U32646 ( .A1(n40598), .A2(n40036), .B1(n40982), .B2(n40029), .C1(
        n826), .C2(n40022), .ZN(n8098) );
  OAI222_X1 U32647 ( .A1(n40604), .A2(n40036), .B1(n40988), .B2(n40029), .C1(
        n825), .C2(n40022), .ZN(n8097) );
  OAI222_X1 U32648 ( .A1(n40610), .A2(n40036), .B1(n40994), .B2(n40029), .C1(
        n824), .C2(n40022), .ZN(n8096) );
  OAI222_X1 U32649 ( .A1(n40616), .A2(n40036), .B1(n41000), .B2(n40029), .C1(
        n823), .C2(n40022), .ZN(n8095) );
  OAI222_X1 U32650 ( .A1(n40659), .A2(n40134), .B1(n41043), .B2(n40127), .C1(
        n25458), .C2(n40117), .ZN(n8408) );
  OAI222_X1 U32651 ( .A1(n40665), .A2(n40134), .B1(n41049), .B2(n40127), .C1(
        n25459), .C2(n40117), .ZN(n8407) );
  OAI222_X1 U32652 ( .A1(n40671), .A2(n40134), .B1(n41055), .B2(n40127), .C1(
        n25460), .C2(n40117), .ZN(n8406) );
  OAI222_X1 U32653 ( .A1(n40677), .A2(n40134), .B1(n41061), .B2(n40127), .C1(
        n25461), .C2(n40117), .ZN(n8405) );
  OAI222_X1 U32654 ( .A1(n40683), .A2(n40134), .B1(n41067), .B2(n40127), .C1(
        n25462), .C2(n40117), .ZN(n8404) );
  OAI222_X1 U32655 ( .A1(n40689), .A2(n40134), .B1(n41073), .B2(n40127), .C1(
        n25463), .C2(n40118), .ZN(n8403) );
  OAI222_X1 U32656 ( .A1(n40695), .A2(n40133), .B1(n41079), .B2(n40126), .C1(
        n25464), .C2(n40117), .ZN(n8402) );
  OAI222_X1 U32657 ( .A1(n40701), .A2(n40133), .B1(n41085), .B2(n40126), .C1(
        n25465), .C2(n40117), .ZN(n8401) );
  OAI222_X1 U32658 ( .A1(n40707), .A2(n40133), .B1(n41091), .B2(n40126), .C1(
        n25466), .C2(n40117), .ZN(n8400) );
  OAI222_X1 U32659 ( .A1(n40713), .A2(n40133), .B1(n41097), .B2(n40126), .C1(
        n25467), .C2(n40117), .ZN(n8399) );
  OAI222_X1 U32660 ( .A1(n40719), .A2(n40133), .B1(n41103), .B2(n40126), .C1(
        n25468), .C2(n40117), .ZN(n8398) );
  OAI222_X1 U32661 ( .A1(n40725), .A2(n40133), .B1(n41109), .B2(n40126), .C1(
        n25469), .C2(n40117), .ZN(n8397) );
  OAI222_X1 U32662 ( .A1(n40731), .A2(n40133), .B1(n41115), .B2(n40126), .C1(
        n25470), .C2(n40117), .ZN(n8396) );
  OAI222_X1 U32663 ( .A1(n40737), .A2(n40133), .B1(n41121), .B2(n40126), .C1(
        n25471), .C2(n40117), .ZN(n8395) );
  OAI222_X1 U32664 ( .A1(n40743), .A2(n40133), .B1(n41127), .B2(n40126), .C1(
        n25472), .C2(n40118), .ZN(n8394) );
  OAI222_X1 U32665 ( .A1(n40749), .A2(n40133), .B1(n41133), .B2(n40126), .C1(
        n25473), .C2(n40118), .ZN(n8393) );
  OAI222_X1 U32666 ( .A1(n40755), .A2(n40133), .B1(n41139), .B2(n40126), .C1(
        n25474), .C2(n40118), .ZN(n8392) );
  OAI222_X1 U32667 ( .A1(n40761), .A2(n40133), .B1(n41145), .B2(n40126), .C1(
        n25475), .C2(n40118), .ZN(n8391) );
  OAI222_X1 U32668 ( .A1(n40767), .A2(n40132), .B1(n41151), .B2(n40125), .C1(
        n25476), .C2(n40118), .ZN(n8390) );
  OAI222_X1 U32669 ( .A1(n40773), .A2(n40132), .B1(n41157), .B2(n40125), .C1(
        n25477), .C2(n40118), .ZN(n8389) );
  OAI222_X1 U32670 ( .A1(n40779), .A2(n40132), .B1(n41163), .B2(n40125), .C1(
        n25478), .C2(n40118), .ZN(n8388) );
  OAI222_X1 U32671 ( .A1(n40785), .A2(n40132), .B1(n41169), .B2(n40125), .C1(
        n25479), .C2(n40118), .ZN(n8387) );
  OAI222_X1 U32672 ( .A1(n40791), .A2(n40132), .B1(n41175), .B2(n40125), .C1(
        n25480), .C2(n40118), .ZN(n8386) );
  OAI222_X1 U32673 ( .A1(n40797), .A2(n40132), .B1(n41181), .B2(n40125), .C1(
        n25481), .C2(n40118), .ZN(n8385) );
  OAI222_X1 U32674 ( .A1(n40803), .A2(n40132), .B1(n41187), .B2(n40125), .C1(
        n25482), .C2(n40118), .ZN(n8384) );
  OAI222_X1 U32675 ( .A1(n40809), .A2(n40132), .B1(n41193), .B2(n40125), .C1(
        n25483), .C2(n40118), .ZN(n8383) );
  OAI222_X1 U32676 ( .A1(n40815), .A2(n40132), .B1(n41199), .B2(n40125), .C1(
        n25484), .C2(n40119), .ZN(n8382) );
  OAI222_X1 U32677 ( .A1(n40821), .A2(n40132), .B1(n41205), .B2(n40125), .C1(
        n25485), .C2(n40119), .ZN(n8381) );
  OAI222_X1 U32678 ( .A1(n40827), .A2(n40132), .B1(n41211), .B2(n40125), .C1(
        n25486), .C2(n40119), .ZN(n8380) );
  OAI222_X1 U32679 ( .A1(n40833), .A2(n40132), .B1(n41217), .B2(n40125), .C1(
        n25487), .C2(n40119), .ZN(n8379) );
  OAI222_X1 U32680 ( .A1(n40839), .A2(n40131), .B1(n41223), .B2(n40124), .C1(
        n25488), .C2(n40119), .ZN(n8378) );
  OAI222_X1 U32681 ( .A1(n40845), .A2(n40131), .B1(n41229), .B2(n40124), .C1(
        n25489), .C2(n40119), .ZN(n8377) );
  OAI222_X1 U32682 ( .A1(n40851), .A2(n40131), .B1(n41235), .B2(n40124), .C1(
        n25490), .C2(n40119), .ZN(n8376) );
  OAI222_X1 U32683 ( .A1(n40857), .A2(n40131), .B1(n41241), .B2(n40124), .C1(
        n25491), .C2(n40119), .ZN(n8375) );
  OAI222_X1 U32684 ( .A1(n40863), .A2(n40131), .B1(n41247), .B2(n40124), .C1(
        n25492), .C2(n40119), .ZN(n8374) );
  OAI222_X1 U32685 ( .A1(n40869), .A2(n40131), .B1(n41253), .B2(n40124), .C1(
        n25493), .C2(n40119), .ZN(n8373) );
  OAI222_X1 U32686 ( .A1(n40875), .A2(n40131), .B1(n41259), .B2(n40124), .C1(
        n25494), .C2(n40119), .ZN(n8372) );
  OAI222_X1 U32687 ( .A1(n40881), .A2(n40131), .B1(n41265), .B2(n40124), .C1(
        n25495), .C2(n40119), .ZN(n8371) );
  OAI222_X1 U32688 ( .A1(n40887), .A2(n40131), .B1(n41271), .B2(n40124), .C1(
        n25496), .C2(n40119), .ZN(n8370) );
  OAI222_X1 U32689 ( .A1(n40893), .A2(n40131), .B1(n41277), .B2(n40124), .C1(
        n25497), .C2(n40120), .ZN(n8369) );
  OAI222_X1 U32690 ( .A1(n40899), .A2(n40131), .B1(n41283), .B2(n40124), .C1(
        n25498), .C2(n40120), .ZN(n8368) );
  OAI222_X1 U32691 ( .A1(n40905), .A2(n40131), .B1(n41289), .B2(n40124), .C1(
        n25499), .C2(n40120), .ZN(n8367) );
  OAI222_X1 U32692 ( .A1(n40911), .A2(n40130), .B1(n41295), .B2(n40123), .C1(
        n25500), .C2(n40120), .ZN(n8366) );
  OAI222_X1 U32693 ( .A1(n40917), .A2(n40130), .B1(n41301), .B2(n40123), .C1(
        n25501), .C2(n40120), .ZN(n8365) );
  OAI222_X1 U32694 ( .A1(n40923), .A2(n40130), .B1(n41307), .B2(n40123), .C1(
        n25502), .C2(n40120), .ZN(n8364) );
  OAI222_X1 U32695 ( .A1(n40929), .A2(n40130), .B1(n41313), .B2(n40123), .C1(
        n25503), .C2(n40120), .ZN(n8363) );
  OAI222_X1 U32696 ( .A1(n40935), .A2(n40130), .B1(n41319), .B2(n40123), .C1(
        n25504), .C2(n40120), .ZN(n8362) );
  OAI222_X1 U32697 ( .A1(n40941), .A2(n40130), .B1(n41325), .B2(n40123), .C1(
        n25505), .C2(n40120), .ZN(n8361) );
  OAI222_X1 U32698 ( .A1(n40947), .A2(n40130), .B1(n41331), .B2(n40123), .C1(
        n25506), .C2(n40120), .ZN(n8360) );
  OAI222_X1 U32699 ( .A1(n40953), .A2(n40130), .B1(n41337), .B2(n40123), .C1(
        n25507), .C2(n40120), .ZN(n8359) );
  OAI222_X1 U32700 ( .A1(n40959), .A2(n40130), .B1(n41343), .B2(n40123), .C1(
        n25508), .C2(n40120), .ZN(n8358) );
  OAI222_X1 U32701 ( .A1(n40965), .A2(n40130), .B1(n41349), .B2(n40123), .C1(
        n25509), .C2(n40121), .ZN(n8357) );
  OAI222_X1 U32702 ( .A1(n40971), .A2(n40130), .B1(n41355), .B2(n40123), .C1(
        n25510), .C2(n40120), .ZN(n8356) );
  OAI222_X1 U32703 ( .A1(n40977), .A2(n40130), .B1(n41361), .B2(n40123), .C1(
        n25511), .C2(n40116), .ZN(n8355) );
  OAI222_X1 U32704 ( .A1(n40599), .A2(n40115), .B1(n40983), .B2(n40108), .C1(
        n25398), .C2(n40101), .ZN(n8354) );
  OAI222_X1 U32705 ( .A1(n40605), .A2(n40115), .B1(n40989), .B2(n40108), .C1(
        n25399), .C2(n40101), .ZN(n8353) );
  OAI222_X1 U32706 ( .A1(n40611), .A2(n40115), .B1(n40995), .B2(n40108), .C1(
        n25400), .C2(n40101), .ZN(n8352) );
  OAI222_X1 U32707 ( .A1(n40617), .A2(n40115), .B1(n41001), .B2(n40108), .C1(
        n25401), .C2(n40101), .ZN(n8351) );
  OAI222_X1 U32708 ( .A1(n40623), .A2(n40114), .B1(n41007), .B2(n40107), .C1(
        n25402), .C2(n40101), .ZN(n8350) );
  OAI222_X1 U32709 ( .A1(n40629), .A2(n40114), .B1(n41013), .B2(n40107), .C1(
        n25403), .C2(n40101), .ZN(n8349) );
  OAI222_X1 U32710 ( .A1(n40635), .A2(n40114), .B1(n41019), .B2(n40107), .C1(
        n25404), .C2(n40101), .ZN(n8348) );
  OAI222_X1 U32711 ( .A1(n40641), .A2(n40114), .B1(n41025), .B2(n40107), .C1(
        n25405), .C2(n40101), .ZN(n8347) );
  OAI222_X1 U32712 ( .A1(n40647), .A2(n40114), .B1(n41031), .B2(n40107), .C1(
        n25406), .C2(n40101), .ZN(n8346) );
  OAI222_X1 U32713 ( .A1(n40653), .A2(n40114), .B1(n41037), .B2(n40107), .C1(
        n25407), .C2(n40101), .ZN(n8345) );
  OAI222_X1 U32714 ( .A1(n40659), .A2(n40114), .B1(n41043), .B2(n40107), .C1(
        n25408), .C2(n40101), .ZN(n8344) );
  OAI222_X1 U32715 ( .A1(n40665), .A2(n40114), .B1(n41049), .B2(n40107), .C1(
        n25409), .C2(n40101), .ZN(n8343) );
  OAI222_X1 U32716 ( .A1(n40671), .A2(n40114), .B1(n41055), .B2(n40107), .C1(
        n25410), .C2(n40101), .ZN(n8342) );
  OAI222_X1 U32717 ( .A1(n40677), .A2(n40114), .B1(n41061), .B2(n40107), .C1(
        n25411), .C2(n40100), .ZN(n8341) );
  OAI222_X1 U32718 ( .A1(n40683), .A2(n40114), .B1(n41067), .B2(n40107), .C1(
        n25412), .C2(n40100), .ZN(n8340) );
  OAI222_X1 U32719 ( .A1(n40689), .A2(n40114), .B1(n41073), .B2(n40107), .C1(
        n25413), .C2(n40100), .ZN(n8339) );
  OAI222_X1 U32720 ( .A1(n40695), .A2(n40113), .B1(n41079), .B2(n40106), .C1(
        n25414), .C2(n40100), .ZN(n8338) );
  OAI222_X1 U32721 ( .A1(n40701), .A2(n40113), .B1(n41085), .B2(n40106), .C1(
        n25415), .C2(n40100), .ZN(n8337) );
  OAI222_X1 U32722 ( .A1(n40707), .A2(n40113), .B1(n41091), .B2(n40106), .C1(
        n25416), .C2(n40100), .ZN(n8336) );
  OAI222_X1 U32723 ( .A1(n40713), .A2(n40113), .B1(n41097), .B2(n40106), .C1(
        n25417), .C2(n40100), .ZN(n8335) );
  OAI222_X1 U32724 ( .A1(n40719), .A2(n40113), .B1(n41103), .B2(n40106), .C1(
        n25418), .C2(n40100), .ZN(n8334) );
  OAI222_X1 U32725 ( .A1(n40725), .A2(n40113), .B1(n41109), .B2(n40106), .C1(
        n25419), .C2(n40100), .ZN(n8333) );
  OAI222_X1 U32726 ( .A1(n40731), .A2(n40113), .B1(n41115), .B2(n40106), .C1(
        n25420), .C2(n40100), .ZN(n8332) );
  OAI222_X1 U32727 ( .A1(n40737), .A2(n40113), .B1(n41121), .B2(n40106), .C1(
        n25421), .C2(n40100), .ZN(n8331) );
  OAI222_X1 U32728 ( .A1(n40743), .A2(n40113), .B1(n41127), .B2(n40106), .C1(
        n25422), .C2(n40100), .ZN(n8330) );
  OAI222_X1 U32729 ( .A1(n40749), .A2(n40113), .B1(n41133), .B2(n40106), .C1(
        n25423), .C2(n40100), .ZN(n8329) );
  OAI222_X1 U32730 ( .A1(n40755), .A2(n40113), .B1(n41139), .B2(n40106), .C1(
        n25424), .C2(n40099), .ZN(n8328) );
  OAI222_X1 U32731 ( .A1(n40761), .A2(n40113), .B1(n41145), .B2(n40106), .C1(
        n25425), .C2(n40099), .ZN(n8327) );
  OAI222_X1 U32732 ( .A1(n40767), .A2(n40112), .B1(n41151), .B2(n40105), .C1(
        n25426), .C2(n40099), .ZN(n8326) );
  OAI222_X1 U32733 ( .A1(n40773), .A2(n40112), .B1(n41157), .B2(n40105), .C1(
        n25427), .C2(n40099), .ZN(n8325) );
  OAI222_X1 U32734 ( .A1(n40779), .A2(n40112), .B1(n41163), .B2(n40105), .C1(
        n25428), .C2(n40099), .ZN(n8324) );
  OAI222_X1 U32735 ( .A1(n40785), .A2(n40112), .B1(n41169), .B2(n40105), .C1(
        n25429), .C2(n40099), .ZN(n8323) );
  OAI222_X1 U32736 ( .A1(n40791), .A2(n40112), .B1(n41175), .B2(n40105), .C1(
        n25430), .C2(n40099), .ZN(n8322) );
  OAI222_X1 U32737 ( .A1(n40797), .A2(n40112), .B1(n41181), .B2(n40105), .C1(
        n25431), .C2(n40099), .ZN(n8321) );
  OAI222_X1 U32738 ( .A1(n40803), .A2(n40112), .B1(n41187), .B2(n40105), .C1(
        n25432), .C2(n40099), .ZN(n8320) );
  OAI222_X1 U32739 ( .A1(n40809), .A2(n40112), .B1(n41193), .B2(n40105), .C1(
        n25433), .C2(n40099), .ZN(n8319) );
  OAI222_X1 U32740 ( .A1(n40815), .A2(n40112), .B1(n41199), .B2(n40105), .C1(
        n25434), .C2(n40099), .ZN(n8318) );
  OAI222_X1 U32741 ( .A1(n40821), .A2(n40112), .B1(n41205), .B2(n40105), .C1(
        n25435), .C2(n40099), .ZN(n8317) );
  OAI222_X1 U32742 ( .A1(n40827), .A2(n40112), .B1(n41211), .B2(n40105), .C1(
        n25436), .C2(n40099), .ZN(n8316) );
  OAI222_X1 U32743 ( .A1(n40833), .A2(n40112), .B1(n41217), .B2(n40105), .C1(
        n25437), .C2(n40098), .ZN(n8315) );
  OAI222_X1 U32744 ( .A1(n40839), .A2(n40111), .B1(n41223), .B2(n40104), .C1(
        n25438), .C2(n40098), .ZN(n8314) );
  OAI222_X1 U32745 ( .A1(n40845), .A2(n40111), .B1(n41229), .B2(n40104), .C1(
        n25439), .C2(n40098), .ZN(n8313) );
  OAI222_X1 U32746 ( .A1(n40851), .A2(n40111), .B1(n41235), .B2(n40104), .C1(
        n25440), .C2(n40098), .ZN(n8312) );
  OAI222_X1 U32747 ( .A1(n40857), .A2(n40111), .B1(n41241), .B2(n40104), .C1(
        n25441), .C2(n40098), .ZN(n8311) );
  OAI222_X1 U32748 ( .A1(n40863), .A2(n40111), .B1(n41247), .B2(n40104), .C1(
        n25442), .C2(n40098), .ZN(n8310) );
  OAI222_X1 U32749 ( .A1(n40869), .A2(n40111), .B1(n41253), .B2(n40104), .C1(
        n25443), .C2(n40098), .ZN(n8309) );
  OAI222_X1 U32750 ( .A1(n40875), .A2(n40111), .B1(n41259), .B2(n40104), .C1(
        n25444), .C2(n40098), .ZN(n8308) );
  OAI222_X1 U32751 ( .A1(n40881), .A2(n40111), .B1(n41265), .B2(n40104), .C1(
        n25445), .C2(n40098), .ZN(n8307) );
  OAI222_X1 U32752 ( .A1(n40887), .A2(n40111), .B1(n41271), .B2(n40104), .C1(
        n25446), .C2(n40098), .ZN(n8306) );
  OAI222_X1 U32753 ( .A1(n40893), .A2(n40111), .B1(n41277), .B2(n40104), .C1(
        n25447), .C2(n40098), .ZN(n8305) );
  OAI222_X1 U32754 ( .A1(n40899), .A2(n40111), .B1(n41283), .B2(n40104), .C1(
        n25448), .C2(n40098), .ZN(n8304) );
  OAI222_X1 U32755 ( .A1(n40905), .A2(n40111), .B1(n41289), .B2(n40104), .C1(
        n25449), .C2(n40098), .ZN(n8303) );
  OAI222_X1 U32756 ( .A1(n40911), .A2(n40110), .B1(n41295), .B2(n40103), .C1(
        n25450), .C2(n40097), .ZN(n8302) );
  OAI222_X1 U32757 ( .A1(n40917), .A2(n40110), .B1(n41301), .B2(n40103), .C1(
        n25451), .C2(n40097), .ZN(n8301) );
  OAI222_X1 U32758 ( .A1(n40923), .A2(n40110), .B1(n41307), .B2(n40103), .C1(
        n25452), .C2(n40097), .ZN(n8300) );
  OAI222_X1 U32759 ( .A1(n40929), .A2(n40110), .B1(n41313), .B2(n40103), .C1(
        n25453), .C2(n40097), .ZN(n8299) );
  OAI222_X1 U32760 ( .A1(n40935), .A2(n40110), .B1(n41319), .B2(n40103), .C1(
        n25454), .C2(n40097), .ZN(n8298) );
  OAI222_X1 U32761 ( .A1(n40941), .A2(n40110), .B1(n41325), .B2(n40103), .C1(
        n25455), .C2(n40097), .ZN(n8297) );
  OAI222_X1 U32762 ( .A1(n40947), .A2(n40110), .B1(n41331), .B2(n40103), .C1(
        n25456), .C2(n40097), .ZN(n8296) );
  OAI222_X1 U32763 ( .A1(n40953), .A2(n40110), .B1(n41337), .B2(n40103), .C1(
        n28840), .C2(n40097), .ZN(n8295) );
  OAI222_X1 U32764 ( .A1(n40959), .A2(n40110), .B1(n41343), .B2(n40103), .C1(
        n25457), .C2(n40097), .ZN(n8294) );
  OAI222_X1 U32765 ( .A1(n40965), .A2(n40110), .B1(n41349), .B2(n40103), .C1(
        n25395), .C2(n40097), .ZN(n8293) );
  OAI222_X1 U32766 ( .A1(n40971), .A2(n40110), .B1(n41355), .B2(n40103), .C1(
        n25396), .C2(n40097), .ZN(n8292) );
  OAI222_X1 U32767 ( .A1(n40977), .A2(n40110), .B1(n41361), .B2(n40103), .C1(
        n25397), .C2(n40097), .ZN(n8291) );
  OAI222_X1 U32768 ( .A1(n40598), .A2(n39820), .B1(n40982), .B2(n39813), .C1(
        n27943), .C2(n39806), .ZN(n7394) );
  OAI222_X1 U32769 ( .A1(n40604), .A2(n39820), .B1(n40988), .B2(n39813), .C1(
        n27942), .C2(n39806), .ZN(n7393) );
  OAI222_X1 U32770 ( .A1(n40610), .A2(n39820), .B1(n40994), .B2(n39813), .C1(
        n27941), .C2(n39806), .ZN(n7392) );
  OAI222_X1 U32771 ( .A1(n40616), .A2(n39820), .B1(n41000), .B2(n39813), .C1(
        n27940), .C2(n39806), .ZN(n7391) );
  OAI222_X1 U32772 ( .A1(n40622), .A2(n39819), .B1(n41006), .B2(n39812), .C1(
        n27939), .C2(n39806), .ZN(n7390) );
  OAI222_X1 U32773 ( .A1(n40628), .A2(n39819), .B1(n41012), .B2(n39812), .C1(
        n27938), .C2(n39806), .ZN(n7389) );
  OAI222_X1 U32774 ( .A1(n40634), .A2(n39819), .B1(n41018), .B2(n39812), .C1(
        n27937), .C2(n39806), .ZN(n7388) );
  OAI222_X1 U32775 ( .A1(n40640), .A2(n39819), .B1(n41024), .B2(n39812), .C1(
        n27936), .C2(n39806), .ZN(n7387) );
  OAI222_X1 U32776 ( .A1(n40646), .A2(n39819), .B1(n41030), .B2(n39812), .C1(
        n27935), .C2(n39806), .ZN(n7386) );
  OAI222_X1 U32777 ( .A1(n40652), .A2(n39819), .B1(n41036), .B2(n39812), .C1(
        n27934), .C2(n39806), .ZN(n7385) );
  OAI222_X1 U32778 ( .A1(n40658), .A2(n39819), .B1(n41042), .B2(n39812), .C1(
        n27933), .C2(n39806), .ZN(n7384) );
  OAI222_X1 U32779 ( .A1(n40664), .A2(n39819), .B1(n41048), .B2(n39812), .C1(
        n27932), .C2(n39806), .ZN(n7383) );
  OAI222_X1 U32780 ( .A1(n40670), .A2(n39819), .B1(n41054), .B2(n39812), .C1(
        n27931), .C2(n39806), .ZN(n7382) );
  OAI222_X1 U32781 ( .A1(n40676), .A2(n39819), .B1(n41060), .B2(n39812), .C1(
        n27930), .C2(n39805), .ZN(n7381) );
  OAI222_X1 U32782 ( .A1(n40682), .A2(n39819), .B1(n41066), .B2(n39812), .C1(
        n27929), .C2(n39805), .ZN(n7380) );
  OAI222_X1 U32783 ( .A1(n40688), .A2(n39819), .B1(n41072), .B2(n39812), .C1(
        n27928), .C2(n39805), .ZN(n7379) );
  OAI222_X1 U32784 ( .A1(n40694), .A2(n39818), .B1(n41078), .B2(n39811), .C1(
        n27927), .C2(n39805), .ZN(n7378) );
  OAI222_X1 U32785 ( .A1(n40700), .A2(n39818), .B1(n41084), .B2(n39811), .C1(
        n27926), .C2(n39805), .ZN(n7377) );
  OAI222_X1 U32786 ( .A1(n40706), .A2(n39818), .B1(n41090), .B2(n39811), .C1(
        n27925), .C2(n39805), .ZN(n7376) );
  OAI222_X1 U32787 ( .A1(n40712), .A2(n39818), .B1(n41096), .B2(n39811), .C1(
        n27924), .C2(n39805), .ZN(n7375) );
  OAI222_X1 U32788 ( .A1(n40718), .A2(n39818), .B1(n41102), .B2(n39811), .C1(
        n27923), .C2(n39805), .ZN(n7374) );
  OAI222_X1 U32789 ( .A1(n40724), .A2(n39818), .B1(n41108), .B2(n39811), .C1(
        n27922), .C2(n39805), .ZN(n7373) );
  OAI222_X1 U32790 ( .A1(n40730), .A2(n39818), .B1(n41114), .B2(n39811), .C1(
        n27921), .C2(n39805), .ZN(n7372) );
  OAI222_X1 U32791 ( .A1(n40912), .A2(n40430), .B1(n41296), .B2(n40423), .C1(
        n40420), .C2(n38794), .ZN(n9326) );
  OAI222_X1 U32792 ( .A1(n40918), .A2(n40430), .B1(n41302), .B2(n40423), .C1(
        n40420), .C2(n38795), .ZN(n9325) );
  OAI222_X1 U32793 ( .A1(n40924), .A2(n40430), .B1(n41308), .B2(n40423), .C1(
        n40420), .C2(n38796), .ZN(n9324) );
  OAI222_X1 U32794 ( .A1(n40930), .A2(n40430), .B1(n41314), .B2(n40423), .C1(
        n40420), .C2(n38797), .ZN(n9323) );
  OAI222_X1 U32795 ( .A1(n40936), .A2(n40430), .B1(n41320), .B2(n40423), .C1(
        n40420), .C2(n38798), .ZN(n9322) );
  OAI222_X1 U32796 ( .A1(n40942), .A2(n40430), .B1(n41326), .B2(n40423), .C1(
        n40420), .C2(n38799), .ZN(n9321) );
  OAI222_X1 U32797 ( .A1(n40948), .A2(n40430), .B1(n41332), .B2(n40423), .C1(
        n40420), .C2(n38800), .ZN(n9320) );
  OAI222_X1 U32798 ( .A1(n40960), .A2(n40430), .B1(n41344), .B2(n40423), .C1(
        n40420), .C2(n38801), .ZN(n9318) );
  OAI222_X1 U32799 ( .A1(n40624), .A2(n40434), .B1(n41008), .B2(n40427), .C1(
        n40416), .C2(n38802), .ZN(n9374) );
  OAI222_X1 U32800 ( .A1(n40630), .A2(n40434), .B1(n41014), .B2(n40427), .C1(
        n40416), .C2(n38803), .ZN(n9373) );
  OAI222_X1 U32801 ( .A1(n40636), .A2(n40434), .B1(n41020), .B2(n40427), .C1(
        n40416), .C2(n38804), .ZN(n9372) );
  OAI222_X1 U32802 ( .A1(n40642), .A2(n40434), .B1(n41026), .B2(n40427), .C1(
        n40416), .C2(n38805), .ZN(n9371) );
  OAI222_X1 U32803 ( .A1(n40648), .A2(n40434), .B1(n41032), .B2(n40427), .C1(
        n40416), .C2(n38806), .ZN(n9370) );
  OAI222_X1 U32804 ( .A1(n40654), .A2(n40434), .B1(n41038), .B2(n40427), .C1(
        n40416), .C2(n38807), .ZN(n9369) );
  OAI222_X1 U32805 ( .A1(n40660), .A2(n40434), .B1(n41044), .B2(n40427), .C1(
        n40416), .C2(n38808), .ZN(n9368) );
  OAI222_X1 U32806 ( .A1(n40666), .A2(n40434), .B1(n41050), .B2(n40427), .C1(
        n40416), .C2(n38809), .ZN(n9367) );
  OAI222_X1 U32807 ( .A1(n40672), .A2(n40434), .B1(n41056), .B2(n40427), .C1(
        n40417), .C2(n38810), .ZN(n9366) );
  OAI222_X1 U32808 ( .A1(n40678), .A2(n40434), .B1(n41062), .B2(n40427), .C1(
        n40417), .C2(n38811), .ZN(n9365) );
  OAI222_X1 U32809 ( .A1(n40684), .A2(n40434), .B1(n41068), .B2(n40427), .C1(
        n40417), .C2(n38812), .ZN(n9364) );
  OAI222_X1 U32810 ( .A1(n40690), .A2(n40434), .B1(n41074), .B2(n40427), .C1(
        n40418), .C2(n38813), .ZN(n9363) );
  OAI222_X1 U32811 ( .A1(n40696), .A2(n40433), .B1(n41080), .B2(n40426), .C1(
        n40417), .C2(n38814), .ZN(n9362) );
  OAI222_X1 U32812 ( .A1(n40702), .A2(n40433), .B1(n41086), .B2(n40426), .C1(
        n40417), .C2(n38815), .ZN(n9361) );
  OAI222_X1 U32813 ( .A1(n40708), .A2(n40433), .B1(n41092), .B2(n40426), .C1(
        n40417), .C2(n38816), .ZN(n9360) );
  OAI222_X1 U32814 ( .A1(n40714), .A2(n40433), .B1(n41098), .B2(n40426), .C1(
        n40417), .C2(n38817), .ZN(n9359) );
  OAI222_X1 U32815 ( .A1(n40720), .A2(n40433), .B1(n41104), .B2(n40426), .C1(
        n40417), .C2(n38818), .ZN(n9358) );
  OAI222_X1 U32816 ( .A1(n40726), .A2(n40433), .B1(n41110), .B2(n40426), .C1(
        n40417), .C2(n38819), .ZN(n9357) );
  OAI222_X1 U32817 ( .A1(n40732), .A2(n40433), .B1(n41116), .B2(n40426), .C1(
        n40417), .C2(n38820), .ZN(n9356) );
  OAI222_X1 U32818 ( .A1(n40738), .A2(n40433), .B1(n41122), .B2(n40426), .C1(
        n40417), .C2(n38821), .ZN(n9355) );
  OAI222_X1 U32819 ( .A1(n40744), .A2(n40433), .B1(n41128), .B2(n40426), .C1(
        n40417), .C2(n38822), .ZN(n9354) );
  OAI222_X1 U32820 ( .A1(n40750), .A2(n40433), .B1(n41134), .B2(n40426), .C1(
        n40418), .C2(n38823), .ZN(n9353) );
  OAI222_X1 U32821 ( .A1(n40756), .A2(n40433), .B1(n41140), .B2(n40426), .C1(
        n40418), .C2(n38824), .ZN(n9352) );
  OAI222_X1 U32822 ( .A1(n40762), .A2(n40433), .B1(n41146), .B2(n40426), .C1(
        n40418), .C2(n38825), .ZN(n9351) );
  OAI222_X1 U32823 ( .A1(n40768), .A2(n40432), .B1(n41152), .B2(n40425), .C1(
        n40418), .C2(n38826), .ZN(n9350) );
  OAI222_X1 U32824 ( .A1(n40774), .A2(n40432), .B1(n41158), .B2(n40425), .C1(
        n40418), .C2(n38827), .ZN(n9349) );
  OAI222_X1 U32825 ( .A1(n40780), .A2(n40432), .B1(n41164), .B2(n40425), .C1(
        n40418), .C2(n38828), .ZN(n9348) );
  OAI222_X1 U32826 ( .A1(n40786), .A2(n40432), .B1(n41170), .B2(n40425), .C1(
        n40418), .C2(n38829), .ZN(n9347) );
  OAI222_X1 U32827 ( .A1(n40792), .A2(n40432), .B1(n41176), .B2(n40425), .C1(
        n40418), .C2(n38830), .ZN(n9346) );
  OAI222_X1 U32828 ( .A1(n40798), .A2(n40432), .B1(n41182), .B2(n40425), .C1(
        n40418), .C2(n38831), .ZN(n9345) );
  OAI222_X1 U32829 ( .A1(n40804), .A2(n40432), .B1(n41188), .B2(n40425), .C1(
        n40418), .C2(n38832), .ZN(n9344) );
  OAI222_X1 U32830 ( .A1(n40810), .A2(n40432), .B1(n41194), .B2(n40425), .C1(
        n40418), .C2(n38833), .ZN(n9343) );
  OAI222_X1 U32831 ( .A1(n40816), .A2(n40432), .B1(n41200), .B2(n40425), .C1(
        n40419), .C2(n38834), .ZN(n9342) );
  OAI222_X1 U32832 ( .A1(n40822), .A2(n40432), .B1(n41206), .B2(n40425), .C1(
        n40419), .C2(n38835), .ZN(n9341) );
  OAI222_X1 U32833 ( .A1(n40828), .A2(n40432), .B1(n41212), .B2(n40425), .C1(
        n40419), .C2(n38836), .ZN(n9340) );
  OAI222_X1 U32834 ( .A1(n40834), .A2(n40432), .B1(n41218), .B2(n40425), .C1(
        n40419), .C2(n38837), .ZN(n9339) );
  OAI222_X1 U32835 ( .A1(n40840), .A2(n40431), .B1(n41224), .B2(n40424), .C1(
        n40419), .C2(n38838), .ZN(n9338) );
  OAI222_X1 U32836 ( .A1(n40846), .A2(n40431), .B1(n41230), .B2(n40424), .C1(
        n40419), .C2(n38839), .ZN(n9337) );
  OAI222_X1 U32837 ( .A1(n40852), .A2(n40431), .B1(n41236), .B2(n40424), .C1(
        n40419), .C2(n38840), .ZN(n9336) );
  OAI222_X1 U32838 ( .A1(n40858), .A2(n40431), .B1(n41242), .B2(n40424), .C1(
        n40419), .C2(n38841), .ZN(n9335) );
  OAI222_X1 U32839 ( .A1(n40864), .A2(n40431), .B1(n41248), .B2(n40424), .C1(
        n40419), .C2(n38842), .ZN(n9334) );
  OAI222_X1 U32840 ( .A1(n40870), .A2(n40431), .B1(n41254), .B2(n40424), .C1(
        n40419), .C2(n38843), .ZN(n9333) );
  OAI222_X1 U32841 ( .A1(n40876), .A2(n40431), .B1(n41260), .B2(n40424), .C1(
        n40419), .C2(n38844), .ZN(n9332) );
  OAI222_X1 U32842 ( .A1(n40882), .A2(n40431), .B1(n41266), .B2(n40424), .C1(
        n40419), .C2(n38845), .ZN(n9331) );
  OAI222_X1 U32843 ( .A1(n40888), .A2(n40431), .B1(n41272), .B2(n40424), .C1(
        n40420), .C2(n38846), .ZN(n9330) );
  OAI222_X1 U32844 ( .A1(n40894), .A2(n40431), .B1(n41278), .B2(n40424), .C1(
        n40420), .C2(n38847), .ZN(n9329) );
  OAI222_X1 U32845 ( .A1(n40900), .A2(n40431), .B1(n41284), .B2(n40424), .C1(
        n40420), .C2(n38848), .ZN(n9328) );
  OAI222_X1 U32846 ( .A1(n40906), .A2(n40431), .B1(n41290), .B2(n40424), .C1(
        n40420), .C2(n38849), .ZN(n9327) );
  OAI222_X1 U32847 ( .A1(n40912), .A2(n40410), .B1(n41296), .B2(n40403), .C1(
        n40400), .C2(n38927), .ZN(n9262) );
  OAI222_X1 U32848 ( .A1(n40918), .A2(n40410), .B1(n41302), .B2(n40403), .C1(
        n40400), .C2(n38928), .ZN(n9261) );
  OAI222_X1 U32849 ( .A1(n40924), .A2(n40410), .B1(n41308), .B2(n40403), .C1(
        n40400), .C2(n38929), .ZN(n9260) );
  OAI222_X1 U32850 ( .A1(n40930), .A2(n40410), .B1(n41314), .B2(n40403), .C1(
        n40400), .C2(n38930), .ZN(n9259) );
  OAI222_X1 U32851 ( .A1(n40936), .A2(n40410), .B1(n41320), .B2(n40403), .C1(
        n40400), .C2(n38931), .ZN(n9258) );
  OAI222_X1 U32852 ( .A1(n40942), .A2(n40410), .B1(n41326), .B2(n40403), .C1(
        n40400), .C2(n38932), .ZN(n9257) );
  OAI222_X1 U32853 ( .A1(n40948), .A2(n40410), .B1(n41332), .B2(n40403), .C1(
        n40400), .C2(n38933), .ZN(n9256) );
  OAI222_X1 U32854 ( .A1(n40960), .A2(n40410), .B1(n41344), .B2(n40403), .C1(
        n40400), .C2(n38934), .ZN(n9254) );
  OAI222_X1 U32855 ( .A1(n40911), .A2(n40210), .B1(n41295), .B2(n40203), .C1(
        n40200), .C2(n33110), .ZN(n8622) );
  OAI222_X1 U32856 ( .A1(n40917), .A2(n40210), .B1(n41301), .B2(n40203), .C1(
        n40200), .C2(n33109), .ZN(n8621) );
  OAI222_X1 U32857 ( .A1(n40923), .A2(n40210), .B1(n41307), .B2(n40203), .C1(
        n40200), .C2(n33108), .ZN(n8620) );
  OAI222_X1 U32858 ( .A1(n40929), .A2(n40210), .B1(n41313), .B2(n40203), .C1(
        n40200), .C2(n33107), .ZN(n8619) );
  OAI222_X1 U32859 ( .A1(n40935), .A2(n40210), .B1(n41319), .B2(n40203), .C1(
        n40200), .C2(n33106), .ZN(n8618) );
  OAI222_X1 U32860 ( .A1(n40941), .A2(n40210), .B1(n41325), .B2(n40203), .C1(
        n40200), .C2(n33105), .ZN(n8617) );
  OAI222_X1 U32861 ( .A1(n40947), .A2(n40210), .B1(n41331), .B2(n40203), .C1(
        n40200), .C2(n33104), .ZN(n8616) );
  OAI222_X1 U32862 ( .A1(n40959), .A2(n40210), .B1(n41343), .B2(n40203), .C1(
        n40200), .C2(n33102), .ZN(n8614) );
  OAI222_X1 U32863 ( .A1(n40911), .A2(n40230), .B1(n41295), .B2(n40223), .C1(
        n40220), .C2(n33098), .ZN(n8686) );
  OAI222_X1 U32864 ( .A1(n40917), .A2(n40230), .B1(n41301), .B2(n40223), .C1(
        n40220), .C2(n33097), .ZN(n8685) );
  OAI222_X1 U32865 ( .A1(n40923), .A2(n40230), .B1(n41307), .B2(n40223), .C1(
        n40220), .C2(n33096), .ZN(n8684) );
  OAI222_X1 U32866 ( .A1(n40929), .A2(n40230), .B1(n41313), .B2(n40223), .C1(
        n40220), .C2(n33095), .ZN(n8683) );
  OAI222_X1 U32867 ( .A1(n40935), .A2(n40230), .B1(n41319), .B2(n40223), .C1(
        n40220), .C2(n33094), .ZN(n8682) );
  OAI222_X1 U32868 ( .A1(n40941), .A2(n40230), .B1(n41325), .B2(n40223), .C1(
        n40220), .C2(n33093), .ZN(n8681) );
  OAI222_X1 U32869 ( .A1(n40947), .A2(n40230), .B1(n41331), .B2(n40223), .C1(
        n40220), .C2(n33092), .ZN(n8680) );
  OAI222_X1 U32870 ( .A1(n40959), .A2(n40230), .B1(n41343), .B2(n40223), .C1(
        n40220), .C2(n33090), .ZN(n8678) );
  OAI222_X1 U32871 ( .A1(n40624), .A2(n40414), .B1(n41008), .B2(n40407), .C1(
        n40396), .C2(n38935), .ZN(n9310) );
  OAI222_X1 U32872 ( .A1(n40630), .A2(n40414), .B1(n41014), .B2(n40407), .C1(
        n40396), .C2(n38936), .ZN(n9309) );
  OAI222_X1 U32873 ( .A1(n40636), .A2(n40414), .B1(n41020), .B2(n40407), .C1(
        n40396), .C2(n38937), .ZN(n9308) );
  OAI222_X1 U32874 ( .A1(n40642), .A2(n40414), .B1(n41026), .B2(n40407), .C1(
        n40396), .C2(n38938), .ZN(n9307) );
  OAI222_X1 U32875 ( .A1(n40648), .A2(n40414), .B1(n41032), .B2(n40407), .C1(
        n40396), .C2(n38939), .ZN(n9306) );
  OAI222_X1 U32876 ( .A1(n40654), .A2(n40414), .B1(n41038), .B2(n40407), .C1(
        n40396), .C2(n38940), .ZN(n9305) );
  OAI222_X1 U32877 ( .A1(n40660), .A2(n40414), .B1(n41044), .B2(n40407), .C1(
        n40396), .C2(n38941), .ZN(n9304) );
  OAI222_X1 U32878 ( .A1(n40666), .A2(n40414), .B1(n41050), .B2(n40407), .C1(
        n40396), .C2(n38942), .ZN(n9303) );
  OAI222_X1 U32879 ( .A1(n40672), .A2(n40414), .B1(n41056), .B2(n40407), .C1(
        n40397), .C2(n38943), .ZN(n9302) );
  OAI222_X1 U32880 ( .A1(n40678), .A2(n40414), .B1(n41062), .B2(n40407), .C1(
        n40397), .C2(n38944), .ZN(n9301) );
  OAI222_X1 U32881 ( .A1(n40684), .A2(n40414), .B1(n41068), .B2(n40407), .C1(
        n40397), .C2(n38945), .ZN(n9300) );
  OAI222_X1 U32882 ( .A1(n40690), .A2(n40414), .B1(n41074), .B2(n40407), .C1(
        n40398), .C2(n38946), .ZN(n9299) );
  OAI222_X1 U32883 ( .A1(n40696), .A2(n40413), .B1(n41080), .B2(n40406), .C1(
        n40397), .C2(n38947), .ZN(n9298) );
  OAI222_X1 U32884 ( .A1(n40702), .A2(n40413), .B1(n41086), .B2(n40406), .C1(
        n40397), .C2(n38948), .ZN(n9297) );
  OAI222_X1 U32885 ( .A1(n40708), .A2(n40413), .B1(n41092), .B2(n40406), .C1(
        n40397), .C2(n38949), .ZN(n9296) );
  OAI222_X1 U32886 ( .A1(n40714), .A2(n40413), .B1(n41098), .B2(n40406), .C1(
        n40397), .C2(n38950), .ZN(n9295) );
  OAI222_X1 U32887 ( .A1(n40720), .A2(n40413), .B1(n41104), .B2(n40406), .C1(
        n40397), .C2(n38951), .ZN(n9294) );
  OAI222_X1 U32888 ( .A1(n40726), .A2(n40413), .B1(n41110), .B2(n40406), .C1(
        n40397), .C2(n38952), .ZN(n9293) );
  OAI222_X1 U32889 ( .A1(n40732), .A2(n40413), .B1(n41116), .B2(n40406), .C1(
        n40397), .C2(n38953), .ZN(n9292) );
  OAI222_X1 U32890 ( .A1(n40738), .A2(n40413), .B1(n41122), .B2(n40406), .C1(
        n40397), .C2(n38954), .ZN(n9291) );
  OAI222_X1 U32891 ( .A1(n40744), .A2(n40413), .B1(n41128), .B2(n40406), .C1(
        n40397), .C2(n38955), .ZN(n9290) );
  OAI222_X1 U32892 ( .A1(n40750), .A2(n40413), .B1(n41134), .B2(n40406), .C1(
        n40398), .C2(n38956), .ZN(n9289) );
  OAI222_X1 U32893 ( .A1(n40756), .A2(n40413), .B1(n41140), .B2(n40406), .C1(
        n40398), .C2(n38957), .ZN(n9288) );
  OAI222_X1 U32894 ( .A1(n40762), .A2(n40413), .B1(n41146), .B2(n40406), .C1(
        n40398), .C2(n38958), .ZN(n9287) );
  OAI222_X1 U32895 ( .A1(n40768), .A2(n40412), .B1(n41152), .B2(n40405), .C1(
        n40398), .C2(n38959), .ZN(n9286) );
  OAI222_X1 U32896 ( .A1(n40774), .A2(n40412), .B1(n41158), .B2(n40405), .C1(
        n40398), .C2(n38960), .ZN(n9285) );
  OAI222_X1 U32897 ( .A1(n40780), .A2(n40412), .B1(n41164), .B2(n40405), .C1(
        n40398), .C2(n38961), .ZN(n9284) );
  OAI222_X1 U32898 ( .A1(n40786), .A2(n40412), .B1(n41170), .B2(n40405), .C1(
        n40398), .C2(n38962), .ZN(n9283) );
  OAI222_X1 U32899 ( .A1(n40792), .A2(n40412), .B1(n41176), .B2(n40405), .C1(
        n40398), .C2(n38963), .ZN(n9282) );
  OAI222_X1 U32900 ( .A1(n40798), .A2(n40412), .B1(n41182), .B2(n40405), .C1(
        n40398), .C2(n38964), .ZN(n9281) );
  OAI222_X1 U32901 ( .A1(n40804), .A2(n40412), .B1(n41188), .B2(n40405), .C1(
        n40398), .C2(n38965), .ZN(n9280) );
  OAI222_X1 U32902 ( .A1(n40810), .A2(n40412), .B1(n41194), .B2(n40405), .C1(
        n40398), .C2(n38966), .ZN(n9279) );
  OAI222_X1 U32903 ( .A1(n40816), .A2(n40412), .B1(n41200), .B2(n40405), .C1(
        n40399), .C2(n38967), .ZN(n9278) );
  OAI222_X1 U32904 ( .A1(n40822), .A2(n40412), .B1(n41206), .B2(n40405), .C1(
        n40399), .C2(n38968), .ZN(n9277) );
  OAI222_X1 U32905 ( .A1(n40828), .A2(n40412), .B1(n41212), .B2(n40405), .C1(
        n40399), .C2(n38969), .ZN(n9276) );
  OAI222_X1 U32906 ( .A1(n40834), .A2(n40412), .B1(n41218), .B2(n40405), .C1(
        n40399), .C2(n38970), .ZN(n9275) );
  OAI222_X1 U32907 ( .A1(n40840), .A2(n40411), .B1(n41224), .B2(n40404), .C1(
        n40399), .C2(n38971), .ZN(n9274) );
  OAI222_X1 U32908 ( .A1(n40846), .A2(n40411), .B1(n41230), .B2(n40404), .C1(
        n40399), .C2(n38972), .ZN(n9273) );
  OAI222_X1 U32909 ( .A1(n40852), .A2(n40411), .B1(n41236), .B2(n40404), .C1(
        n40399), .C2(n38973), .ZN(n9272) );
  OAI222_X1 U32910 ( .A1(n40858), .A2(n40411), .B1(n41242), .B2(n40404), .C1(
        n40399), .C2(n38974), .ZN(n9271) );
  OAI222_X1 U32911 ( .A1(n40864), .A2(n40411), .B1(n41248), .B2(n40404), .C1(
        n40399), .C2(n38975), .ZN(n9270) );
  OAI222_X1 U32912 ( .A1(n40870), .A2(n40411), .B1(n41254), .B2(n40404), .C1(
        n40399), .C2(n38976), .ZN(n9269) );
  OAI222_X1 U32913 ( .A1(n40876), .A2(n40411), .B1(n41260), .B2(n40404), .C1(
        n40399), .C2(n38977), .ZN(n9268) );
  OAI222_X1 U32914 ( .A1(n40882), .A2(n40411), .B1(n41266), .B2(n40404), .C1(
        n40399), .C2(n38978), .ZN(n9267) );
  OAI222_X1 U32915 ( .A1(n40888), .A2(n40411), .B1(n41272), .B2(n40404), .C1(
        n40400), .C2(n38979), .ZN(n9266) );
  OAI222_X1 U32916 ( .A1(n40894), .A2(n40411), .B1(n41278), .B2(n40404), .C1(
        n40400), .C2(n38980), .ZN(n9265) );
  OAI222_X1 U32917 ( .A1(n40900), .A2(n40411), .B1(n41284), .B2(n40404), .C1(
        n40400), .C2(n38981), .ZN(n9264) );
  OAI222_X1 U32918 ( .A1(n40906), .A2(n40411), .B1(n41290), .B2(n40404), .C1(
        n40400), .C2(n38982), .ZN(n9263) );
  OAI222_X1 U32919 ( .A1(n40623), .A2(n40214), .B1(n41007), .B2(n40207), .C1(
        n40196), .C2(n32942), .ZN(n8670) );
  OAI222_X1 U32920 ( .A1(n40629), .A2(n40214), .B1(n41013), .B2(n40207), .C1(
        n40196), .C2(n32941), .ZN(n8669) );
  OAI222_X1 U32921 ( .A1(n40635), .A2(n40214), .B1(n41019), .B2(n40207), .C1(
        n40196), .C2(n32940), .ZN(n8668) );
  OAI222_X1 U32922 ( .A1(n40641), .A2(n40214), .B1(n41025), .B2(n40207), .C1(
        n40196), .C2(n32939), .ZN(n8667) );
  OAI222_X1 U32923 ( .A1(n40647), .A2(n40214), .B1(n41031), .B2(n40207), .C1(
        n40196), .C2(n32938), .ZN(n8666) );
  OAI222_X1 U32924 ( .A1(n40653), .A2(n40214), .B1(n41037), .B2(n40207), .C1(
        n40196), .C2(n32937), .ZN(n8665) );
  OAI222_X1 U32925 ( .A1(n40659), .A2(n40214), .B1(n41043), .B2(n40207), .C1(
        n40196), .C2(n32936), .ZN(n8664) );
  OAI222_X1 U32926 ( .A1(n40665), .A2(n40214), .B1(n41049), .B2(n40207), .C1(
        n40196), .C2(n32935), .ZN(n8663) );
  OAI222_X1 U32927 ( .A1(n40671), .A2(n40214), .B1(n41055), .B2(n40207), .C1(
        n40197), .C2(n32934), .ZN(n8662) );
  OAI222_X1 U32928 ( .A1(n40677), .A2(n40214), .B1(n41061), .B2(n40207), .C1(
        n40197), .C2(n32933), .ZN(n8661) );
  OAI222_X1 U32929 ( .A1(n40683), .A2(n40214), .B1(n41067), .B2(n40207), .C1(
        n40197), .C2(n32932), .ZN(n8660) );
  OAI222_X1 U32930 ( .A1(n40689), .A2(n40214), .B1(n41073), .B2(n40207), .C1(
        n40198), .C2(n32931), .ZN(n8659) );
  OAI222_X1 U32931 ( .A1(n40695), .A2(n40213), .B1(n41079), .B2(n40206), .C1(
        n40197), .C2(n32930), .ZN(n8658) );
  OAI222_X1 U32932 ( .A1(n40701), .A2(n40213), .B1(n41085), .B2(n40206), .C1(
        n40197), .C2(n32929), .ZN(n8657) );
  OAI222_X1 U32933 ( .A1(n40707), .A2(n40213), .B1(n41091), .B2(n40206), .C1(
        n40197), .C2(n32928), .ZN(n8656) );
  OAI222_X1 U32934 ( .A1(n40713), .A2(n40213), .B1(n41097), .B2(n40206), .C1(
        n40197), .C2(n32927), .ZN(n8655) );
  OAI222_X1 U32935 ( .A1(n40719), .A2(n40213), .B1(n41103), .B2(n40206), .C1(
        n40197), .C2(n32926), .ZN(n8654) );
  OAI222_X1 U32936 ( .A1(n40725), .A2(n40213), .B1(n41109), .B2(n40206), .C1(
        n40197), .C2(n32925), .ZN(n8653) );
  OAI222_X1 U32937 ( .A1(n40731), .A2(n40213), .B1(n41115), .B2(n40206), .C1(
        n40197), .C2(n32924), .ZN(n8652) );
  OAI222_X1 U32938 ( .A1(n40737), .A2(n40213), .B1(n41121), .B2(n40206), .C1(
        n40197), .C2(n32923), .ZN(n8651) );
  OAI222_X1 U32939 ( .A1(n40743), .A2(n40213), .B1(n41127), .B2(n40206), .C1(
        n40197), .C2(n32922), .ZN(n8650) );
  OAI222_X1 U32940 ( .A1(n40749), .A2(n40213), .B1(n41133), .B2(n40206), .C1(
        n40198), .C2(n32921), .ZN(n8649) );
  OAI222_X1 U32941 ( .A1(n40755), .A2(n40213), .B1(n41139), .B2(n40206), .C1(
        n40198), .C2(n32920), .ZN(n8648) );
  OAI222_X1 U32942 ( .A1(n40761), .A2(n40213), .B1(n41145), .B2(n40206), .C1(
        n40198), .C2(n32919), .ZN(n8647) );
  OAI222_X1 U32943 ( .A1(n40767), .A2(n40212), .B1(n41151), .B2(n40205), .C1(
        n40198), .C2(n32918), .ZN(n8646) );
  OAI222_X1 U32944 ( .A1(n40773), .A2(n40212), .B1(n41157), .B2(n40205), .C1(
        n40198), .C2(n32917), .ZN(n8645) );
  OAI222_X1 U32945 ( .A1(n40779), .A2(n40212), .B1(n41163), .B2(n40205), .C1(
        n40198), .C2(n32916), .ZN(n8644) );
  OAI222_X1 U32946 ( .A1(n40785), .A2(n40212), .B1(n41169), .B2(n40205), .C1(
        n40198), .C2(n32915), .ZN(n8643) );
  OAI222_X1 U32947 ( .A1(n40791), .A2(n40212), .B1(n41175), .B2(n40205), .C1(
        n40198), .C2(n32914), .ZN(n8642) );
  OAI222_X1 U32948 ( .A1(n40797), .A2(n40212), .B1(n41181), .B2(n40205), .C1(
        n40198), .C2(n32913), .ZN(n8641) );
  OAI222_X1 U32949 ( .A1(n40803), .A2(n40212), .B1(n41187), .B2(n40205), .C1(
        n40198), .C2(n32912), .ZN(n8640) );
  OAI222_X1 U32950 ( .A1(n40809), .A2(n40212), .B1(n41193), .B2(n40205), .C1(
        n40198), .C2(n32911), .ZN(n8639) );
  OAI222_X1 U32951 ( .A1(n40815), .A2(n40212), .B1(n41199), .B2(n40205), .C1(
        n40199), .C2(n32910), .ZN(n8638) );
  OAI222_X1 U32952 ( .A1(n40821), .A2(n40212), .B1(n41205), .B2(n40205), .C1(
        n40199), .C2(n32909), .ZN(n8637) );
  OAI222_X1 U32953 ( .A1(n40827), .A2(n40212), .B1(n41211), .B2(n40205), .C1(
        n40199), .C2(n32908), .ZN(n8636) );
  OAI222_X1 U32954 ( .A1(n40833), .A2(n40212), .B1(n41217), .B2(n40205), .C1(
        n40199), .C2(n32907), .ZN(n8635) );
  OAI222_X1 U32955 ( .A1(n40839), .A2(n40211), .B1(n41223), .B2(n40204), .C1(
        n40199), .C2(n32906), .ZN(n8634) );
  OAI222_X1 U32956 ( .A1(n40845), .A2(n40211), .B1(n41229), .B2(n40204), .C1(
        n40199), .C2(n32905), .ZN(n8633) );
  OAI222_X1 U32957 ( .A1(n40851), .A2(n40211), .B1(n41235), .B2(n40204), .C1(
        n40199), .C2(n32904), .ZN(n8632) );
  OAI222_X1 U32958 ( .A1(n40857), .A2(n40211), .B1(n41241), .B2(n40204), .C1(
        n40199), .C2(n32903), .ZN(n8631) );
  OAI222_X1 U32959 ( .A1(n40863), .A2(n40211), .B1(n41247), .B2(n40204), .C1(
        n40199), .C2(n32902), .ZN(n8630) );
  OAI222_X1 U32960 ( .A1(n40869), .A2(n40211), .B1(n41253), .B2(n40204), .C1(
        n40199), .C2(n32901), .ZN(n8629) );
  OAI222_X1 U32961 ( .A1(n40875), .A2(n40211), .B1(n41259), .B2(n40204), .C1(
        n40199), .C2(n32900), .ZN(n8628) );
  OAI222_X1 U32962 ( .A1(n40881), .A2(n40211), .B1(n41265), .B2(n40204), .C1(
        n40199), .C2(n32899), .ZN(n8627) );
  OAI222_X1 U32963 ( .A1(n40887), .A2(n40211), .B1(n41271), .B2(n40204), .C1(
        n40200), .C2(n32898), .ZN(n8626) );
  OAI222_X1 U32964 ( .A1(n40893), .A2(n40211), .B1(n41277), .B2(n40204), .C1(
        n40200), .C2(n32897), .ZN(n8625) );
  OAI222_X1 U32965 ( .A1(n40899), .A2(n40211), .B1(n41283), .B2(n40204), .C1(
        n40200), .C2(n32896), .ZN(n8624) );
  OAI222_X1 U32966 ( .A1(n40905), .A2(n40211), .B1(n41289), .B2(n40204), .C1(
        n40200), .C2(n32895), .ZN(n8623) );
  OAI222_X1 U32967 ( .A1(n40623), .A2(n40234), .B1(n41007), .B2(n40227), .C1(
        n40216), .C2(n32894), .ZN(n8734) );
  OAI222_X1 U32968 ( .A1(n40629), .A2(n40234), .B1(n41013), .B2(n40227), .C1(
        n40216), .C2(n32893), .ZN(n8733) );
  OAI222_X1 U32969 ( .A1(n40635), .A2(n40234), .B1(n41019), .B2(n40227), .C1(
        n40216), .C2(n32892), .ZN(n8732) );
  OAI222_X1 U32970 ( .A1(n40641), .A2(n40234), .B1(n41025), .B2(n40227), .C1(
        n40216), .C2(n32891), .ZN(n8731) );
  OAI222_X1 U32971 ( .A1(n40647), .A2(n40234), .B1(n41031), .B2(n40227), .C1(
        n40216), .C2(n32890), .ZN(n8730) );
  OAI222_X1 U32972 ( .A1(n40653), .A2(n40234), .B1(n41037), .B2(n40227), .C1(
        n40216), .C2(n32889), .ZN(n8729) );
  OAI222_X1 U32973 ( .A1(n40659), .A2(n40234), .B1(n41043), .B2(n40227), .C1(
        n40216), .C2(n32888), .ZN(n8728) );
  OAI222_X1 U32974 ( .A1(n40665), .A2(n40234), .B1(n41049), .B2(n40227), .C1(
        n40216), .C2(n32887), .ZN(n8727) );
  OAI222_X1 U32975 ( .A1(n40671), .A2(n40234), .B1(n41055), .B2(n40227), .C1(
        n40217), .C2(n32886), .ZN(n8726) );
  OAI222_X1 U32976 ( .A1(n40677), .A2(n40234), .B1(n41061), .B2(n40227), .C1(
        n40217), .C2(n32885), .ZN(n8725) );
  OAI222_X1 U32977 ( .A1(n40683), .A2(n40234), .B1(n41067), .B2(n40227), .C1(
        n40217), .C2(n32884), .ZN(n8724) );
  OAI222_X1 U32978 ( .A1(n40689), .A2(n40234), .B1(n41073), .B2(n40227), .C1(
        n40218), .C2(n32883), .ZN(n8723) );
  OAI222_X1 U32979 ( .A1(n40695), .A2(n40233), .B1(n41079), .B2(n40226), .C1(
        n40217), .C2(n32882), .ZN(n8722) );
  OAI222_X1 U32980 ( .A1(n40701), .A2(n40233), .B1(n41085), .B2(n40226), .C1(
        n40217), .C2(n32881), .ZN(n8721) );
  OAI222_X1 U32981 ( .A1(n40707), .A2(n40233), .B1(n41091), .B2(n40226), .C1(
        n40217), .C2(n32880), .ZN(n8720) );
  OAI222_X1 U32982 ( .A1(n40713), .A2(n40233), .B1(n41097), .B2(n40226), .C1(
        n40217), .C2(n32879), .ZN(n8719) );
  OAI222_X1 U32983 ( .A1(n40719), .A2(n40233), .B1(n41103), .B2(n40226), .C1(
        n40217), .C2(n32878), .ZN(n8718) );
  OAI222_X1 U32984 ( .A1(n40725), .A2(n40233), .B1(n41109), .B2(n40226), .C1(
        n40217), .C2(n32877), .ZN(n8717) );
  OAI222_X1 U32985 ( .A1(n40731), .A2(n40233), .B1(n41115), .B2(n40226), .C1(
        n40217), .C2(n32876), .ZN(n8716) );
  OAI222_X1 U32986 ( .A1(n40737), .A2(n40233), .B1(n41121), .B2(n40226), .C1(
        n40217), .C2(n32875), .ZN(n8715) );
  OAI222_X1 U32987 ( .A1(n40743), .A2(n40233), .B1(n41127), .B2(n40226), .C1(
        n40217), .C2(n32874), .ZN(n8714) );
  OAI222_X1 U32988 ( .A1(n40749), .A2(n40233), .B1(n41133), .B2(n40226), .C1(
        n40218), .C2(n32873), .ZN(n8713) );
  OAI222_X1 U32989 ( .A1(n40755), .A2(n40233), .B1(n41139), .B2(n40226), .C1(
        n40218), .C2(n32872), .ZN(n8712) );
  OAI222_X1 U32990 ( .A1(n40761), .A2(n40233), .B1(n41145), .B2(n40226), .C1(
        n40218), .C2(n32871), .ZN(n8711) );
  OAI222_X1 U32991 ( .A1(n40767), .A2(n40232), .B1(n41151), .B2(n40225), .C1(
        n40218), .C2(n32870), .ZN(n8710) );
  OAI222_X1 U32992 ( .A1(n40773), .A2(n40232), .B1(n41157), .B2(n40225), .C1(
        n40218), .C2(n32869), .ZN(n8709) );
  OAI222_X1 U32993 ( .A1(n40779), .A2(n40232), .B1(n41163), .B2(n40225), .C1(
        n40218), .C2(n32868), .ZN(n8708) );
  OAI222_X1 U32994 ( .A1(n40785), .A2(n40232), .B1(n41169), .B2(n40225), .C1(
        n40218), .C2(n32867), .ZN(n8707) );
  OAI222_X1 U32995 ( .A1(n40791), .A2(n40232), .B1(n41175), .B2(n40225), .C1(
        n40218), .C2(n32866), .ZN(n8706) );
  OAI222_X1 U32996 ( .A1(n40797), .A2(n40232), .B1(n41181), .B2(n40225), .C1(
        n40218), .C2(n32865), .ZN(n8705) );
  OAI222_X1 U32997 ( .A1(n40803), .A2(n40232), .B1(n41187), .B2(n40225), .C1(
        n40218), .C2(n32864), .ZN(n8704) );
  OAI222_X1 U32998 ( .A1(n40809), .A2(n40232), .B1(n41193), .B2(n40225), .C1(
        n40218), .C2(n32863), .ZN(n8703) );
  OAI222_X1 U32999 ( .A1(n40815), .A2(n40232), .B1(n41199), .B2(n40225), .C1(
        n40219), .C2(n32862), .ZN(n8702) );
  OAI222_X1 U33000 ( .A1(n40821), .A2(n40232), .B1(n41205), .B2(n40225), .C1(
        n40219), .C2(n32861), .ZN(n8701) );
  OAI222_X1 U33001 ( .A1(n40827), .A2(n40232), .B1(n41211), .B2(n40225), .C1(
        n40219), .C2(n32860), .ZN(n8700) );
  OAI222_X1 U33002 ( .A1(n40833), .A2(n40232), .B1(n41217), .B2(n40225), .C1(
        n40219), .C2(n32859), .ZN(n8699) );
  OAI222_X1 U33003 ( .A1(n40839), .A2(n40231), .B1(n41223), .B2(n40224), .C1(
        n40219), .C2(n32858), .ZN(n8698) );
  OAI222_X1 U33004 ( .A1(n40845), .A2(n40231), .B1(n41229), .B2(n40224), .C1(
        n40219), .C2(n32857), .ZN(n8697) );
  OAI222_X1 U33005 ( .A1(n40851), .A2(n40231), .B1(n41235), .B2(n40224), .C1(
        n40219), .C2(n32856), .ZN(n8696) );
  OAI222_X1 U33006 ( .A1(n40857), .A2(n40231), .B1(n41241), .B2(n40224), .C1(
        n40219), .C2(n32855), .ZN(n8695) );
  OAI222_X1 U33007 ( .A1(n40863), .A2(n40231), .B1(n41247), .B2(n40224), .C1(
        n40219), .C2(n32854), .ZN(n8694) );
  OAI222_X1 U33008 ( .A1(n40869), .A2(n40231), .B1(n41253), .B2(n40224), .C1(
        n40219), .C2(n32853), .ZN(n8693) );
  OAI222_X1 U33009 ( .A1(n40875), .A2(n40231), .B1(n41259), .B2(n40224), .C1(
        n40219), .C2(n32852), .ZN(n8692) );
  OAI222_X1 U33010 ( .A1(n40881), .A2(n40231), .B1(n41265), .B2(n40224), .C1(
        n40219), .C2(n32851), .ZN(n8691) );
  OAI222_X1 U33011 ( .A1(n40887), .A2(n40231), .B1(n41271), .B2(n40224), .C1(
        n40220), .C2(n32850), .ZN(n8690) );
  OAI222_X1 U33012 ( .A1(n40893), .A2(n40231), .B1(n41277), .B2(n40224), .C1(
        n40220), .C2(n32849), .ZN(n8689) );
  OAI222_X1 U33013 ( .A1(n40899), .A2(n40231), .B1(n41283), .B2(n40224), .C1(
        n40220), .C2(n32848), .ZN(n8688) );
  OAI222_X1 U33014 ( .A1(n40905), .A2(n40231), .B1(n41289), .B2(n40224), .C1(
        n40220), .C2(n32847), .ZN(n8687) );
  OAI222_X1 U33015 ( .A1(n40912), .A2(n40310), .B1(n41296), .B2(n40303), .C1(
        n40300), .C2(n32726), .ZN(n8942) );
  OAI222_X1 U33016 ( .A1(n40918), .A2(n40310), .B1(n41302), .B2(n40303), .C1(
        n40300), .C2(n32725), .ZN(n8941) );
  OAI222_X1 U33017 ( .A1(n40924), .A2(n40310), .B1(n41308), .B2(n40303), .C1(
        n40300), .C2(n32724), .ZN(n8940) );
  OAI222_X1 U33018 ( .A1(n40930), .A2(n40310), .B1(n41314), .B2(n40303), .C1(
        n40300), .C2(n32723), .ZN(n8939) );
  OAI222_X1 U33019 ( .A1(n40936), .A2(n40310), .B1(n41320), .B2(n40303), .C1(
        n40300), .C2(n32722), .ZN(n8938) );
  OAI222_X1 U33020 ( .A1(n40942), .A2(n40310), .B1(n41326), .B2(n40303), .C1(
        n40300), .C2(n32721), .ZN(n8937) );
  OAI222_X1 U33021 ( .A1(n40948), .A2(n40310), .B1(n41332), .B2(n40303), .C1(
        n40300), .C2(n32720), .ZN(n8936) );
  OAI222_X1 U33022 ( .A1(n40960), .A2(n40310), .B1(n41344), .B2(n40303), .C1(
        n40300), .C2(n32718), .ZN(n8934) );
  OAI222_X1 U33023 ( .A1(n40912), .A2(n40330), .B1(n41296), .B2(n40323), .C1(
        n40320), .C2(n32714), .ZN(n9006) );
  OAI222_X1 U33024 ( .A1(n40918), .A2(n40330), .B1(n41302), .B2(n40323), .C1(
        n40320), .C2(n32713), .ZN(n9005) );
  OAI222_X1 U33025 ( .A1(n40924), .A2(n40330), .B1(n41308), .B2(n40323), .C1(
        n40320), .C2(n32712), .ZN(n9004) );
  OAI222_X1 U33026 ( .A1(n40930), .A2(n40330), .B1(n41314), .B2(n40323), .C1(
        n40320), .C2(n32711), .ZN(n9003) );
  OAI222_X1 U33027 ( .A1(n40936), .A2(n40330), .B1(n41320), .B2(n40323), .C1(
        n40320), .C2(n32710), .ZN(n9002) );
  OAI222_X1 U33028 ( .A1(n40942), .A2(n40330), .B1(n41326), .B2(n40323), .C1(
        n40320), .C2(n32709), .ZN(n9001) );
  OAI222_X1 U33029 ( .A1(n40948), .A2(n40330), .B1(n41332), .B2(n40323), .C1(
        n40320), .C2(n32708), .ZN(n9000) );
  OAI222_X1 U33030 ( .A1(n40960), .A2(n40330), .B1(n41344), .B2(n40323), .C1(
        n40320), .C2(n32706), .ZN(n8998) );
  OAI222_X1 U33031 ( .A1(n40910), .A2(n39835), .B1(n41294), .B2(n39828), .C1(
        n39825), .C2(n32702), .ZN(n7406) );
  OAI222_X1 U33032 ( .A1(n40916), .A2(n39835), .B1(n41300), .B2(n39828), .C1(
        n39825), .C2(n32701), .ZN(n7405) );
  OAI222_X1 U33033 ( .A1(n40922), .A2(n39835), .B1(n41306), .B2(n39828), .C1(
        n39825), .C2(n32700), .ZN(n7404) );
  OAI222_X1 U33034 ( .A1(n40928), .A2(n39835), .B1(n41312), .B2(n39828), .C1(
        n39825), .C2(n32699), .ZN(n7403) );
  OAI222_X1 U33035 ( .A1(n40934), .A2(n39835), .B1(n41318), .B2(n39828), .C1(
        n39825), .C2(n32698), .ZN(n7402) );
  OAI222_X1 U33036 ( .A1(n40940), .A2(n39835), .B1(n41324), .B2(n39828), .C1(
        n39825), .C2(n32697), .ZN(n7401) );
  OAI222_X1 U33037 ( .A1(n40946), .A2(n39835), .B1(n41330), .B2(n39828), .C1(
        n39825), .C2(n32696), .ZN(n7400) );
  OAI222_X1 U33038 ( .A1(n40958), .A2(n39835), .B1(n41342), .B2(n39828), .C1(
        n39825), .C2(n32694), .ZN(n7398) );
  OAI222_X1 U33039 ( .A1(n40624), .A2(n40314), .B1(n41008), .B2(n40307), .C1(
        n40296), .C2(n32690), .ZN(n8990) );
  OAI222_X1 U33040 ( .A1(n40630), .A2(n40314), .B1(n41014), .B2(n40307), .C1(
        n40296), .C2(n32689), .ZN(n8989) );
  OAI222_X1 U33041 ( .A1(n40636), .A2(n40314), .B1(n41020), .B2(n40307), .C1(
        n40296), .C2(n32688), .ZN(n8988) );
  OAI222_X1 U33042 ( .A1(n40642), .A2(n40314), .B1(n41026), .B2(n40307), .C1(
        n40296), .C2(n32687), .ZN(n8987) );
  OAI222_X1 U33043 ( .A1(n40648), .A2(n40314), .B1(n41032), .B2(n40307), .C1(
        n40296), .C2(n32686), .ZN(n8986) );
  OAI222_X1 U33044 ( .A1(n40654), .A2(n40314), .B1(n41038), .B2(n40307), .C1(
        n40296), .C2(n32685), .ZN(n8985) );
  OAI222_X1 U33045 ( .A1(n40660), .A2(n40314), .B1(n41044), .B2(n40307), .C1(
        n40296), .C2(n32684), .ZN(n8984) );
  OAI222_X1 U33046 ( .A1(n40666), .A2(n40314), .B1(n41050), .B2(n40307), .C1(
        n40296), .C2(n32683), .ZN(n8983) );
  OAI222_X1 U33047 ( .A1(n40672), .A2(n40314), .B1(n41056), .B2(n40307), .C1(
        n40297), .C2(n32682), .ZN(n8982) );
  OAI222_X1 U33048 ( .A1(n40678), .A2(n40314), .B1(n41062), .B2(n40307), .C1(
        n40297), .C2(n32681), .ZN(n8981) );
  OAI222_X1 U33049 ( .A1(n40684), .A2(n40314), .B1(n41068), .B2(n40307), .C1(
        n40297), .C2(n32680), .ZN(n8980) );
  OAI222_X1 U33050 ( .A1(n40690), .A2(n40314), .B1(n41074), .B2(n40307), .C1(
        n40298), .C2(n32679), .ZN(n8979) );
  OAI222_X1 U33051 ( .A1(n40696), .A2(n40313), .B1(n41080), .B2(n40306), .C1(
        n40297), .C2(n32678), .ZN(n8978) );
  OAI222_X1 U33052 ( .A1(n40702), .A2(n40313), .B1(n41086), .B2(n40306), .C1(
        n40297), .C2(n32677), .ZN(n8977) );
  OAI222_X1 U33053 ( .A1(n40708), .A2(n40313), .B1(n41092), .B2(n40306), .C1(
        n40297), .C2(n32676), .ZN(n8976) );
  OAI222_X1 U33054 ( .A1(n40714), .A2(n40313), .B1(n41098), .B2(n40306), .C1(
        n40297), .C2(n32675), .ZN(n8975) );
  OAI222_X1 U33055 ( .A1(n40720), .A2(n40313), .B1(n41104), .B2(n40306), .C1(
        n40297), .C2(n32674), .ZN(n8974) );
  OAI222_X1 U33056 ( .A1(n40726), .A2(n40313), .B1(n41110), .B2(n40306), .C1(
        n40297), .C2(n32673), .ZN(n8973) );
  OAI222_X1 U33057 ( .A1(n40732), .A2(n40313), .B1(n41116), .B2(n40306), .C1(
        n40297), .C2(n32672), .ZN(n8972) );
  OAI222_X1 U33058 ( .A1(n40738), .A2(n40313), .B1(n41122), .B2(n40306), .C1(
        n40297), .C2(n32671), .ZN(n8971) );
  OAI222_X1 U33059 ( .A1(n40744), .A2(n40313), .B1(n41128), .B2(n40306), .C1(
        n40297), .C2(n32670), .ZN(n8970) );
  OAI222_X1 U33060 ( .A1(n40750), .A2(n40313), .B1(n41134), .B2(n40306), .C1(
        n40298), .C2(n32669), .ZN(n8969) );
  OAI222_X1 U33061 ( .A1(n40756), .A2(n40313), .B1(n41140), .B2(n40306), .C1(
        n40298), .C2(n32668), .ZN(n8968) );
  OAI222_X1 U33062 ( .A1(n40762), .A2(n40313), .B1(n41146), .B2(n40306), .C1(
        n40298), .C2(n32667), .ZN(n8967) );
  OAI222_X1 U33063 ( .A1(n40768), .A2(n40312), .B1(n41152), .B2(n40305), .C1(
        n40298), .C2(n32666), .ZN(n8966) );
  OAI222_X1 U33064 ( .A1(n40774), .A2(n40312), .B1(n41158), .B2(n40305), .C1(
        n40298), .C2(n32665), .ZN(n8965) );
  OAI222_X1 U33065 ( .A1(n40780), .A2(n40312), .B1(n41164), .B2(n40305), .C1(
        n40298), .C2(n32664), .ZN(n8964) );
  OAI222_X1 U33066 ( .A1(n40786), .A2(n40312), .B1(n41170), .B2(n40305), .C1(
        n40298), .C2(n32663), .ZN(n8963) );
  OAI222_X1 U33067 ( .A1(n40792), .A2(n40312), .B1(n41176), .B2(n40305), .C1(
        n40298), .C2(n32662), .ZN(n8962) );
  OAI222_X1 U33068 ( .A1(n40798), .A2(n40312), .B1(n41182), .B2(n40305), .C1(
        n40298), .C2(n32661), .ZN(n8961) );
  OAI222_X1 U33069 ( .A1(n40804), .A2(n40312), .B1(n41188), .B2(n40305), .C1(
        n40298), .C2(n32660), .ZN(n8960) );
  OAI222_X1 U33070 ( .A1(n40810), .A2(n40312), .B1(n41194), .B2(n40305), .C1(
        n40298), .C2(n32659), .ZN(n8959) );
  OAI222_X1 U33071 ( .A1(n40816), .A2(n40312), .B1(n41200), .B2(n40305), .C1(
        n40299), .C2(n32658), .ZN(n8958) );
  OAI222_X1 U33072 ( .A1(n40822), .A2(n40312), .B1(n41206), .B2(n40305), .C1(
        n40299), .C2(n32657), .ZN(n8957) );
  OAI222_X1 U33073 ( .A1(n40828), .A2(n40312), .B1(n41212), .B2(n40305), .C1(
        n40299), .C2(n32656), .ZN(n8956) );
  OAI222_X1 U33074 ( .A1(n40834), .A2(n40312), .B1(n41218), .B2(n40305), .C1(
        n40299), .C2(n32655), .ZN(n8955) );
  OAI222_X1 U33075 ( .A1(n40840), .A2(n40311), .B1(n41224), .B2(n40304), .C1(
        n40299), .C2(n32654), .ZN(n8954) );
  OAI222_X1 U33076 ( .A1(n40846), .A2(n40311), .B1(n41230), .B2(n40304), .C1(
        n40299), .C2(n32653), .ZN(n8953) );
  OAI222_X1 U33077 ( .A1(n40852), .A2(n40311), .B1(n41236), .B2(n40304), .C1(
        n40299), .C2(n32652), .ZN(n8952) );
  OAI222_X1 U33078 ( .A1(n40858), .A2(n40311), .B1(n41242), .B2(n40304), .C1(
        n40299), .C2(n32651), .ZN(n8951) );
  OAI222_X1 U33079 ( .A1(n40864), .A2(n40311), .B1(n41248), .B2(n40304), .C1(
        n40299), .C2(n32650), .ZN(n8950) );
  OAI222_X1 U33080 ( .A1(n40870), .A2(n40311), .B1(n41254), .B2(n40304), .C1(
        n40299), .C2(n32649), .ZN(n8949) );
  OAI222_X1 U33081 ( .A1(n40876), .A2(n40311), .B1(n41260), .B2(n40304), .C1(
        n40299), .C2(n32648), .ZN(n8948) );
  OAI222_X1 U33082 ( .A1(n40882), .A2(n40311), .B1(n41266), .B2(n40304), .C1(
        n40299), .C2(n32647), .ZN(n8947) );
  OAI222_X1 U33083 ( .A1(n40888), .A2(n40311), .B1(n41272), .B2(n40304), .C1(
        n40300), .C2(n32646), .ZN(n8946) );
  OAI222_X1 U33084 ( .A1(n40894), .A2(n40311), .B1(n41278), .B2(n40304), .C1(
        n40300), .C2(n32645), .ZN(n8945) );
  OAI222_X1 U33085 ( .A1(n40900), .A2(n40311), .B1(n41284), .B2(n40304), .C1(
        n40300), .C2(n32644), .ZN(n8944) );
  OAI222_X1 U33086 ( .A1(n40906), .A2(n40311), .B1(n41290), .B2(n40304), .C1(
        n40300), .C2(n32643), .ZN(n8943) );
  OAI222_X1 U33087 ( .A1(n40624), .A2(n40334), .B1(n41008), .B2(n40327), .C1(
        n40316), .C2(n32642), .ZN(n9054) );
  OAI222_X1 U33088 ( .A1(n40630), .A2(n40334), .B1(n41014), .B2(n40327), .C1(
        n40316), .C2(n32641), .ZN(n9053) );
  OAI222_X1 U33089 ( .A1(n40636), .A2(n40334), .B1(n41020), .B2(n40327), .C1(
        n40316), .C2(n32640), .ZN(n9052) );
  OAI222_X1 U33090 ( .A1(n40642), .A2(n40334), .B1(n41026), .B2(n40327), .C1(
        n40316), .C2(n32639), .ZN(n9051) );
  OAI222_X1 U33091 ( .A1(n40648), .A2(n40334), .B1(n41032), .B2(n40327), .C1(
        n40316), .C2(n32638), .ZN(n9050) );
  OAI222_X1 U33092 ( .A1(n40654), .A2(n40334), .B1(n41038), .B2(n40327), .C1(
        n40316), .C2(n32637), .ZN(n9049) );
  OAI222_X1 U33093 ( .A1(n40660), .A2(n40334), .B1(n41044), .B2(n40327), .C1(
        n40316), .C2(n32636), .ZN(n9048) );
  OAI222_X1 U33094 ( .A1(n40666), .A2(n40334), .B1(n41050), .B2(n40327), .C1(
        n40316), .C2(n32635), .ZN(n9047) );
  OAI222_X1 U33095 ( .A1(n40672), .A2(n40334), .B1(n41056), .B2(n40327), .C1(
        n40317), .C2(n32634), .ZN(n9046) );
  OAI222_X1 U33096 ( .A1(n40678), .A2(n40334), .B1(n41062), .B2(n40327), .C1(
        n40317), .C2(n32633), .ZN(n9045) );
  OAI222_X1 U33097 ( .A1(n40684), .A2(n40334), .B1(n41068), .B2(n40327), .C1(
        n40317), .C2(n32632), .ZN(n9044) );
  OAI222_X1 U33098 ( .A1(n40690), .A2(n40334), .B1(n41074), .B2(n40327), .C1(
        n40318), .C2(n32631), .ZN(n9043) );
  OAI222_X1 U33099 ( .A1(n40696), .A2(n40333), .B1(n41080), .B2(n40326), .C1(
        n40317), .C2(n32630), .ZN(n9042) );
  OAI222_X1 U33100 ( .A1(n40702), .A2(n40333), .B1(n41086), .B2(n40326), .C1(
        n40317), .C2(n32629), .ZN(n9041) );
  OAI222_X1 U33101 ( .A1(n40708), .A2(n40333), .B1(n41092), .B2(n40326), .C1(
        n40317), .C2(n32628), .ZN(n9040) );
  OAI222_X1 U33102 ( .A1(n40714), .A2(n40333), .B1(n41098), .B2(n40326), .C1(
        n40317), .C2(n32627), .ZN(n9039) );
  OAI222_X1 U33103 ( .A1(n40720), .A2(n40333), .B1(n41104), .B2(n40326), .C1(
        n40317), .C2(n32626), .ZN(n9038) );
  OAI222_X1 U33104 ( .A1(n40726), .A2(n40333), .B1(n41110), .B2(n40326), .C1(
        n40317), .C2(n32625), .ZN(n9037) );
  OAI222_X1 U33105 ( .A1(n40732), .A2(n40333), .B1(n41116), .B2(n40326), .C1(
        n40317), .C2(n32624), .ZN(n9036) );
  OAI222_X1 U33106 ( .A1(n40738), .A2(n40333), .B1(n41122), .B2(n40326), .C1(
        n40317), .C2(n32623), .ZN(n9035) );
  OAI222_X1 U33107 ( .A1(n40744), .A2(n40333), .B1(n41128), .B2(n40326), .C1(
        n40317), .C2(n32622), .ZN(n9034) );
  OAI222_X1 U33108 ( .A1(n40750), .A2(n40333), .B1(n41134), .B2(n40326), .C1(
        n40318), .C2(n32621), .ZN(n9033) );
  OAI222_X1 U33109 ( .A1(n40756), .A2(n40333), .B1(n41140), .B2(n40326), .C1(
        n40318), .C2(n32620), .ZN(n9032) );
  OAI222_X1 U33110 ( .A1(n40762), .A2(n40333), .B1(n41146), .B2(n40326), .C1(
        n40318), .C2(n32619), .ZN(n9031) );
  OAI222_X1 U33111 ( .A1(n40768), .A2(n40332), .B1(n41152), .B2(n40325), .C1(
        n40318), .C2(n32618), .ZN(n9030) );
  OAI222_X1 U33112 ( .A1(n40774), .A2(n40332), .B1(n41158), .B2(n40325), .C1(
        n40318), .C2(n32617), .ZN(n9029) );
  OAI222_X1 U33113 ( .A1(n40780), .A2(n40332), .B1(n41164), .B2(n40325), .C1(
        n40318), .C2(n32616), .ZN(n9028) );
  OAI222_X1 U33114 ( .A1(n40786), .A2(n40332), .B1(n41170), .B2(n40325), .C1(
        n40318), .C2(n32615), .ZN(n9027) );
  OAI222_X1 U33115 ( .A1(n40792), .A2(n40332), .B1(n41176), .B2(n40325), .C1(
        n40318), .C2(n32614), .ZN(n9026) );
  OAI222_X1 U33116 ( .A1(n40798), .A2(n40332), .B1(n41182), .B2(n40325), .C1(
        n40318), .C2(n32613), .ZN(n9025) );
  OAI222_X1 U33117 ( .A1(n40804), .A2(n40332), .B1(n41188), .B2(n40325), .C1(
        n40318), .C2(n32612), .ZN(n9024) );
  OAI222_X1 U33118 ( .A1(n40810), .A2(n40332), .B1(n41194), .B2(n40325), .C1(
        n40318), .C2(n32611), .ZN(n9023) );
  OAI222_X1 U33119 ( .A1(n40816), .A2(n40332), .B1(n41200), .B2(n40325), .C1(
        n40319), .C2(n32610), .ZN(n9022) );
  OAI222_X1 U33120 ( .A1(n40822), .A2(n40332), .B1(n41206), .B2(n40325), .C1(
        n40319), .C2(n32609), .ZN(n9021) );
  OAI222_X1 U33121 ( .A1(n40828), .A2(n40332), .B1(n41212), .B2(n40325), .C1(
        n40319), .C2(n32608), .ZN(n9020) );
  OAI222_X1 U33122 ( .A1(n40834), .A2(n40332), .B1(n41218), .B2(n40325), .C1(
        n40319), .C2(n32607), .ZN(n9019) );
  OAI222_X1 U33123 ( .A1(n40840), .A2(n40331), .B1(n41224), .B2(n40324), .C1(
        n40319), .C2(n32606), .ZN(n9018) );
  OAI222_X1 U33124 ( .A1(n40846), .A2(n40331), .B1(n41230), .B2(n40324), .C1(
        n40319), .C2(n32605), .ZN(n9017) );
  OAI222_X1 U33125 ( .A1(n40852), .A2(n40331), .B1(n41236), .B2(n40324), .C1(
        n40319), .C2(n32604), .ZN(n9016) );
  OAI222_X1 U33126 ( .A1(n40858), .A2(n40331), .B1(n41242), .B2(n40324), .C1(
        n40319), .C2(n32603), .ZN(n9015) );
  OAI222_X1 U33127 ( .A1(n40864), .A2(n40331), .B1(n41248), .B2(n40324), .C1(
        n40319), .C2(n32602), .ZN(n9014) );
  OAI222_X1 U33128 ( .A1(n40870), .A2(n40331), .B1(n41254), .B2(n40324), .C1(
        n40319), .C2(n32601), .ZN(n9013) );
  OAI222_X1 U33129 ( .A1(n40876), .A2(n40331), .B1(n41260), .B2(n40324), .C1(
        n40319), .C2(n32600), .ZN(n9012) );
  OAI222_X1 U33130 ( .A1(n40882), .A2(n40331), .B1(n41266), .B2(n40324), .C1(
        n40319), .C2(n32599), .ZN(n9011) );
  OAI222_X1 U33131 ( .A1(n40888), .A2(n40331), .B1(n41272), .B2(n40324), .C1(
        n40320), .C2(n32598), .ZN(n9010) );
  OAI222_X1 U33132 ( .A1(n40894), .A2(n40331), .B1(n41278), .B2(n40324), .C1(
        n40320), .C2(n32597), .ZN(n9009) );
  OAI222_X1 U33133 ( .A1(n40900), .A2(n40331), .B1(n41284), .B2(n40324), .C1(
        n40320), .C2(n32596), .ZN(n9008) );
  OAI222_X1 U33134 ( .A1(n40906), .A2(n40331), .B1(n41290), .B2(n40324), .C1(
        n40320), .C2(n32595), .ZN(n9007) );
  OAI222_X1 U33135 ( .A1(n40622), .A2(n39839), .B1(n41006), .B2(n39832), .C1(
        n39821), .C2(n32594), .ZN(n7454) );
  OAI222_X1 U33136 ( .A1(n40628), .A2(n39839), .B1(n41012), .B2(n39832), .C1(
        n39821), .C2(n32593), .ZN(n7453) );
  OAI222_X1 U33137 ( .A1(n40634), .A2(n39839), .B1(n41018), .B2(n39832), .C1(
        n39821), .C2(n32592), .ZN(n7452) );
  OAI222_X1 U33138 ( .A1(n40640), .A2(n39839), .B1(n41024), .B2(n39832), .C1(
        n39821), .C2(n32591), .ZN(n7451) );
  OAI222_X1 U33139 ( .A1(n40646), .A2(n39839), .B1(n41030), .B2(n39832), .C1(
        n39821), .C2(n32590), .ZN(n7450) );
  OAI222_X1 U33140 ( .A1(n40652), .A2(n39839), .B1(n41036), .B2(n39832), .C1(
        n39821), .C2(n32589), .ZN(n7449) );
  OAI222_X1 U33141 ( .A1(n40658), .A2(n39839), .B1(n41042), .B2(n39832), .C1(
        n39821), .C2(n32588), .ZN(n7448) );
  OAI222_X1 U33142 ( .A1(n40664), .A2(n39839), .B1(n41048), .B2(n39832), .C1(
        n39821), .C2(n32587), .ZN(n7447) );
  OAI222_X1 U33143 ( .A1(n40670), .A2(n39839), .B1(n41054), .B2(n39832), .C1(
        n39822), .C2(n32586), .ZN(n7446) );
  OAI222_X1 U33144 ( .A1(n40676), .A2(n39839), .B1(n41060), .B2(n39832), .C1(
        n39822), .C2(n32585), .ZN(n7445) );
  OAI222_X1 U33145 ( .A1(n40682), .A2(n39839), .B1(n41066), .B2(n39832), .C1(
        n39822), .C2(n32584), .ZN(n7444) );
  OAI222_X1 U33146 ( .A1(n40688), .A2(n39839), .B1(n41072), .B2(n39832), .C1(
        n39823), .C2(n32583), .ZN(n7443) );
  OAI222_X1 U33147 ( .A1(n40694), .A2(n39838), .B1(n41078), .B2(n39831), .C1(
        n39822), .C2(n32582), .ZN(n7442) );
  OAI222_X1 U33148 ( .A1(n40700), .A2(n39838), .B1(n41084), .B2(n39831), .C1(
        n39822), .C2(n32581), .ZN(n7441) );
  OAI222_X1 U33149 ( .A1(n40706), .A2(n39838), .B1(n41090), .B2(n39831), .C1(
        n39822), .C2(n32580), .ZN(n7440) );
  OAI222_X1 U33150 ( .A1(n40712), .A2(n39838), .B1(n41096), .B2(n39831), .C1(
        n39822), .C2(n32579), .ZN(n7439) );
  OAI222_X1 U33151 ( .A1(n40718), .A2(n39838), .B1(n41102), .B2(n39831), .C1(
        n39822), .C2(n32578), .ZN(n7438) );
  OAI222_X1 U33152 ( .A1(n40724), .A2(n39838), .B1(n41108), .B2(n39831), .C1(
        n39822), .C2(n32577), .ZN(n7437) );
  OAI222_X1 U33153 ( .A1(n40730), .A2(n39838), .B1(n41114), .B2(n39831), .C1(
        n39822), .C2(n32576), .ZN(n7436) );
  OAI222_X1 U33154 ( .A1(n40736), .A2(n39838), .B1(n41120), .B2(n39831), .C1(
        n39822), .C2(n32575), .ZN(n7435) );
  OAI222_X1 U33155 ( .A1(n40742), .A2(n39838), .B1(n41126), .B2(n39831), .C1(
        n39822), .C2(n32574), .ZN(n7434) );
  OAI222_X1 U33156 ( .A1(n40748), .A2(n39838), .B1(n41132), .B2(n39831), .C1(
        n39823), .C2(n32573), .ZN(n7433) );
  OAI222_X1 U33157 ( .A1(n40754), .A2(n39838), .B1(n41138), .B2(n39831), .C1(
        n39823), .C2(n32572), .ZN(n7432) );
  OAI222_X1 U33158 ( .A1(n40760), .A2(n39838), .B1(n41144), .B2(n39831), .C1(
        n39823), .C2(n32571), .ZN(n7431) );
  OAI222_X1 U33159 ( .A1(n40766), .A2(n39837), .B1(n41150), .B2(n39830), .C1(
        n39823), .C2(n32570), .ZN(n7430) );
  OAI222_X1 U33160 ( .A1(n40772), .A2(n39837), .B1(n41156), .B2(n39830), .C1(
        n39823), .C2(n32569), .ZN(n7429) );
  OAI222_X1 U33161 ( .A1(n40778), .A2(n39837), .B1(n41162), .B2(n39830), .C1(
        n39823), .C2(n32568), .ZN(n7428) );
  OAI222_X1 U33162 ( .A1(n40784), .A2(n39837), .B1(n41168), .B2(n39830), .C1(
        n39823), .C2(n32567), .ZN(n7427) );
  OAI222_X1 U33163 ( .A1(n40790), .A2(n39837), .B1(n41174), .B2(n39830), .C1(
        n39823), .C2(n32566), .ZN(n7426) );
  OAI222_X1 U33164 ( .A1(n40796), .A2(n39837), .B1(n41180), .B2(n39830), .C1(
        n39823), .C2(n32565), .ZN(n7425) );
  OAI222_X1 U33165 ( .A1(n40802), .A2(n39837), .B1(n41186), .B2(n39830), .C1(
        n39823), .C2(n32564), .ZN(n7424) );
  OAI222_X1 U33166 ( .A1(n40808), .A2(n39837), .B1(n41192), .B2(n39830), .C1(
        n39823), .C2(n32563), .ZN(n7423) );
  OAI222_X1 U33167 ( .A1(n40814), .A2(n39837), .B1(n41198), .B2(n39830), .C1(
        n39824), .C2(n32562), .ZN(n7422) );
  OAI222_X1 U33168 ( .A1(n40820), .A2(n39837), .B1(n41204), .B2(n39830), .C1(
        n39824), .C2(n32561), .ZN(n7421) );
  OAI222_X1 U33169 ( .A1(n40826), .A2(n39837), .B1(n41210), .B2(n39830), .C1(
        n39824), .C2(n32560), .ZN(n7420) );
  OAI222_X1 U33170 ( .A1(n40832), .A2(n39837), .B1(n41216), .B2(n39830), .C1(
        n39824), .C2(n32559), .ZN(n7419) );
  OAI222_X1 U33171 ( .A1(n40838), .A2(n39836), .B1(n41222), .B2(n39829), .C1(
        n39824), .C2(n32558), .ZN(n7418) );
  OAI222_X1 U33172 ( .A1(n40844), .A2(n39836), .B1(n41228), .B2(n39829), .C1(
        n39824), .C2(n32557), .ZN(n7417) );
  OAI222_X1 U33173 ( .A1(n40850), .A2(n39836), .B1(n41234), .B2(n39829), .C1(
        n39824), .C2(n32556), .ZN(n7416) );
  OAI222_X1 U33174 ( .A1(n40856), .A2(n39836), .B1(n41240), .B2(n39829), .C1(
        n39824), .C2(n32555), .ZN(n7415) );
  OAI222_X1 U33175 ( .A1(n40862), .A2(n39836), .B1(n41246), .B2(n39829), .C1(
        n39824), .C2(n32554), .ZN(n7414) );
  OAI222_X1 U33176 ( .A1(n40868), .A2(n39836), .B1(n41252), .B2(n39829), .C1(
        n39824), .C2(n32553), .ZN(n7413) );
  OAI222_X1 U33177 ( .A1(n40874), .A2(n39836), .B1(n41258), .B2(n39829), .C1(
        n39824), .C2(n32552), .ZN(n7412) );
  OAI222_X1 U33178 ( .A1(n40880), .A2(n39836), .B1(n41264), .B2(n39829), .C1(
        n39824), .C2(n32551), .ZN(n7411) );
  OAI222_X1 U33179 ( .A1(n40886), .A2(n39836), .B1(n41270), .B2(n39829), .C1(
        n39825), .C2(n32550), .ZN(n7410) );
  OAI222_X1 U33180 ( .A1(n40892), .A2(n39836), .B1(n41276), .B2(n39829), .C1(
        n39825), .C2(n32549), .ZN(n7409) );
  OAI222_X1 U33181 ( .A1(n40898), .A2(n39836), .B1(n41282), .B2(n39829), .C1(
        n39825), .C2(n32548), .ZN(n7408) );
  OAI222_X1 U33182 ( .A1(n40904), .A2(n39836), .B1(n41288), .B2(n39829), .C1(
        n39825), .C2(n32547), .ZN(n7407) );
  OAI222_X1 U33183 ( .A1(n40635), .A2(n40134), .B1(n41019), .B2(n40127), .C1(
        n40116), .C2(n38850), .ZN(n8412) );
  OAI222_X1 U33184 ( .A1(n40623), .A2(n40134), .B1(n41007), .B2(n40127), .C1(
        n40116), .C2(n38851), .ZN(n8414) );
  OAI222_X1 U33185 ( .A1(n40629), .A2(n40134), .B1(n41013), .B2(n40127), .C1(
        n40116), .C2(n38852), .ZN(n8413) );
  OAI222_X1 U33186 ( .A1(n40641), .A2(n40134), .B1(n41025), .B2(n40127), .C1(
        n40116), .C2(n38853), .ZN(n8411) );
  OAI222_X1 U33187 ( .A1(n40647), .A2(n40134), .B1(n41031), .B2(n40127), .C1(
        n40116), .C2(n38854), .ZN(n8410) );
  OAI222_X1 U33188 ( .A1(n40653), .A2(n40134), .B1(n41037), .B2(n40127), .C1(
        n40116), .C2(n38855), .ZN(n8409) );
  OAI222_X1 U33189 ( .A1(n40600), .A2(n40435), .B1(n40984), .B2(n40428), .C1(
        n40416), .C2(n38856), .ZN(n9378) );
  OAI222_X1 U33190 ( .A1(n40606), .A2(n40435), .B1(n40990), .B2(n40428), .C1(
        n40416), .C2(n38857), .ZN(n9377) );
  OAI222_X1 U33191 ( .A1(n40612), .A2(n40435), .B1(n40996), .B2(n40428), .C1(
        n40416), .C2(n38858), .ZN(n9376) );
  OAI222_X1 U33192 ( .A1(n40618), .A2(n40435), .B1(n41002), .B2(n40428), .C1(
        n40416), .C2(n38859), .ZN(n9375) );
  OAI222_X1 U33193 ( .A1(n40600), .A2(n40415), .B1(n40984), .B2(n40408), .C1(
        n40396), .C2(n38983), .ZN(n9314) );
  OAI222_X1 U33194 ( .A1(n40606), .A2(n40415), .B1(n40990), .B2(n40408), .C1(
        n40396), .C2(n38984), .ZN(n9313) );
  OAI222_X1 U33195 ( .A1(n40612), .A2(n40415), .B1(n40996), .B2(n40408), .C1(
        n40396), .C2(n38985), .ZN(n9312) );
  OAI222_X1 U33196 ( .A1(n40618), .A2(n40415), .B1(n41002), .B2(n40408), .C1(
        n40396), .C2(n38986), .ZN(n9311) );
  OAI222_X1 U33197 ( .A1(n40599), .A2(n40215), .B1(n40983), .B2(n40208), .C1(
        n40196), .C2(n32483), .ZN(n8674) );
  OAI222_X1 U33198 ( .A1(n40605), .A2(n40215), .B1(n40989), .B2(n40208), .C1(
        n40196), .C2(n32482), .ZN(n8673) );
  OAI222_X1 U33199 ( .A1(n40611), .A2(n40215), .B1(n40995), .B2(n40208), .C1(
        n40196), .C2(n32481), .ZN(n8672) );
  OAI222_X1 U33200 ( .A1(n40617), .A2(n40215), .B1(n41001), .B2(n40208), .C1(
        n40196), .C2(n32480), .ZN(n8671) );
  OAI222_X1 U33201 ( .A1(n40599), .A2(n40235), .B1(n40983), .B2(n40228), .C1(
        n40216), .C2(n32479), .ZN(n8738) );
  OAI222_X1 U33202 ( .A1(n40605), .A2(n40235), .B1(n40989), .B2(n40228), .C1(
        n40216), .C2(n32478), .ZN(n8737) );
  OAI222_X1 U33203 ( .A1(n40611), .A2(n40235), .B1(n40995), .B2(n40228), .C1(
        n40216), .C2(n32477), .ZN(n8736) );
  OAI222_X1 U33204 ( .A1(n40617), .A2(n40235), .B1(n41001), .B2(n40228), .C1(
        n40216), .C2(n32476), .ZN(n8735) );
  OAI222_X1 U33205 ( .A1(n40600), .A2(n40315), .B1(n40984), .B2(n40308), .C1(
        n40296), .C2(n32467), .ZN(n8994) );
  OAI222_X1 U33206 ( .A1(n40606), .A2(n40315), .B1(n40990), .B2(n40308), .C1(
        n40296), .C2(n32466), .ZN(n8993) );
  OAI222_X1 U33207 ( .A1(n40612), .A2(n40315), .B1(n40996), .B2(n40308), .C1(
        n40296), .C2(n32465), .ZN(n8992) );
  OAI222_X1 U33208 ( .A1(n40618), .A2(n40315), .B1(n41002), .B2(n40308), .C1(
        n40296), .C2(n32464), .ZN(n8991) );
  OAI222_X1 U33209 ( .A1(n40600), .A2(n40335), .B1(n40984), .B2(n40328), .C1(
        n40316), .C2(n32463), .ZN(n9058) );
  OAI222_X1 U33210 ( .A1(n40606), .A2(n40335), .B1(n40990), .B2(n40328), .C1(
        n40316), .C2(n32462), .ZN(n9057) );
  OAI222_X1 U33211 ( .A1(n40612), .A2(n40335), .B1(n40996), .B2(n40328), .C1(
        n40316), .C2(n32461), .ZN(n9056) );
  OAI222_X1 U33212 ( .A1(n40618), .A2(n40335), .B1(n41002), .B2(n40328), .C1(
        n40316), .C2(n32460), .ZN(n9055) );
  OAI222_X1 U33213 ( .A1(n40598), .A2(n39840), .B1(n40982), .B2(n39833), .C1(
        n39821), .C2(n32459), .ZN(n7458) );
  OAI222_X1 U33214 ( .A1(n40604), .A2(n39840), .B1(n40988), .B2(n39833), .C1(
        n39821), .C2(n32458), .ZN(n7457) );
  OAI222_X1 U33215 ( .A1(n40610), .A2(n39840), .B1(n40994), .B2(n39833), .C1(
        n39821), .C2(n32457), .ZN(n7456) );
  OAI222_X1 U33216 ( .A1(n40616), .A2(n39840), .B1(n41000), .B2(n39833), .C1(
        n39821), .C2(n32456), .ZN(n7455) );
  OAI222_X1 U33217 ( .A1(n40599), .A2(n40135), .B1(n40983), .B2(n40128), .C1(
        n40116), .C2(n38860), .ZN(n8418) );
  OAI222_X1 U33218 ( .A1(n40605), .A2(n40135), .B1(n40989), .B2(n40128), .C1(
        n40116), .C2(n38861), .ZN(n8417) );
  OAI222_X1 U33219 ( .A1(n40611), .A2(n40135), .B1(n40995), .B2(n40128), .C1(
        n40116), .C2(n38862), .ZN(n8416) );
  OAI222_X1 U33220 ( .A1(n40617), .A2(n40135), .B1(n41001), .B2(n40128), .C1(
        n40116), .C2(n38863), .ZN(n8415) );
  OAI222_X1 U33221 ( .A1(n40913), .A2(n40530), .B1(n41297), .B2(n40523), .C1(
        n40520), .C2(n38864), .ZN(n9646) );
  OAI222_X1 U33222 ( .A1(n40919), .A2(n40530), .B1(n41303), .B2(n40523), .C1(
        n40520), .C2(n38865), .ZN(n9645) );
  OAI222_X1 U33223 ( .A1(n40925), .A2(n40530), .B1(n41309), .B2(n40523), .C1(
        n40520), .C2(n38866), .ZN(n9644) );
  OAI222_X1 U33224 ( .A1(n40931), .A2(n40530), .B1(n41315), .B2(n40523), .C1(
        n40520), .C2(n38867), .ZN(n9643) );
  OAI222_X1 U33225 ( .A1(n40937), .A2(n40530), .B1(n41321), .B2(n40523), .C1(
        n40520), .C2(n38868), .ZN(n9642) );
  OAI222_X1 U33226 ( .A1(n40943), .A2(n40530), .B1(n41327), .B2(n40523), .C1(
        n40520), .C2(n38869), .ZN(n9641) );
  OAI222_X1 U33227 ( .A1(n40949), .A2(n40530), .B1(n41333), .B2(n40523), .C1(
        n40520), .C2(n38870), .ZN(n9640) );
  OAI222_X1 U33228 ( .A1(n40961), .A2(n40530), .B1(n41345), .B2(n40523), .C1(
        n40520), .C2(n38871), .ZN(n9638) );
  OAI222_X1 U33229 ( .A1(n40625), .A2(n40534), .B1(n41009), .B2(n40527), .C1(
        n40516), .C2(n38872), .ZN(n9694) );
  OAI222_X1 U33230 ( .A1(n40631), .A2(n40534), .B1(n41015), .B2(n40527), .C1(
        n40516), .C2(n38873), .ZN(n9693) );
  OAI222_X1 U33231 ( .A1(n40637), .A2(n40534), .B1(n41021), .B2(n40527), .C1(
        n40516), .C2(n38874), .ZN(n9692) );
  OAI222_X1 U33232 ( .A1(n40643), .A2(n40534), .B1(n41027), .B2(n40527), .C1(
        n40516), .C2(n38875), .ZN(n9691) );
  OAI222_X1 U33233 ( .A1(n40649), .A2(n40534), .B1(n41033), .B2(n40527), .C1(
        n40516), .C2(n38876), .ZN(n9690) );
  OAI222_X1 U33234 ( .A1(n40655), .A2(n40534), .B1(n41039), .B2(n40527), .C1(
        n40516), .C2(n38877), .ZN(n9689) );
  OAI222_X1 U33235 ( .A1(n40661), .A2(n40534), .B1(n41045), .B2(n40527), .C1(
        n40516), .C2(n38878), .ZN(n9688) );
  OAI222_X1 U33236 ( .A1(n40667), .A2(n40534), .B1(n41051), .B2(n40527), .C1(
        n40516), .C2(n38879), .ZN(n9687) );
  OAI222_X1 U33237 ( .A1(n40673), .A2(n40534), .B1(n41057), .B2(n40527), .C1(
        n40517), .C2(n38880), .ZN(n9686) );
  OAI222_X1 U33238 ( .A1(n40679), .A2(n40534), .B1(n41063), .B2(n40527), .C1(
        n40517), .C2(n38881), .ZN(n9685) );
  OAI222_X1 U33239 ( .A1(n40685), .A2(n40534), .B1(n41069), .B2(n40527), .C1(
        n40517), .C2(n38882), .ZN(n9684) );
  OAI222_X1 U33240 ( .A1(n40691), .A2(n40534), .B1(n41075), .B2(n40527), .C1(
        n40518), .C2(n38883), .ZN(n9683) );
  OAI222_X1 U33241 ( .A1(n40697), .A2(n40533), .B1(n41081), .B2(n40526), .C1(
        n40517), .C2(n38884), .ZN(n9682) );
  OAI222_X1 U33242 ( .A1(n40703), .A2(n40533), .B1(n41087), .B2(n40526), .C1(
        n40517), .C2(n38885), .ZN(n9681) );
  OAI222_X1 U33243 ( .A1(n40709), .A2(n40533), .B1(n41093), .B2(n40526), .C1(
        n40517), .C2(n38886), .ZN(n9680) );
  OAI222_X1 U33244 ( .A1(n40715), .A2(n40533), .B1(n41099), .B2(n40526), .C1(
        n40517), .C2(n38887), .ZN(n9679) );
  OAI222_X1 U33245 ( .A1(n40721), .A2(n40533), .B1(n41105), .B2(n40526), .C1(
        n40517), .C2(n38888), .ZN(n9678) );
  OAI222_X1 U33246 ( .A1(n40727), .A2(n40533), .B1(n41111), .B2(n40526), .C1(
        n40517), .C2(n38889), .ZN(n9677) );
  OAI222_X1 U33247 ( .A1(n40733), .A2(n40533), .B1(n41117), .B2(n40526), .C1(
        n40517), .C2(n38890), .ZN(n9676) );
  OAI222_X1 U33248 ( .A1(n40739), .A2(n40533), .B1(n41123), .B2(n40526), .C1(
        n40517), .C2(n38891), .ZN(n9675) );
  OAI222_X1 U33249 ( .A1(n40745), .A2(n40533), .B1(n41129), .B2(n40526), .C1(
        n40517), .C2(n38892), .ZN(n9674) );
  OAI222_X1 U33250 ( .A1(n40751), .A2(n40533), .B1(n41135), .B2(n40526), .C1(
        n40518), .C2(n38893), .ZN(n9673) );
  OAI222_X1 U33251 ( .A1(n40757), .A2(n40533), .B1(n41141), .B2(n40526), .C1(
        n40518), .C2(n38894), .ZN(n9672) );
  OAI222_X1 U33252 ( .A1(n40763), .A2(n40533), .B1(n41147), .B2(n40526), .C1(
        n40518), .C2(n38895), .ZN(n9671) );
  OAI222_X1 U33253 ( .A1(n40769), .A2(n40532), .B1(n41153), .B2(n40525), .C1(
        n40518), .C2(n38896), .ZN(n9670) );
  OAI222_X1 U33254 ( .A1(n40775), .A2(n40532), .B1(n41159), .B2(n40525), .C1(
        n40518), .C2(n38897), .ZN(n9669) );
  OAI222_X1 U33255 ( .A1(n40781), .A2(n40532), .B1(n41165), .B2(n40525), .C1(
        n40518), .C2(n38898), .ZN(n9668) );
  OAI222_X1 U33256 ( .A1(n40787), .A2(n40532), .B1(n41171), .B2(n40525), .C1(
        n40518), .C2(n38899), .ZN(n9667) );
  OAI222_X1 U33257 ( .A1(n40793), .A2(n40532), .B1(n41177), .B2(n40525), .C1(
        n40518), .C2(n38900), .ZN(n9666) );
  OAI222_X1 U33258 ( .A1(n40799), .A2(n40532), .B1(n41183), .B2(n40525), .C1(
        n40518), .C2(n38901), .ZN(n9665) );
  OAI222_X1 U33259 ( .A1(n40805), .A2(n40532), .B1(n41189), .B2(n40525), .C1(
        n40518), .C2(n38902), .ZN(n9664) );
  OAI222_X1 U33260 ( .A1(n40811), .A2(n40532), .B1(n41195), .B2(n40525), .C1(
        n40518), .C2(n38903), .ZN(n9663) );
  OAI222_X1 U33261 ( .A1(n40817), .A2(n40532), .B1(n41201), .B2(n40525), .C1(
        n40519), .C2(n38904), .ZN(n9662) );
  OAI222_X1 U33262 ( .A1(n40823), .A2(n40532), .B1(n41207), .B2(n40525), .C1(
        n40519), .C2(n38905), .ZN(n9661) );
  OAI222_X1 U33263 ( .A1(n40829), .A2(n40532), .B1(n41213), .B2(n40525), .C1(
        n40519), .C2(n38906), .ZN(n9660) );
  OAI222_X1 U33264 ( .A1(n40835), .A2(n40532), .B1(n41219), .B2(n40525), .C1(
        n40519), .C2(n38907), .ZN(n9659) );
  OAI222_X1 U33265 ( .A1(n40841), .A2(n40531), .B1(n41225), .B2(n40524), .C1(
        n40519), .C2(n38908), .ZN(n9658) );
  OAI222_X1 U33266 ( .A1(n40847), .A2(n40531), .B1(n41231), .B2(n40524), .C1(
        n40519), .C2(n38909), .ZN(n9657) );
  OAI222_X1 U33267 ( .A1(n40853), .A2(n40531), .B1(n41237), .B2(n40524), .C1(
        n40519), .C2(n38910), .ZN(n9656) );
  OAI222_X1 U33268 ( .A1(n40859), .A2(n40531), .B1(n41243), .B2(n40524), .C1(
        n40519), .C2(n38911), .ZN(n9655) );
  OAI222_X1 U33269 ( .A1(n40865), .A2(n40531), .B1(n41249), .B2(n40524), .C1(
        n40519), .C2(n38912), .ZN(n9654) );
  OAI222_X1 U33270 ( .A1(n40871), .A2(n40531), .B1(n41255), .B2(n40524), .C1(
        n40519), .C2(n38913), .ZN(n9653) );
  OAI222_X1 U33271 ( .A1(n40877), .A2(n40531), .B1(n41261), .B2(n40524), .C1(
        n40519), .C2(n38914), .ZN(n9652) );
  OAI222_X1 U33272 ( .A1(n40883), .A2(n40531), .B1(n41267), .B2(n40524), .C1(
        n40519), .C2(n38915), .ZN(n9651) );
  OAI222_X1 U33273 ( .A1(n40889), .A2(n40531), .B1(n41273), .B2(n40524), .C1(
        n40520), .C2(n38916), .ZN(n9650) );
  OAI222_X1 U33274 ( .A1(n40895), .A2(n40531), .B1(n41279), .B2(n40524), .C1(
        n40520), .C2(n38917), .ZN(n9649) );
  OAI222_X1 U33275 ( .A1(n40901), .A2(n40531), .B1(n41285), .B2(n40524), .C1(
        n40520), .C2(n38918), .ZN(n9648) );
  OAI222_X1 U33276 ( .A1(n40907), .A2(n40531), .B1(n41291), .B2(n40524), .C1(
        n40520), .C2(n38919), .ZN(n9647) );
  OAI222_X1 U33277 ( .A1(n40912), .A2(n40510), .B1(n41296), .B2(n40503), .C1(
        n40500), .C2(n38987), .ZN(n9582) );
  OAI222_X1 U33278 ( .A1(n40918), .A2(n40510), .B1(n41302), .B2(n40503), .C1(
        n40500), .C2(n38988), .ZN(n9581) );
  OAI222_X1 U33279 ( .A1(n40924), .A2(n40510), .B1(n41308), .B2(n40503), .C1(
        n40500), .C2(n38989), .ZN(n9580) );
  OAI222_X1 U33280 ( .A1(n40930), .A2(n40510), .B1(n41314), .B2(n40503), .C1(
        n40500), .C2(n38990), .ZN(n9579) );
  OAI222_X1 U33281 ( .A1(n40936), .A2(n40510), .B1(n41320), .B2(n40503), .C1(
        n40500), .C2(n38991), .ZN(n9578) );
  OAI222_X1 U33282 ( .A1(n40942), .A2(n40510), .B1(n41326), .B2(n40503), .C1(
        n40500), .C2(n38992), .ZN(n9577) );
  OAI222_X1 U33283 ( .A1(n40948), .A2(n40510), .B1(n41332), .B2(n40503), .C1(
        n40500), .C2(n38993), .ZN(n9576) );
  OAI222_X1 U33284 ( .A1(n40960), .A2(n40510), .B1(n41344), .B2(n40503), .C1(
        n40500), .C2(n38994), .ZN(n9574) );
  OAI222_X1 U33285 ( .A1(n40624), .A2(n40514), .B1(n41008), .B2(n40507), .C1(
        n40496), .C2(n38995), .ZN(n9630) );
  OAI222_X1 U33286 ( .A1(n40630), .A2(n40514), .B1(n41014), .B2(n40507), .C1(
        n40496), .C2(n38996), .ZN(n9629) );
  OAI222_X1 U33287 ( .A1(n40636), .A2(n40514), .B1(n41020), .B2(n40507), .C1(
        n40496), .C2(n38997), .ZN(n9628) );
  OAI222_X1 U33288 ( .A1(n40642), .A2(n40514), .B1(n41026), .B2(n40507), .C1(
        n40496), .C2(n38998), .ZN(n9627) );
  OAI222_X1 U33289 ( .A1(n40648), .A2(n40514), .B1(n41032), .B2(n40507), .C1(
        n40496), .C2(n38999), .ZN(n9626) );
  OAI222_X1 U33290 ( .A1(n40654), .A2(n40514), .B1(n41038), .B2(n40507), .C1(
        n40496), .C2(n39000), .ZN(n9625) );
  OAI222_X1 U33291 ( .A1(n40660), .A2(n40514), .B1(n41044), .B2(n40507), .C1(
        n40496), .C2(n39001), .ZN(n9624) );
  OAI222_X1 U33292 ( .A1(n40666), .A2(n40514), .B1(n41050), .B2(n40507), .C1(
        n40496), .C2(n39002), .ZN(n9623) );
  OAI222_X1 U33293 ( .A1(n40672), .A2(n40514), .B1(n41056), .B2(n40507), .C1(
        n40497), .C2(n39003), .ZN(n9622) );
  OAI222_X1 U33294 ( .A1(n40678), .A2(n40514), .B1(n41062), .B2(n40507), .C1(
        n40497), .C2(n39004), .ZN(n9621) );
  OAI222_X1 U33295 ( .A1(n40684), .A2(n40514), .B1(n41068), .B2(n40507), .C1(
        n40497), .C2(n39005), .ZN(n9620) );
  OAI222_X1 U33296 ( .A1(n40690), .A2(n40514), .B1(n41074), .B2(n40507), .C1(
        n40498), .C2(n39006), .ZN(n9619) );
  OAI222_X1 U33297 ( .A1(n40696), .A2(n40513), .B1(n41080), .B2(n40506), .C1(
        n40497), .C2(n39007), .ZN(n9618) );
  OAI222_X1 U33298 ( .A1(n40702), .A2(n40513), .B1(n41086), .B2(n40506), .C1(
        n40497), .C2(n39008), .ZN(n9617) );
  OAI222_X1 U33299 ( .A1(n40708), .A2(n40513), .B1(n41092), .B2(n40506), .C1(
        n40497), .C2(n39009), .ZN(n9616) );
  OAI222_X1 U33300 ( .A1(n40714), .A2(n40513), .B1(n41098), .B2(n40506), .C1(
        n40497), .C2(n39010), .ZN(n9615) );
  OAI222_X1 U33301 ( .A1(n40720), .A2(n40513), .B1(n41104), .B2(n40506), .C1(
        n40497), .C2(n39011), .ZN(n9614) );
  OAI222_X1 U33302 ( .A1(n40726), .A2(n40513), .B1(n41110), .B2(n40506), .C1(
        n40497), .C2(n39012), .ZN(n9613) );
  OAI222_X1 U33303 ( .A1(n40732), .A2(n40513), .B1(n41116), .B2(n40506), .C1(
        n40497), .C2(n39013), .ZN(n9612) );
  OAI222_X1 U33304 ( .A1(n40738), .A2(n40513), .B1(n41122), .B2(n40506), .C1(
        n40497), .C2(n39014), .ZN(n9611) );
  OAI222_X1 U33305 ( .A1(n40744), .A2(n40513), .B1(n41128), .B2(n40506), .C1(
        n40497), .C2(n39015), .ZN(n9610) );
  OAI222_X1 U33306 ( .A1(n40750), .A2(n40513), .B1(n41134), .B2(n40506), .C1(
        n40498), .C2(n39016), .ZN(n9609) );
  OAI222_X1 U33307 ( .A1(n40756), .A2(n40513), .B1(n41140), .B2(n40506), .C1(
        n40498), .C2(n39017), .ZN(n9608) );
  OAI222_X1 U33308 ( .A1(n40762), .A2(n40513), .B1(n41146), .B2(n40506), .C1(
        n40498), .C2(n39018), .ZN(n9607) );
  OAI222_X1 U33309 ( .A1(n40768), .A2(n40512), .B1(n41152), .B2(n40505), .C1(
        n40498), .C2(n39019), .ZN(n9606) );
  OAI222_X1 U33310 ( .A1(n40774), .A2(n40512), .B1(n41158), .B2(n40505), .C1(
        n40498), .C2(n39020), .ZN(n9605) );
  OAI222_X1 U33311 ( .A1(n40780), .A2(n40512), .B1(n41164), .B2(n40505), .C1(
        n40498), .C2(n39021), .ZN(n9604) );
  OAI222_X1 U33312 ( .A1(n40786), .A2(n40512), .B1(n41170), .B2(n40505), .C1(
        n40498), .C2(n39022), .ZN(n9603) );
  OAI222_X1 U33313 ( .A1(n40792), .A2(n40512), .B1(n41176), .B2(n40505), .C1(
        n40498), .C2(n39023), .ZN(n9602) );
  OAI222_X1 U33314 ( .A1(n40798), .A2(n40512), .B1(n41182), .B2(n40505), .C1(
        n40498), .C2(n39024), .ZN(n9601) );
  OAI222_X1 U33315 ( .A1(n40804), .A2(n40512), .B1(n41188), .B2(n40505), .C1(
        n40498), .C2(n39025), .ZN(n9600) );
  OAI222_X1 U33316 ( .A1(n40810), .A2(n40512), .B1(n41194), .B2(n40505), .C1(
        n40498), .C2(n39026), .ZN(n9599) );
  OAI222_X1 U33317 ( .A1(n40816), .A2(n40512), .B1(n41200), .B2(n40505), .C1(
        n40499), .C2(n39027), .ZN(n9598) );
  OAI222_X1 U33318 ( .A1(n40822), .A2(n40512), .B1(n41206), .B2(n40505), .C1(
        n40499), .C2(n39028), .ZN(n9597) );
  OAI222_X1 U33319 ( .A1(n40828), .A2(n40512), .B1(n41212), .B2(n40505), .C1(
        n40499), .C2(n39029), .ZN(n9596) );
  OAI222_X1 U33320 ( .A1(n40834), .A2(n40512), .B1(n41218), .B2(n40505), .C1(
        n40499), .C2(n39030), .ZN(n9595) );
  OAI222_X1 U33321 ( .A1(n40840), .A2(n40511), .B1(n41224), .B2(n40504), .C1(
        n40499), .C2(n39031), .ZN(n9594) );
  OAI222_X1 U33322 ( .A1(n40846), .A2(n40511), .B1(n41230), .B2(n40504), .C1(
        n40499), .C2(n39032), .ZN(n9593) );
  OAI222_X1 U33323 ( .A1(n40852), .A2(n40511), .B1(n41236), .B2(n40504), .C1(
        n40499), .C2(n39033), .ZN(n9592) );
  OAI222_X1 U33324 ( .A1(n40858), .A2(n40511), .B1(n41242), .B2(n40504), .C1(
        n40499), .C2(n39034), .ZN(n9591) );
  OAI222_X1 U33325 ( .A1(n40864), .A2(n40511), .B1(n41248), .B2(n40504), .C1(
        n40499), .C2(n39035), .ZN(n9590) );
  OAI222_X1 U33326 ( .A1(n40870), .A2(n40511), .B1(n41254), .B2(n40504), .C1(
        n40499), .C2(n39036), .ZN(n9589) );
  OAI222_X1 U33327 ( .A1(n40876), .A2(n40511), .B1(n41260), .B2(n40504), .C1(
        n40499), .C2(n39037), .ZN(n9588) );
  OAI222_X1 U33328 ( .A1(n40882), .A2(n40511), .B1(n41266), .B2(n40504), .C1(
        n40499), .C2(n39038), .ZN(n9587) );
  OAI222_X1 U33329 ( .A1(n40888), .A2(n40511), .B1(n41272), .B2(n40504), .C1(
        n40500), .C2(n39039), .ZN(n9586) );
  OAI222_X1 U33330 ( .A1(n40894), .A2(n40511), .B1(n41278), .B2(n40504), .C1(
        n40500), .C2(n39040), .ZN(n9585) );
  OAI222_X1 U33331 ( .A1(n40900), .A2(n40511), .B1(n41284), .B2(n40504), .C1(
        n40500), .C2(n39041), .ZN(n9584) );
  OAI222_X1 U33332 ( .A1(n40906), .A2(n40511), .B1(n41290), .B2(n40504), .C1(
        n40500), .C2(n39042), .ZN(n9583) );
  OAI222_X1 U33333 ( .A1(n40601), .A2(n40535), .B1(n40985), .B2(n40528), .C1(
        n40516), .C2(n38920), .ZN(n9698) );
  OAI222_X1 U33334 ( .A1(n40607), .A2(n40535), .B1(n40991), .B2(n40528), .C1(
        n40516), .C2(n38921), .ZN(n9697) );
  OAI222_X1 U33335 ( .A1(n40613), .A2(n40535), .B1(n40997), .B2(n40528), .C1(
        n40516), .C2(n38922), .ZN(n9696) );
  OAI222_X1 U33336 ( .A1(n40619), .A2(n40535), .B1(n41003), .B2(n40528), .C1(
        n40516), .C2(n38923), .ZN(n9695) );
  OAI222_X1 U33337 ( .A1(n40600), .A2(n40515), .B1(n40984), .B2(n40508), .C1(
        n40496), .C2(n39043), .ZN(n9634) );
  OAI222_X1 U33338 ( .A1(n40606), .A2(n40515), .B1(n40990), .B2(n40508), .C1(
        n40496), .C2(n39044), .ZN(n9633) );
  OAI222_X1 U33339 ( .A1(n40612), .A2(n40515), .B1(n40996), .B2(n40508), .C1(
        n40496), .C2(n39045), .ZN(n9632) );
  OAI222_X1 U33340 ( .A1(n40618), .A2(n40515), .B1(n41002), .B2(n40508), .C1(
        n40496), .C2(n39046), .ZN(n9631) );
  AOI221_X1 U33341 ( .B1(n39222), .B2(n29415), .C1(n39216), .C2(n29479), .A(
        n37018), .ZN(n37013) );
  OAI222_X1 U33342 ( .A1(n31675), .A2(n39210), .B1(n31739), .B2(n39204), .C1(
        n31611), .C2(n39198), .ZN(n37018) );
  AOI221_X1 U33343 ( .B1(n39223), .B2(n29414), .C1(n39217), .C2(n29478), .A(
        n36999), .ZN(n36994) );
  OAI222_X1 U33344 ( .A1(n31674), .A2(n39211), .B1(n31738), .B2(n39205), .C1(
        n31610), .C2(n39199), .ZN(n36999) );
  AOI221_X1 U33345 ( .B1(n39223), .B2(n29413), .C1(n39217), .C2(n29477), .A(
        n36980), .ZN(n36975) );
  OAI222_X1 U33346 ( .A1(n31673), .A2(n39211), .B1(n31737), .B2(n39205), .C1(
        n31609), .C2(n39199), .ZN(n36980) );
  AOI221_X1 U33347 ( .B1(n39223), .B2(n29412), .C1(n39217), .C2(n29476), .A(
        n36961), .ZN(n36956) );
  OAI222_X1 U33348 ( .A1(n31672), .A2(n39211), .B1(n31736), .B2(n39205), .C1(
        n31608), .C2(n39199), .ZN(n36961) );
  AOI221_X1 U33349 ( .B1(n39223), .B2(n29411), .C1(n39217), .C2(n29475), .A(
        n36942), .ZN(n36937) );
  OAI222_X1 U33350 ( .A1(n31671), .A2(n39211), .B1(n31735), .B2(n39205), .C1(
        n31607), .C2(n39199), .ZN(n36942) );
  AOI221_X1 U33351 ( .B1(n39223), .B2(n29410), .C1(n39217), .C2(n29474), .A(
        n36923), .ZN(n36918) );
  OAI222_X1 U33352 ( .A1(n31670), .A2(n39211), .B1(n31734), .B2(n39205), .C1(
        n31606), .C2(n39199), .ZN(n36923) );
  AOI221_X1 U33353 ( .B1(n39223), .B2(n29409), .C1(n39217), .C2(n29473), .A(
        n36904), .ZN(n36899) );
  OAI222_X1 U33354 ( .A1(n31669), .A2(n39211), .B1(n31733), .B2(n39205), .C1(
        n31605), .C2(n39199), .ZN(n36904) );
  AOI221_X1 U33355 ( .B1(n39223), .B2(n29408), .C1(n39217), .C2(n29472), .A(
        n36885), .ZN(n36880) );
  OAI222_X1 U33356 ( .A1(n31668), .A2(n39211), .B1(n31732), .B2(n39205), .C1(
        n31604), .C2(n39199), .ZN(n36885) );
  AOI221_X1 U33357 ( .B1(n39223), .B2(n29407), .C1(n39217), .C2(n29471), .A(
        n36866), .ZN(n36861) );
  OAI222_X1 U33358 ( .A1(n31667), .A2(n39211), .B1(n31731), .B2(n39205), .C1(
        n31603), .C2(n39199), .ZN(n36866) );
  AOI221_X1 U33359 ( .B1(n39223), .B2(n29406), .C1(n39217), .C2(n29470), .A(
        n36847), .ZN(n36842) );
  OAI222_X1 U33360 ( .A1(n31666), .A2(n39211), .B1(n31730), .B2(n39205), .C1(
        n31602), .C2(n39199), .ZN(n36847) );
  AOI221_X1 U33361 ( .B1(n39223), .B2(n29405), .C1(n39217), .C2(n29469), .A(
        n36828), .ZN(n36823) );
  OAI222_X1 U33362 ( .A1(n31665), .A2(n39211), .B1(n31729), .B2(n39205), .C1(
        n31601), .C2(n39199), .ZN(n36828) );
  AOI221_X1 U33363 ( .B1(n39223), .B2(n29404), .C1(n39217), .C2(n29468), .A(
        n36809), .ZN(n36804) );
  OAI222_X1 U33364 ( .A1(n31664), .A2(n39211), .B1(n31728), .B2(n39205), .C1(
        n31600), .C2(n39199), .ZN(n36809) );
  AOI221_X1 U33365 ( .B1(n39223), .B2(n29403), .C1(n39217), .C2(n29467), .A(
        n36790), .ZN(n36785) );
  OAI222_X1 U33366 ( .A1(n31663), .A2(n39211), .B1(n31727), .B2(n39205), .C1(
        n31599), .C2(n39199), .ZN(n36790) );
  AOI221_X1 U33367 ( .B1(n39224), .B2(n29402), .C1(n39218), .C2(n29466), .A(
        n36771), .ZN(n36766) );
  OAI222_X1 U33368 ( .A1(n31662), .A2(n39212), .B1(n31726), .B2(n39206), .C1(
        n31598), .C2(n39200), .ZN(n36771) );
  AOI221_X1 U33369 ( .B1(n39224), .B2(n29401), .C1(n39218), .C2(n29465), .A(
        n36752), .ZN(n36747) );
  OAI222_X1 U33370 ( .A1(n31661), .A2(n39212), .B1(n31725), .B2(n39206), .C1(
        n31597), .C2(n39200), .ZN(n36752) );
  AOI221_X1 U33371 ( .B1(n39224), .B2(n29400), .C1(n39218), .C2(n29464), .A(
        n36733), .ZN(n36728) );
  OAI222_X1 U33372 ( .A1(n31660), .A2(n39212), .B1(n31724), .B2(n39206), .C1(
        n31596), .C2(n39200), .ZN(n36733) );
  AOI221_X1 U33373 ( .B1(n39224), .B2(n29399), .C1(n39218), .C2(n29463), .A(
        n36714), .ZN(n36709) );
  OAI222_X1 U33374 ( .A1(n31659), .A2(n39212), .B1(n31723), .B2(n39206), .C1(
        n31595), .C2(n39200), .ZN(n36714) );
  AOI221_X1 U33375 ( .B1(n39224), .B2(n29398), .C1(n39218), .C2(n29462), .A(
        n36695), .ZN(n36690) );
  OAI222_X1 U33376 ( .A1(n31658), .A2(n39212), .B1(n31722), .B2(n39206), .C1(
        n31594), .C2(n39200), .ZN(n36695) );
  AOI221_X1 U33377 ( .B1(n39224), .B2(n29397), .C1(n39218), .C2(n29461), .A(
        n36676), .ZN(n36671) );
  OAI222_X1 U33378 ( .A1(n31657), .A2(n39212), .B1(n31721), .B2(n39206), .C1(
        n31593), .C2(n39200), .ZN(n36676) );
  AOI221_X1 U33379 ( .B1(n39224), .B2(n29396), .C1(n39218), .C2(n29460), .A(
        n36657), .ZN(n36652) );
  OAI222_X1 U33380 ( .A1(n31656), .A2(n39212), .B1(n31720), .B2(n39206), .C1(
        n31592), .C2(n39200), .ZN(n36657) );
  AOI221_X1 U33381 ( .B1(n39224), .B2(n29395), .C1(n39218), .C2(n29459), .A(
        n36638), .ZN(n36633) );
  OAI222_X1 U33382 ( .A1(n31655), .A2(n39212), .B1(n31719), .B2(n39206), .C1(
        n31591), .C2(n39200), .ZN(n36638) );
  AOI221_X1 U33383 ( .B1(n39224), .B2(n29394), .C1(n39218), .C2(n29458), .A(
        n36619), .ZN(n36614) );
  OAI222_X1 U33384 ( .A1(n31654), .A2(n39212), .B1(n31718), .B2(n39206), .C1(
        n31590), .C2(n39200), .ZN(n36619) );
  AOI221_X1 U33385 ( .B1(n39224), .B2(n29393), .C1(n39218), .C2(n29457), .A(
        n36600), .ZN(n36595) );
  OAI222_X1 U33386 ( .A1(n31653), .A2(n39212), .B1(n31717), .B2(n39206), .C1(
        n31589), .C2(n39200), .ZN(n36600) );
  AOI221_X1 U33387 ( .B1(n39224), .B2(n29392), .C1(n39218), .C2(n29456), .A(
        n36581), .ZN(n36576) );
  OAI222_X1 U33388 ( .A1(n31652), .A2(n39212), .B1(n31716), .B2(n39206), .C1(
        n31588), .C2(n39200), .ZN(n36581) );
  AOI221_X1 U33389 ( .B1(n39224), .B2(n29391), .C1(n39218), .C2(n29455), .A(
        n36562), .ZN(n36557) );
  OAI222_X1 U33390 ( .A1(n31651), .A2(n39212), .B1(n31715), .B2(n39206), .C1(
        n31587), .C2(n39200), .ZN(n36562) );
  AOI221_X1 U33391 ( .B1(n39225), .B2(n29390), .C1(n39219), .C2(n29454), .A(
        n36543), .ZN(n36538) );
  OAI222_X1 U33392 ( .A1(n31650), .A2(n39213), .B1(n31714), .B2(n39207), .C1(
        n31586), .C2(n39201), .ZN(n36543) );
  AOI221_X1 U33393 ( .B1(n39225), .B2(n29389), .C1(n39219), .C2(n29453), .A(
        n36524), .ZN(n36519) );
  OAI222_X1 U33394 ( .A1(n31649), .A2(n39213), .B1(n31713), .B2(n39207), .C1(
        n31585), .C2(n39201), .ZN(n36524) );
  AOI221_X1 U33395 ( .B1(n39225), .B2(n29388), .C1(n39219), .C2(n29452), .A(
        n36505), .ZN(n36500) );
  OAI222_X1 U33396 ( .A1(n31648), .A2(n39213), .B1(n31712), .B2(n39207), .C1(
        n31584), .C2(n39201), .ZN(n36505) );
  AOI221_X1 U33397 ( .B1(n39225), .B2(n29387), .C1(n39219), .C2(n29451), .A(
        n36486), .ZN(n36481) );
  OAI222_X1 U33398 ( .A1(n31647), .A2(n39213), .B1(n31711), .B2(n39207), .C1(
        n31583), .C2(n39201), .ZN(n36486) );
  AOI221_X1 U33399 ( .B1(n39225), .B2(n29386), .C1(n39219), .C2(n29450), .A(
        n36467), .ZN(n36462) );
  OAI222_X1 U33400 ( .A1(n31646), .A2(n39213), .B1(n31710), .B2(n39207), .C1(
        n31582), .C2(n39201), .ZN(n36467) );
  AOI221_X1 U33401 ( .B1(n39225), .B2(n29385), .C1(n39219), .C2(n29449), .A(
        n36448), .ZN(n36443) );
  OAI222_X1 U33402 ( .A1(n31645), .A2(n39213), .B1(n31709), .B2(n39207), .C1(
        n31581), .C2(n39201), .ZN(n36448) );
  AOI221_X1 U33403 ( .B1(n39225), .B2(n29384), .C1(n39219), .C2(n29448), .A(
        n36429), .ZN(n36424) );
  OAI222_X1 U33404 ( .A1(n31644), .A2(n39213), .B1(n31708), .B2(n39207), .C1(
        n31580), .C2(n39201), .ZN(n36429) );
  AOI221_X1 U33405 ( .B1(n39225), .B2(n29383), .C1(n39219), .C2(n29447), .A(
        n36410), .ZN(n36405) );
  OAI222_X1 U33406 ( .A1(n31643), .A2(n39213), .B1(n31707), .B2(n39207), .C1(
        n31579), .C2(n39201), .ZN(n36410) );
  AOI221_X1 U33407 ( .B1(n39225), .B2(n29382), .C1(n39219), .C2(n29446), .A(
        n36391), .ZN(n36386) );
  OAI222_X1 U33408 ( .A1(n31642), .A2(n39213), .B1(n31706), .B2(n39207), .C1(
        n31578), .C2(n39201), .ZN(n36391) );
  AOI221_X1 U33409 ( .B1(n39225), .B2(n29381), .C1(n39219), .C2(n29445), .A(
        n36372), .ZN(n36367) );
  OAI222_X1 U33410 ( .A1(n31641), .A2(n39213), .B1(n31705), .B2(n39207), .C1(
        n31577), .C2(n39201), .ZN(n36372) );
  AOI221_X1 U33411 ( .B1(n39225), .B2(n29380), .C1(n39219), .C2(n29444), .A(
        n36353), .ZN(n36348) );
  OAI222_X1 U33412 ( .A1(n31640), .A2(n39213), .B1(n31704), .B2(n39207), .C1(
        n31576), .C2(n39201), .ZN(n36353) );
  AOI221_X1 U33413 ( .B1(n39225), .B2(n29379), .C1(n39219), .C2(n29443), .A(
        n36334), .ZN(n36329) );
  OAI222_X1 U33414 ( .A1(n31639), .A2(n39213), .B1(n31703), .B2(n39207), .C1(
        n31575), .C2(n39201), .ZN(n36334) );
  AOI221_X1 U33415 ( .B1(n39226), .B2(n29378), .C1(n39220), .C2(n29442), .A(
        n36315), .ZN(n36310) );
  OAI222_X1 U33416 ( .A1(n31638), .A2(n39214), .B1(n31702), .B2(n39208), .C1(
        n31574), .C2(n39202), .ZN(n36315) );
  AOI221_X1 U33417 ( .B1(n39226), .B2(n29377), .C1(n39220), .C2(n29441), .A(
        n36296), .ZN(n36291) );
  OAI222_X1 U33418 ( .A1(n31637), .A2(n39214), .B1(n31701), .B2(n39208), .C1(
        n31573), .C2(n39202), .ZN(n36296) );
  AOI221_X1 U33419 ( .B1(n39226), .B2(n29376), .C1(n39220), .C2(n29440), .A(
        n36277), .ZN(n36272) );
  OAI222_X1 U33420 ( .A1(n31636), .A2(n39214), .B1(n31700), .B2(n39208), .C1(
        n31572), .C2(n39202), .ZN(n36277) );
  AOI221_X1 U33421 ( .B1(n39226), .B2(n29375), .C1(n39220), .C2(n29439), .A(
        n36258), .ZN(n36253) );
  OAI222_X1 U33422 ( .A1(n31635), .A2(n39214), .B1(n31699), .B2(n39208), .C1(
        n31571), .C2(n39202), .ZN(n36258) );
  AOI221_X1 U33423 ( .B1(n39226), .B2(n29374), .C1(n39220), .C2(n29438), .A(
        n36239), .ZN(n36234) );
  OAI222_X1 U33424 ( .A1(n31634), .A2(n39214), .B1(n31698), .B2(n39208), .C1(
        n31570), .C2(n39202), .ZN(n36239) );
  AOI221_X1 U33425 ( .B1(n39226), .B2(n29373), .C1(n39220), .C2(n29437), .A(
        n36220), .ZN(n36215) );
  OAI222_X1 U33426 ( .A1(n31633), .A2(n39214), .B1(n31697), .B2(n39208), .C1(
        n31569), .C2(n39202), .ZN(n36220) );
  AOI221_X1 U33427 ( .B1(n39222), .B2(n29425), .C1(n39216), .C2(n29489), .A(
        n37208), .ZN(n37203) );
  OAI222_X1 U33428 ( .A1(n31685), .A2(n39210), .B1(n31749), .B2(n39204), .C1(
        n31621), .C2(n39198), .ZN(n37208) );
  AOI221_X1 U33429 ( .B1(n39222), .B2(n29424), .C1(n39216), .C2(n29488), .A(
        n37189), .ZN(n37184) );
  OAI222_X1 U33430 ( .A1(n31684), .A2(n39210), .B1(n31748), .B2(n39204), .C1(
        n31620), .C2(n39198), .ZN(n37189) );
  AOI221_X1 U33431 ( .B1(n39222), .B2(n29423), .C1(n39216), .C2(n29487), .A(
        n37170), .ZN(n37165) );
  OAI222_X1 U33432 ( .A1(n31683), .A2(n39210), .B1(n31747), .B2(n39204), .C1(
        n31619), .C2(n39198), .ZN(n37170) );
  AOI221_X1 U33433 ( .B1(n39222), .B2(n29422), .C1(n39216), .C2(n29486), .A(
        n37151), .ZN(n37146) );
  OAI222_X1 U33434 ( .A1(n31682), .A2(n39210), .B1(n31746), .B2(n39204), .C1(
        n31618), .C2(n39198), .ZN(n37151) );
  AOI221_X1 U33435 ( .B1(n39222), .B2(n29421), .C1(n39216), .C2(n29485), .A(
        n37132), .ZN(n37127) );
  OAI222_X1 U33436 ( .A1(n31681), .A2(n39210), .B1(n31745), .B2(n39204), .C1(
        n31617), .C2(n39198), .ZN(n37132) );
  AOI221_X1 U33437 ( .B1(n39227), .B2(n29366), .C1(n39221), .C2(n29430), .A(
        n36087), .ZN(n36082) );
  OAI222_X1 U33438 ( .A1(n31626), .A2(n39215), .B1(n31690), .B2(n39209), .C1(
        n31562), .C2(n39203), .ZN(n36087) );
  AOI221_X1 U33439 ( .B1(n39227), .B2(n29365), .C1(n39221), .C2(n29429), .A(
        n36068), .ZN(n36063) );
  OAI222_X1 U33440 ( .A1(n31625), .A2(n39215), .B1(n31689), .B2(n39209), .C1(
        n31561), .C2(n39203), .ZN(n36068) );
  AOI221_X1 U33441 ( .B1(n39227), .B2(n29364), .C1(n39221), .C2(n29428), .A(
        n36049), .ZN(n36044) );
  OAI222_X1 U33442 ( .A1(n31624), .A2(n39215), .B1(n31688), .B2(n39209), .C1(
        n31560), .C2(n39203), .ZN(n36049) );
  AOI221_X1 U33443 ( .B1(n39227), .B2(n29363), .C1(n39221), .C2(n29427), .A(
        n36002), .ZN(n35985) );
  OAI222_X1 U33444 ( .A1(n31623), .A2(n39215), .B1(n31687), .B2(n39209), .C1(
        n31559), .C2(n39203), .ZN(n36002) );
  AOI221_X1 U33445 ( .B1(n39222), .B2(n29426), .C1(n39216), .C2(n29490), .A(
        n37237), .ZN(n37222) );
  OAI222_X1 U33446 ( .A1(n31686), .A2(n39210), .B1(n31750), .B2(n39204), .C1(
        n31622), .C2(n39198), .ZN(n37237) );
  AOI221_X1 U33447 ( .B1(n39222), .B2(n29420), .C1(n39216), .C2(n29484), .A(
        n37113), .ZN(n37108) );
  OAI222_X1 U33448 ( .A1(n31680), .A2(n39210), .B1(n31744), .B2(n39204), .C1(
        n31616), .C2(n39198), .ZN(n37113) );
  AOI221_X1 U33449 ( .B1(n39222), .B2(n29419), .C1(n39216), .C2(n29483), .A(
        n37094), .ZN(n37089) );
  OAI222_X1 U33450 ( .A1(n31679), .A2(n39210), .B1(n31743), .B2(n39204), .C1(
        n31615), .C2(n39198), .ZN(n37094) );
  AOI221_X1 U33451 ( .B1(n39222), .B2(n29418), .C1(n39216), .C2(n29482), .A(
        n37075), .ZN(n37070) );
  OAI222_X1 U33452 ( .A1(n31678), .A2(n39210), .B1(n31742), .B2(n39204), .C1(
        n31614), .C2(n39198), .ZN(n37075) );
  AOI221_X1 U33453 ( .B1(n39222), .B2(n29417), .C1(n39216), .C2(n29481), .A(
        n37056), .ZN(n37051) );
  OAI222_X1 U33454 ( .A1(n31677), .A2(n39210), .B1(n31741), .B2(n39204), .C1(
        n31613), .C2(n39198), .ZN(n37056) );
  AOI221_X1 U33455 ( .B1(n39222), .B2(n29416), .C1(n39216), .C2(n29480), .A(
        n37037), .ZN(n37032) );
  OAI222_X1 U33456 ( .A1(n31676), .A2(n39210), .B1(n31740), .B2(n39204), .C1(
        n31612), .C2(n39198), .ZN(n37037) );
  AOI221_X1 U33457 ( .B1(n39226), .B2(n29372), .C1(n39220), .C2(n29436), .A(
        n36201), .ZN(n36196) );
  OAI222_X1 U33458 ( .A1(n31632), .A2(n39214), .B1(n31696), .B2(n39208), .C1(
        n31568), .C2(n39202), .ZN(n36201) );
  AOI221_X1 U33459 ( .B1(n39226), .B2(n29371), .C1(n39220), .C2(n29435), .A(
        n36182), .ZN(n36177) );
  OAI222_X1 U33460 ( .A1(n31631), .A2(n39214), .B1(n31695), .B2(n39208), .C1(
        n31567), .C2(n39202), .ZN(n36182) );
  AOI221_X1 U33461 ( .B1(n39226), .B2(n29370), .C1(n39220), .C2(n29434), .A(
        n36163), .ZN(n36158) );
  OAI222_X1 U33462 ( .A1(n31630), .A2(n39214), .B1(n31694), .B2(n39208), .C1(
        n31566), .C2(n39202), .ZN(n36163) );
  AOI221_X1 U33463 ( .B1(n39226), .B2(n29369), .C1(n39220), .C2(n29433), .A(
        n36144), .ZN(n36139) );
  OAI222_X1 U33464 ( .A1(n31629), .A2(n39214), .B1(n31693), .B2(n39208), .C1(
        n31565), .C2(n39202), .ZN(n36144) );
  AOI221_X1 U33465 ( .B1(n39226), .B2(n29368), .C1(n39220), .C2(n29432), .A(
        n36125), .ZN(n36120) );
  OAI222_X1 U33466 ( .A1(n31628), .A2(n39214), .B1(n31692), .B2(n39208), .C1(
        n31564), .C2(n39202), .ZN(n36125) );
  AOI221_X1 U33467 ( .B1(n39226), .B2(n29367), .C1(n39220), .C2(n29431), .A(
        n36106), .ZN(n36101) );
  OAI222_X1 U33468 ( .A1(n31627), .A2(n39214), .B1(n31691), .B2(n39208), .C1(
        n31563), .C2(n39202), .ZN(n36106) );
  AOI221_X1 U33469 ( .B1(n39729), .B2(n29426), .C1(n39723), .C2(n29490), .A(
        n33447), .ZN(n33430) );
  OAI222_X1 U33470 ( .A1(n31686), .A2(n39717), .B1(n31750), .B2(n39711), .C1(
        n31622), .C2(n39705), .ZN(n33447) );
  AOI221_X1 U33471 ( .B1(n39477), .B2(n29426), .C1(n39471), .C2(n29490), .A(
        n34721), .ZN(n34704) );
  OAI222_X1 U33472 ( .A1(n31686), .A2(n39465), .B1(n31750), .B2(n39459), .C1(
        n31622), .C2(n39453), .ZN(n34721) );
  AOI221_X1 U33473 ( .B1(n39729), .B2(n29425), .C1(n39723), .C2(n29489), .A(
        n33494), .ZN(n33489) );
  OAI222_X1 U33474 ( .A1(n31685), .A2(n39717), .B1(n31749), .B2(n39711), .C1(
        n31621), .C2(n39705), .ZN(n33494) );
  AOI221_X1 U33475 ( .B1(n39477), .B2(n29425), .C1(n39471), .C2(n29489), .A(
        n34768), .ZN(n34763) );
  OAI222_X1 U33476 ( .A1(n31685), .A2(n39465), .B1(n31749), .B2(n39459), .C1(
        n31621), .C2(n39453), .ZN(n34768) );
  AOI221_X1 U33477 ( .B1(n39729), .B2(n29424), .C1(n39723), .C2(n29488), .A(
        n33513), .ZN(n33508) );
  OAI222_X1 U33478 ( .A1(n31684), .A2(n39717), .B1(n31748), .B2(n39711), .C1(
        n31620), .C2(n39705), .ZN(n33513) );
  AOI221_X1 U33479 ( .B1(n39477), .B2(n29424), .C1(n39471), .C2(n29488), .A(
        n34787), .ZN(n34782) );
  OAI222_X1 U33480 ( .A1(n31684), .A2(n39465), .B1(n31748), .B2(n39459), .C1(
        n31620), .C2(n39453), .ZN(n34787) );
  AOI221_X1 U33481 ( .B1(n39729), .B2(n29423), .C1(n39723), .C2(n29487), .A(
        n33532), .ZN(n33527) );
  OAI222_X1 U33482 ( .A1(n31683), .A2(n39717), .B1(n31747), .B2(n39711), .C1(
        n31619), .C2(n39705), .ZN(n33532) );
  AOI221_X1 U33483 ( .B1(n39477), .B2(n29423), .C1(n39471), .C2(n29487), .A(
        n34806), .ZN(n34801) );
  OAI222_X1 U33484 ( .A1(n31683), .A2(n39465), .B1(n31747), .B2(n39459), .C1(
        n31619), .C2(n39453), .ZN(n34806) );
  AOI221_X1 U33485 ( .B1(n39728), .B2(n29422), .C1(n39722), .C2(n29486), .A(
        n33551), .ZN(n33546) );
  OAI222_X1 U33486 ( .A1(n31682), .A2(n39716), .B1(n31746), .B2(n39710), .C1(
        n31618), .C2(n39704), .ZN(n33551) );
  AOI221_X1 U33487 ( .B1(n39476), .B2(n29422), .C1(n39470), .C2(n29486), .A(
        n34825), .ZN(n34820) );
  OAI222_X1 U33488 ( .A1(n31682), .A2(n39464), .B1(n31746), .B2(n39458), .C1(
        n31618), .C2(n39452), .ZN(n34825) );
  AOI221_X1 U33489 ( .B1(n39728), .B2(n29421), .C1(n39722), .C2(n29485), .A(
        n33570), .ZN(n33565) );
  OAI222_X1 U33490 ( .A1(n31681), .A2(n39716), .B1(n31745), .B2(n39710), .C1(
        n31617), .C2(n39704), .ZN(n33570) );
  AOI221_X1 U33491 ( .B1(n39476), .B2(n29421), .C1(n39470), .C2(n29485), .A(
        n34844), .ZN(n34839) );
  OAI222_X1 U33492 ( .A1(n31681), .A2(n39464), .B1(n31745), .B2(n39458), .C1(
        n31617), .C2(n39452), .ZN(n34844) );
  AOI221_X1 U33493 ( .B1(n39728), .B2(n29420), .C1(n39722), .C2(n29484), .A(
        n33589), .ZN(n33584) );
  OAI222_X1 U33494 ( .A1(n31680), .A2(n39716), .B1(n31744), .B2(n39710), .C1(
        n31616), .C2(n39704), .ZN(n33589) );
  AOI221_X1 U33495 ( .B1(n39476), .B2(n29420), .C1(n39470), .C2(n29484), .A(
        n34863), .ZN(n34858) );
  OAI222_X1 U33496 ( .A1(n31680), .A2(n39464), .B1(n31744), .B2(n39458), .C1(
        n31616), .C2(n39452), .ZN(n34863) );
  AOI221_X1 U33497 ( .B1(n39728), .B2(n29419), .C1(n39722), .C2(n29483), .A(
        n33608), .ZN(n33603) );
  OAI222_X1 U33498 ( .A1(n31679), .A2(n39716), .B1(n31743), .B2(n39710), .C1(
        n31615), .C2(n39704), .ZN(n33608) );
  AOI221_X1 U33499 ( .B1(n39476), .B2(n29419), .C1(n39470), .C2(n29483), .A(
        n34882), .ZN(n34877) );
  OAI222_X1 U33500 ( .A1(n31679), .A2(n39464), .B1(n31743), .B2(n39458), .C1(
        n31615), .C2(n39452), .ZN(n34882) );
  AOI221_X1 U33501 ( .B1(n39728), .B2(n29418), .C1(n39722), .C2(n29482), .A(
        n33627), .ZN(n33622) );
  OAI222_X1 U33502 ( .A1(n31678), .A2(n39716), .B1(n31742), .B2(n39710), .C1(
        n31614), .C2(n39704), .ZN(n33627) );
  AOI221_X1 U33503 ( .B1(n39476), .B2(n29418), .C1(n39470), .C2(n29482), .A(
        n34901), .ZN(n34896) );
  OAI222_X1 U33504 ( .A1(n31678), .A2(n39464), .B1(n31742), .B2(n39458), .C1(
        n31614), .C2(n39452), .ZN(n34901) );
  AOI221_X1 U33505 ( .B1(n39728), .B2(n29417), .C1(n39722), .C2(n29481), .A(
        n33646), .ZN(n33641) );
  OAI222_X1 U33506 ( .A1(n31677), .A2(n39716), .B1(n31741), .B2(n39710), .C1(
        n31613), .C2(n39704), .ZN(n33646) );
  AOI221_X1 U33507 ( .B1(n39476), .B2(n29417), .C1(n39470), .C2(n29481), .A(
        n34920), .ZN(n34915) );
  OAI222_X1 U33508 ( .A1(n31677), .A2(n39464), .B1(n31741), .B2(n39458), .C1(
        n31613), .C2(n39452), .ZN(n34920) );
  AOI221_X1 U33509 ( .B1(n39728), .B2(n29416), .C1(n39722), .C2(n29480), .A(
        n33665), .ZN(n33660) );
  OAI222_X1 U33510 ( .A1(n31676), .A2(n39716), .B1(n31740), .B2(n39710), .C1(
        n31612), .C2(n39704), .ZN(n33665) );
  AOI221_X1 U33511 ( .B1(n39476), .B2(n29416), .C1(n39470), .C2(n29480), .A(
        n34939), .ZN(n34934) );
  OAI222_X1 U33512 ( .A1(n31676), .A2(n39464), .B1(n31740), .B2(n39458), .C1(
        n31612), .C2(n39452), .ZN(n34939) );
  AOI221_X1 U33513 ( .B1(n39728), .B2(n29415), .C1(n39722), .C2(n29479), .A(
        n33684), .ZN(n33679) );
  OAI222_X1 U33514 ( .A1(n31675), .A2(n39716), .B1(n31739), .B2(n39710), .C1(
        n31611), .C2(n39704), .ZN(n33684) );
  AOI221_X1 U33515 ( .B1(n39476), .B2(n29415), .C1(n39470), .C2(n29479), .A(
        n34958), .ZN(n34953) );
  OAI222_X1 U33516 ( .A1(n31675), .A2(n39464), .B1(n31739), .B2(n39458), .C1(
        n31611), .C2(n39452), .ZN(n34958) );
  AOI221_X1 U33517 ( .B1(n39728), .B2(n29414), .C1(n39722), .C2(n29478), .A(
        n33703), .ZN(n33698) );
  OAI222_X1 U33518 ( .A1(n31674), .A2(n39716), .B1(n31738), .B2(n39710), .C1(
        n31610), .C2(n39704), .ZN(n33703) );
  AOI221_X1 U33519 ( .B1(n39476), .B2(n29414), .C1(n39470), .C2(n29478), .A(
        n34977), .ZN(n34972) );
  OAI222_X1 U33520 ( .A1(n31674), .A2(n39464), .B1(n31738), .B2(n39458), .C1(
        n31610), .C2(n39452), .ZN(n34977) );
  AOI221_X1 U33521 ( .B1(n39728), .B2(n29413), .C1(n39722), .C2(n29477), .A(
        n33722), .ZN(n33717) );
  OAI222_X1 U33522 ( .A1(n31673), .A2(n39716), .B1(n31737), .B2(n39710), .C1(
        n31609), .C2(n39704), .ZN(n33722) );
  AOI221_X1 U33523 ( .B1(n39476), .B2(n29413), .C1(n39470), .C2(n29477), .A(
        n34996), .ZN(n34991) );
  OAI222_X1 U33524 ( .A1(n31673), .A2(n39464), .B1(n31737), .B2(n39458), .C1(
        n31609), .C2(n39452), .ZN(n34996) );
  AOI221_X1 U33525 ( .B1(n39728), .B2(n29412), .C1(n39722), .C2(n29476), .A(
        n33741), .ZN(n33736) );
  OAI222_X1 U33526 ( .A1(n31672), .A2(n39716), .B1(n31736), .B2(n39710), .C1(
        n31608), .C2(n39704), .ZN(n33741) );
  AOI221_X1 U33527 ( .B1(n39476), .B2(n29412), .C1(n39470), .C2(n29476), .A(
        n35015), .ZN(n35010) );
  OAI222_X1 U33528 ( .A1(n31672), .A2(n39464), .B1(n31736), .B2(n39458), .C1(
        n31608), .C2(n39452), .ZN(n35015) );
  AOI221_X1 U33529 ( .B1(n39728), .B2(n29411), .C1(n39722), .C2(n29475), .A(
        n33760), .ZN(n33755) );
  OAI222_X1 U33530 ( .A1(n31671), .A2(n39716), .B1(n31735), .B2(n39710), .C1(
        n31607), .C2(n39704), .ZN(n33760) );
  AOI221_X1 U33531 ( .B1(n39476), .B2(n29411), .C1(n39470), .C2(n29475), .A(
        n35034), .ZN(n35029) );
  OAI222_X1 U33532 ( .A1(n31671), .A2(n39464), .B1(n31735), .B2(n39458), .C1(
        n31607), .C2(n39452), .ZN(n35034) );
  AOI221_X1 U33533 ( .B1(n39727), .B2(n29410), .C1(n39721), .C2(n29474), .A(
        n33779), .ZN(n33774) );
  OAI222_X1 U33534 ( .A1(n31670), .A2(n39715), .B1(n31734), .B2(n39709), .C1(
        n31606), .C2(n39703), .ZN(n33779) );
  AOI221_X1 U33535 ( .B1(n39475), .B2(n29410), .C1(n39469), .C2(n29474), .A(
        n35053), .ZN(n35048) );
  OAI222_X1 U33536 ( .A1(n31670), .A2(n39463), .B1(n31734), .B2(n39457), .C1(
        n31606), .C2(n39451), .ZN(n35053) );
  AOI221_X1 U33537 ( .B1(n39727), .B2(n29409), .C1(n39721), .C2(n29473), .A(
        n33798), .ZN(n33793) );
  OAI222_X1 U33538 ( .A1(n31669), .A2(n39715), .B1(n31733), .B2(n39709), .C1(
        n31605), .C2(n39703), .ZN(n33798) );
  AOI221_X1 U33539 ( .B1(n39475), .B2(n29409), .C1(n39469), .C2(n29473), .A(
        n35072), .ZN(n35067) );
  OAI222_X1 U33540 ( .A1(n31669), .A2(n39463), .B1(n31733), .B2(n39457), .C1(
        n31605), .C2(n39451), .ZN(n35072) );
  AOI221_X1 U33541 ( .B1(n39727), .B2(n29408), .C1(n39721), .C2(n29472), .A(
        n33817), .ZN(n33812) );
  OAI222_X1 U33542 ( .A1(n31668), .A2(n39715), .B1(n31732), .B2(n39709), .C1(
        n31604), .C2(n39703), .ZN(n33817) );
  AOI221_X1 U33543 ( .B1(n39475), .B2(n29408), .C1(n39469), .C2(n29472), .A(
        n35091), .ZN(n35086) );
  OAI222_X1 U33544 ( .A1(n31668), .A2(n39463), .B1(n31732), .B2(n39457), .C1(
        n31604), .C2(n39451), .ZN(n35091) );
  AOI221_X1 U33545 ( .B1(n39727), .B2(n29407), .C1(n39721), .C2(n29471), .A(
        n33836), .ZN(n33831) );
  OAI222_X1 U33546 ( .A1(n31667), .A2(n39715), .B1(n31731), .B2(n39709), .C1(
        n31603), .C2(n39703), .ZN(n33836) );
  AOI221_X1 U33547 ( .B1(n39475), .B2(n29407), .C1(n39469), .C2(n29471), .A(
        n35110), .ZN(n35105) );
  OAI222_X1 U33548 ( .A1(n31667), .A2(n39463), .B1(n31731), .B2(n39457), .C1(
        n31603), .C2(n39451), .ZN(n35110) );
  AOI221_X1 U33549 ( .B1(n39727), .B2(n29406), .C1(n39721), .C2(n29470), .A(
        n33855), .ZN(n33850) );
  OAI222_X1 U33550 ( .A1(n31666), .A2(n39715), .B1(n31730), .B2(n39709), .C1(
        n31602), .C2(n39703), .ZN(n33855) );
  AOI221_X1 U33551 ( .B1(n39475), .B2(n29406), .C1(n39469), .C2(n29470), .A(
        n35129), .ZN(n35124) );
  OAI222_X1 U33552 ( .A1(n31666), .A2(n39463), .B1(n31730), .B2(n39457), .C1(
        n31602), .C2(n39451), .ZN(n35129) );
  AOI221_X1 U33553 ( .B1(n39727), .B2(n29405), .C1(n39721), .C2(n29469), .A(
        n33874), .ZN(n33869) );
  OAI222_X1 U33554 ( .A1(n31665), .A2(n39715), .B1(n31729), .B2(n39709), .C1(
        n31601), .C2(n39703), .ZN(n33874) );
  AOI221_X1 U33555 ( .B1(n39475), .B2(n29405), .C1(n39469), .C2(n29469), .A(
        n35148), .ZN(n35143) );
  OAI222_X1 U33556 ( .A1(n31665), .A2(n39463), .B1(n31729), .B2(n39457), .C1(
        n31601), .C2(n39451), .ZN(n35148) );
  AOI221_X1 U33557 ( .B1(n39727), .B2(n29404), .C1(n39721), .C2(n29468), .A(
        n33893), .ZN(n33888) );
  OAI222_X1 U33558 ( .A1(n31664), .A2(n39715), .B1(n31728), .B2(n39709), .C1(
        n31600), .C2(n39703), .ZN(n33893) );
  AOI221_X1 U33559 ( .B1(n39475), .B2(n29404), .C1(n39469), .C2(n29468), .A(
        n35167), .ZN(n35162) );
  OAI222_X1 U33560 ( .A1(n31664), .A2(n39463), .B1(n31728), .B2(n39457), .C1(
        n31600), .C2(n39451), .ZN(n35167) );
  AOI221_X1 U33561 ( .B1(n39727), .B2(n29403), .C1(n39721), .C2(n29467), .A(
        n33912), .ZN(n33907) );
  OAI222_X1 U33562 ( .A1(n31663), .A2(n39715), .B1(n31727), .B2(n39709), .C1(
        n31599), .C2(n39703), .ZN(n33912) );
  AOI221_X1 U33563 ( .B1(n39475), .B2(n29403), .C1(n39469), .C2(n29467), .A(
        n35186), .ZN(n35181) );
  OAI222_X1 U33564 ( .A1(n31663), .A2(n39463), .B1(n31727), .B2(n39457), .C1(
        n31599), .C2(n39451), .ZN(n35186) );
  AOI221_X1 U33565 ( .B1(n39727), .B2(n29402), .C1(n39721), .C2(n29466), .A(
        n33931), .ZN(n33926) );
  OAI222_X1 U33566 ( .A1(n31662), .A2(n39715), .B1(n31726), .B2(n39709), .C1(
        n31598), .C2(n39703), .ZN(n33931) );
  AOI221_X1 U33567 ( .B1(n39475), .B2(n29402), .C1(n39469), .C2(n29466), .A(
        n35205), .ZN(n35200) );
  OAI222_X1 U33568 ( .A1(n31662), .A2(n39463), .B1(n31726), .B2(n39457), .C1(
        n31598), .C2(n39451), .ZN(n35205) );
  AOI221_X1 U33569 ( .B1(n39727), .B2(n29401), .C1(n39721), .C2(n29465), .A(
        n33950), .ZN(n33945) );
  OAI222_X1 U33570 ( .A1(n31661), .A2(n39715), .B1(n31725), .B2(n39709), .C1(
        n31597), .C2(n39703), .ZN(n33950) );
  AOI221_X1 U33571 ( .B1(n39475), .B2(n29401), .C1(n39469), .C2(n29465), .A(
        n35224), .ZN(n35219) );
  OAI222_X1 U33572 ( .A1(n31661), .A2(n39463), .B1(n31725), .B2(n39457), .C1(
        n31597), .C2(n39451), .ZN(n35224) );
  AOI221_X1 U33573 ( .B1(n39727), .B2(n29400), .C1(n39721), .C2(n29464), .A(
        n33969), .ZN(n33964) );
  OAI222_X1 U33574 ( .A1(n31660), .A2(n39715), .B1(n31724), .B2(n39709), .C1(
        n31596), .C2(n39703), .ZN(n33969) );
  AOI221_X1 U33575 ( .B1(n39475), .B2(n29400), .C1(n39469), .C2(n29464), .A(
        n35243), .ZN(n35238) );
  OAI222_X1 U33576 ( .A1(n31660), .A2(n39463), .B1(n31724), .B2(n39457), .C1(
        n31596), .C2(n39451), .ZN(n35243) );
  AOI221_X1 U33577 ( .B1(n39727), .B2(n29399), .C1(n39721), .C2(n29463), .A(
        n33988), .ZN(n33983) );
  OAI222_X1 U33578 ( .A1(n31659), .A2(n39715), .B1(n31723), .B2(n39709), .C1(
        n31595), .C2(n39703), .ZN(n33988) );
  AOI221_X1 U33579 ( .B1(n39475), .B2(n29399), .C1(n39469), .C2(n29463), .A(
        n35262), .ZN(n35257) );
  OAI222_X1 U33580 ( .A1(n31659), .A2(n39463), .B1(n31723), .B2(n39457), .C1(
        n31595), .C2(n39451), .ZN(n35262) );
  AOI221_X1 U33581 ( .B1(n39726), .B2(n29398), .C1(n39720), .C2(n29462), .A(
        n34007), .ZN(n34002) );
  OAI222_X1 U33582 ( .A1(n31658), .A2(n39714), .B1(n31722), .B2(n39708), .C1(
        n31594), .C2(n39702), .ZN(n34007) );
  AOI221_X1 U33583 ( .B1(n39474), .B2(n29398), .C1(n39468), .C2(n29462), .A(
        n35281), .ZN(n35276) );
  OAI222_X1 U33584 ( .A1(n31658), .A2(n39462), .B1(n31722), .B2(n39456), .C1(
        n31594), .C2(n39450), .ZN(n35281) );
  AOI221_X1 U33585 ( .B1(n39726), .B2(n29397), .C1(n39720), .C2(n29461), .A(
        n34026), .ZN(n34021) );
  OAI222_X1 U33586 ( .A1(n31657), .A2(n39714), .B1(n31721), .B2(n39708), .C1(
        n31593), .C2(n39702), .ZN(n34026) );
  AOI221_X1 U33587 ( .B1(n39474), .B2(n29397), .C1(n39468), .C2(n29461), .A(
        n35300), .ZN(n35295) );
  OAI222_X1 U33588 ( .A1(n31657), .A2(n39462), .B1(n31721), .B2(n39456), .C1(
        n31593), .C2(n39450), .ZN(n35300) );
  AOI221_X1 U33589 ( .B1(n39726), .B2(n29396), .C1(n39720), .C2(n29460), .A(
        n34045), .ZN(n34040) );
  OAI222_X1 U33590 ( .A1(n31656), .A2(n39714), .B1(n31720), .B2(n39708), .C1(
        n31592), .C2(n39702), .ZN(n34045) );
  AOI221_X1 U33591 ( .B1(n39474), .B2(n29396), .C1(n39468), .C2(n29460), .A(
        n35319), .ZN(n35314) );
  OAI222_X1 U33592 ( .A1(n31656), .A2(n39462), .B1(n31720), .B2(n39456), .C1(
        n31592), .C2(n39450), .ZN(n35319) );
  AOI221_X1 U33593 ( .B1(n39726), .B2(n29395), .C1(n39720), .C2(n29459), .A(
        n34064), .ZN(n34059) );
  OAI222_X1 U33594 ( .A1(n31655), .A2(n39714), .B1(n31719), .B2(n39708), .C1(
        n31591), .C2(n39702), .ZN(n34064) );
  AOI221_X1 U33595 ( .B1(n39474), .B2(n29395), .C1(n39468), .C2(n29459), .A(
        n35338), .ZN(n35333) );
  OAI222_X1 U33596 ( .A1(n31655), .A2(n39462), .B1(n31719), .B2(n39456), .C1(
        n31591), .C2(n39450), .ZN(n35338) );
  AOI221_X1 U33597 ( .B1(n39726), .B2(n29394), .C1(n39720), .C2(n29458), .A(
        n34083), .ZN(n34078) );
  OAI222_X1 U33598 ( .A1(n31654), .A2(n39714), .B1(n31718), .B2(n39708), .C1(
        n31590), .C2(n39702), .ZN(n34083) );
  AOI221_X1 U33599 ( .B1(n39474), .B2(n29394), .C1(n39468), .C2(n29458), .A(
        n35357), .ZN(n35352) );
  OAI222_X1 U33600 ( .A1(n31654), .A2(n39462), .B1(n31718), .B2(n39456), .C1(
        n31590), .C2(n39450), .ZN(n35357) );
  AOI221_X1 U33601 ( .B1(n39726), .B2(n29393), .C1(n39720), .C2(n29457), .A(
        n34102), .ZN(n34097) );
  OAI222_X1 U33602 ( .A1(n31653), .A2(n39714), .B1(n31717), .B2(n39708), .C1(
        n31589), .C2(n39702), .ZN(n34102) );
  AOI221_X1 U33603 ( .B1(n39474), .B2(n29393), .C1(n39468), .C2(n29457), .A(
        n35376), .ZN(n35371) );
  OAI222_X1 U33604 ( .A1(n31653), .A2(n39462), .B1(n31717), .B2(n39456), .C1(
        n31589), .C2(n39450), .ZN(n35376) );
  AOI221_X1 U33605 ( .B1(n39726), .B2(n29392), .C1(n39720), .C2(n29456), .A(
        n34121), .ZN(n34116) );
  OAI222_X1 U33606 ( .A1(n31652), .A2(n39714), .B1(n31716), .B2(n39708), .C1(
        n31588), .C2(n39702), .ZN(n34121) );
  AOI221_X1 U33607 ( .B1(n39474), .B2(n29392), .C1(n39468), .C2(n29456), .A(
        n35395), .ZN(n35390) );
  OAI222_X1 U33608 ( .A1(n31652), .A2(n39462), .B1(n31716), .B2(n39456), .C1(
        n31588), .C2(n39450), .ZN(n35395) );
  AOI221_X1 U33609 ( .B1(n39726), .B2(n29391), .C1(n39720), .C2(n29455), .A(
        n34140), .ZN(n34135) );
  OAI222_X1 U33610 ( .A1(n31651), .A2(n39714), .B1(n31715), .B2(n39708), .C1(
        n31587), .C2(n39702), .ZN(n34140) );
  AOI221_X1 U33611 ( .B1(n39474), .B2(n29391), .C1(n39468), .C2(n29455), .A(
        n35414), .ZN(n35409) );
  OAI222_X1 U33612 ( .A1(n31651), .A2(n39462), .B1(n31715), .B2(n39456), .C1(
        n31587), .C2(n39450), .ZN(n35414) );
  AOI221_X1 U33613 ( .B1(n39726), .B2(n29390), .C1(n39720), .C2(n29454), .A(
        n34159), .ZN(n34154) );
  OAI222_X1 U33614 ( .A1(n31650), .A2(n39714), .B1(n31714), .B2(n39708), .C1(
        n31586), .C2(n39702), .ZN(n34159) );
  AOI221_X1 U33615 ( .B1(n39474), .B2(n29390), .C1(n39468), .C2(n29454), .A(
        n35433), .ZN(n35428) );
  OAI222_X1 U33616 ( .A1(n31650), .A2(n39462), .B1(n31714), .B2(n39456), .C1(
        n31586), .C2(n39450), .ZN(n35433) );
  AOI221_X1 U33617 ( .B1(n39726), .B2(n29389), .C1(n39720), .C2(n29453), .A(
        n34178), .ZN(n34173) );
  OAI222_X1 U33618 ( .A1(n31649), .A2(n39714), .B1(n31713), .B2(n39708), .C1(
        n31585), .C2(n39702), .ZN(n34178) );
  AOI221_X1 U33619 ( .B1(n39474), .B2(n29389), .C1(n39468), .C2(n29453), .A(
        n35452), .ZN(n35447) );
  OAI222_X1 U33620 ( .A1(n31649), .A2(n39462), .B1(n31713), .B2(n39456), .C1(
        n31585), .C2(n39450), .ZN(n35452) );
  AOI221_X1 U33621 ( .B1(n39726), .B2(n29388), .C1(n39720), .C2(n29452), .A(
        n34197), .ZN(n34192) );
  OAI222_X1 U33622 ( .A1(n31648), .A2(n39714), .B1(n31712), .B2(n39708), .C1(
        n31584), .C2(n39702), .ZN(n34197) );
  AOI221_X1 U33623 ( .B1(n39474), .B2(n29388), .C1(n39468), .C2(n29452), .A(
        n35471), .ZN(n35466) );
  OAI222_X1 U33624 ( .A1(n31648), .A2(n39462), .B1(n31712), .B2(n39456), .C1(
        n31584), .C2(n39450), .ZN(n35471) );
  AOI221_X1 U33625 ( .B1(n39726), .B2(n29387), .C1(n39720), .C2(n29451), .A(
        n34216), .ZN(n34211) );
  OAI222_X1 U33626 ( .A1(n31647), .A2(n39714), .B1(n31711), .B2(n39708), .C1(
        n31583), .C2(n39702), .ZN(n34216) );
  AOI221_X1 U33627 ( .B1(n39474), .B2(n29387), .C1(n39468), .C2(n29451), .A(
        n35490), .ZN(n35485) );
  OAI222_X1 U33628 ( .A1(n31647), .A2(n39462), .B1(n31711), .B2(n39456), .C1(
        n31583), .C2(n39450), .ZN(n35490) );
  AOI221_X1 U33629 ( .B1(n39725), .B2(n29386), .C1(n39719), .C2(n29450), .A(
        n34235), .ZN(n34230) );
  OAI222_X1 U33630 ( .A1(n31646), .A2(n39713), .B1(n31710), .B2(n39707), .C1(
        n31582), .C2(n39701), .ZN(n34235) );
  AOI221_X1 U33631 ( .B1(n39473), .B2(n29386), .C1(n39467), .C2(n29450), .A(
        n35509), .ZN(n35504) );
  OAI222_X1 U33632 ( .A1(n31646), .A2(n39461), .B1(n31710), .B2(n39455), .C1(
        n31582), .C2(n39449), .ZN(n35509) );
  AOI221_X1 U33633 ( .B1(n39725), .B2(n29385), .C1(n39719), .C2(n29449), .A(
        n34254), .ZN(n34249) );
  OAI222_X1 U33634 ( .A1(n31645), .A2(n39713), .B1(n31709), .B2(n39707), .C1(
        n31581), .C2(n39701), .ZN(n34254) );
  AOI221_X1 U33635 ( .B1(n39473), .B2(n29385), .C1(n39467), .C2(n29449), .A(
        n35528), .ZN(n35523) );
  OAI222_X1 U33636 ( .A1(n31645), .A2(n39461), .B1(n31709), .B2(n39455), .C1(
        n31581), .C2(n39449), .ZN(n35528) );
  AOI221_X1 U33637 ( .B1(n39725), .B2(n29384), .C1(n39719), .C2(n29448), .A(
        n34273), .ZN(n34268) );
  OAI222_X1 U33638 ( .A1(n31644), .A2(n39713), .B1(n31708), .B2(n39707), .C1(
        n31580), .C2(n39701), .ZN(n34273) );
  AOI221_X1 U33639 ( .B1(n39473), .B2(n29384), .C1(n39467), .C2(n29448), .A(
        n35547), .ZN(n35542) );
  OAI222_X1 U33640 ( .A1(n31644), .A2(n39461), .B1(n31708), .B2(n39455), .C1(
        n31580), .C2(n39449), .ZN(n35547) );
  AOI221_X1 U33641 ( .B1(n39725), .B2(n29383), .C1(n39719), .C2(n29447), .A(
        n34292), .ZN(n34287) );
  OAI222_X1 U33642 ( .A1(n31643), .A2(n39713), .B1(n31707), .B2(n39707), .C1(
        n31579), .C2(n39701), .ZN(n34292) );
  AOI221_X1 U33643 ( .B1(n39473), .B2(n29383), .C1(n39467), .C2(n29447), .A(
        n35566), .ZN(n35561) );
  OAI222_X1 U33644 ( .A1(n31643), .A2(n39461), .B1(n31707), .B2(n39455), .C1(
        n31579), .C2(n39449), .ZN(n35566) );
  AOI221_X1 U33645 ( .B1(n39725), .B2(n29382), .C1(n39719), .C2(n29446), .A(
        n34311), .ZN(n34306) );
  OAI222_X1 U33646 ( .A1(n31642), .A2(n39713), .B1(n31706), .B2(n39707), .C1(
        n31578), .C2(n39701), .ZN(n34311) );
  AOI221_X1 U33647 ( .B1(n39473), .B2(n29382), .C1(n39467), .C2(n29446), .A(
        n35585), .ZN(n35580) );
  OAI222_X1 U33648 ( .A1(n31642), .A2(n39461), .B1(n31706), .B2(n39455), .C1(
        n31578), .C2(n39449), .ZN(n35585) );
  AOI221_X1 U33649 ( .B1(n39725), .B2(n29381), .C1(n39719), .C2(n29445), .A(
        n34330), .ZN(n34325) );
  OAI222_X1 U33650 ( .A1(n31641), .A2(n39713), .B1(n31705), .B2(n39707), .C1(
        n31577), .C2(n39701), .ZN(n34330) );
  AOI221_X1 U33651 ( .B1(n39473), .B2(n29381), .C1(n39467), .C2(n29445), .A(
        n35604), .ZN(n35599) );
  OAI222_X1 U33652 ( .A1(n31641), .A2(n39461), .B1(n31705), .B2(n39455), .C1(
        n31577), .C2(n39449), .ZN(n35604) );
  AOI221_X1 U33653 ( .B1(n39725), .B2(n29380), .C1(n39719), .C2(n29444), .A(
        n34349), .ZN(n34344) );
  OAI222_X1 U33654 ( .A1(n31640), .A2(n39713), .B1(n31704), .B2(n39707), .C1(
        n31576), .C2(n39701), .ZN(n34349) );
  AOI221_X1 U33655 ( .B1(n39473), .B2(n29380), .C1(n39467), .C2(n29444), .A(
        n35623), .ZN(n35618) );
  OAI222_X1 U33656 ( .A1(n31640), .A2(n39461), .B1(n31704), .B2(n39455), .C1(
        n31576), .C2(n39449), .ZN(n35623) );
  AOI221_X1 U33657 ( .B1(n39725), .B2(n29379), .C1(n39719), .C2(n29443), .A(
        n34368), .ZN(n34363) );
  OAI222_X1 U33658 ( .A1(n31639), .A2(n39713), .B1(n31703), .B2(n39707), .C1(
        n31575), .C2(n39701), .ZN(n34368) );
  AOI221_X1 U33659 ( .B1(n39473), .B2(n29379), .C1(n39467), .C2(n29443), .A(
        n35642), .ZN(n35637) );
  OAI222_X1 U33660 ( .A1(n31639), .A2(n39461), .B1(n31703), .B2(n39455), .C1(
        n31575), .C2(n39449), .ZN(n35642) );
  AOI221_X1 U33661 ( .B1(n39725), .B2(n29378), .C1(n39719), .C2(n29442), .A(
        n34387), .ZN(n34382) );
  OAI222_X1 U33662 ( .A1(n31638), .A2(n39713), .B1(n31702), .B2(n39707), .C1(
        n31574), .C2(n39701), .ZN(n34387) );
  AOI221_X1 U33663 ( .B1(n39473), .B2(n29378), .C1(n39467), .C2(n29442), .A(
        n35661), .ZN(n35656) );
  OAI222_X1 U33664 ( .A1(n31638), .A2(n39461), .B1(n31702), .B2(n39455), .C1(
        n31574), .C2(n39449), .ZN(n35661) );
  AOI221_X1 U33665 ( .B1(n39725), .B2(n29377), .C1(n39719), .C2(n29441), .A(
        n34406), .ZN(n34401) );
  OAI222_X1 U33666 ( .A1(n31637), .A2(n39713), .B1(n31701), .B2(n39707), .C1(
        n31573), .C2(n39701), .ZN(n34406) );
  AOI221_X1 U33667 ( .B1(n39473), .B2(n29377), .C1(n39467), .C2(n29441), .A(
        n35680), .ZN(n35675) );
  OAI222_X1 U33668 ( .A1(n31637), .A2(n39461), .B1(n31701), .B2(n39455), .C1(
        n31573), .C2(n39449), .ZN(n35680) );
  AOI221_X1 U33669 ( .B1(n39725), .B2(n29376), .C1(n39719), .C2(n29440), .A(
        n34425), .ZN(n34420) );
  OAI222_X1 U33670 ( .A1(n31636), .A2(n39713), .B1(n31700), .B2(n39707), .C1(
        n31572), .C2(n39701), .ZN(n34425) );
  AOI221_X1 U33671 ( .B1(n39473), .B2(n29376), .C1(n39467), .C2(n29440), .A(
        n35699), .ZN(n35694) );
  OAI222_X1 U33672 ( .A1(n31636), .A2(n39461), .B1(n31700), .B2(n39455), .C1(
        n31572), .C2(n39449), .ZN(n35699) );
  AOI221_X1 U33673 ( .B1(n39725), .B2(n29375), .C1(n39719), .C2(n29439), .A(
        n34444), .ZN(n34439) );
  OAI222_X1 U33674 ( .A1(n31635), .A2(n39713), .B1(n31699), .B2(n39707), .C1(
        n31571), .C2(n39701), .ZN(n34444) );
  AOI221_X1 U33675 ( .B1(n39473), .B2(n29375), .C1(n39467), .C2(n29439), .A(
        n35718), .ZN(n35713) );
  OAI222_X1 U33676 ( .A1(n31635), .A2(n39461), .B1(n31699), .B2(n39455), .C1(
        n31571), .C2(n39449), .ZN(n35718) );
  AOI221_X1 U33677 ( .B1(n39724), .B2(n29374), .C1(n39718), .C2(n29438), .A(
        n34463), .ZN(n34458) );
  OAI222_X1 U33678 ( .A1(n31634), .A2(n39712), .B1(n31698), .B2(n39706), .C1(
        n31570), .C2(n39700), .ZN(n34463) );
  AOI221_X1 U33679 ( .B1(n39472), .B2(n29374), .C1(n39466), .C2(n29438), .A(
        n35737), .ZN(n35732) );
  OAI222_X1 U33680 ( .A1(n31634), .A2(n39460), .B1(n31698), .B2(n39454), .C1(
        n31570), .C2(n39448), .ZN(n35737) );
  AOI221_X1 U33681 ( .B1(n39724), .B2(n29373), .C1(n39718), .C2(n29437), .A(
        n34482), .ZN(n34477) );
  OAI222_X1 U33682 ( .A1(n31633), .A2(n39712), .B1(n31697), .B2(n39706), .C1(
        n31569), .C2(n39700), .ZN(n34482) );
  AOI221_X1 U33683 ( .B1(n39472), .B2(n29373), .C1(n39466), .C2(n29437), .A(
        n35756), .ZN(n35751) );
  OAI222_X1 U33684 ( .A1(n31633), .A2(n39460), .B1(n31697), .B2(n39454), .C1(
        n31569), .C2(n39448), .ZN(n35756) );
  AOI221_X1 U33685 ( .B1(n39724), .B2(n29372), .C1(n39718), .C2(n29436), .A(
        n34501), .ZN(n34496) );
  OAI222_X1 U33686 ( .A1(n31632), .A2(n39712), .B1(n31696), .B2(n39706), .C1(
        n31568), .C2(n39700), .ZN(n34501) );
  AOI221_X1 U33687 ( .B1(n39472), .B2(n29372), .C1(n39466), .C2(n29436), .A(
        n35775), .ZN(n35770) );
  OAI222_X1 U33688 ( .A1(n31632), .A2(n39460), .B1(n31696), .B2(n39454), .C1(
        n31568), .C2(n39448), .ZN(n35775) );
  AOI221_X1 U33689 ( .B1(n39724), .B2(n29371), .C1(n39718), .C2(n29435), .A(
        n34520), .ZN(n34515) );
  OAI222_X1 U33690 ( .A1(n31631), .A2(n39712), .B1(n31695), .B2(n39706), .C1(
        n31567), .C2(n39700), .ZN(n34520) );
  AOI221_X1 U33691 ( .B1(n39472), .B2(n29371), .C1(n39466), .C2(n29435), .A(
        n35794), .ZN(n35789) );
  OAI222_X1 U33692 ( .A1(n31631), .A2(n39460), .B1(n31695), .B2(n39454), .C1(
        n31567), .C2(n39448), .ZN(n35794) );
  AOI221_X1 U33693 ( .B1(n39724), .B2(n29370), .C1(n39718), .C2(n29434), .A(
        n34539), .ZN(n34534) );
  OAI222_X1 U33694 ( .A1(n31630), .A2(n39712), .B1(n31694), .B2(n39706), .C1(
        n31566), .C2(n39700), .ZN(n34539) );
  AOI221_X1 U33695 ( .B1(n39472), .B2(n29370), .C1(n39466), .C2(n29434), .A(
        n35813), .ZN(n35808) );
  OAI222_X1 U33696 ( .A1(n31630), .A2(n39460), .B1(n31694), .B2(n39454), .C1(
        n31566), .C2(n39448), .ZN(n35813) );
  AOI221_X1 U33697 ( .B1(n39724), .B2(n29369), .C1(n39718), .C2(n29433), .A(
        n34558), .ZN(n34553) );
  OAI222_X1 U33698 ( .A1(n31629), .A2(n39712), .B1(n31693), .B2(n39706), .C1(
        n31565), .C2(n39700), .ZN(n34558) );
  AOI221_X1 U33699 ( .B1(n39472), .B2(n29369), .C1(n39466), .C2(n29433), .A(
        n35832), .ZN(n35827) );
  OAI222_X1 U33700 ( .A1(n31629), .A2(n39460), .B1(n31693), .B2(n39454), .C1(
        n31565), .C2(n39448), .ZN(n35832) );
  AOI221_X1 U33701 ( .B1(n39724), .B2(n29368), .C1(n39718), .C2(n29432), .A(
        n34577), .ZN(n34572) );
  OAI222_X1 U33702 ( .A1(n31628), .A2(n39712), .B1(n31692), .B2(n39706), .C1(
        n31564), .C2(n39700), .ZN(n34577) );
  AOI221_X1 U33703 ( .B1(n39472), .B2(n29368), .C1(n39466), .C2(n29432), .A(
        n35851), .ZN(n35846) );
  OAI222_X1 U33704 ( .A1(n31628), .A2(n39460), .B1(n31692), .B2(n39454), .C1(
        n31564), .C2(n39448), .ZN(n35851) );
  AOI221_X1 U33705 ( .B1(n39724), .B2(n29367), .C1(n39718), .C2(n29431), .A(
        n34596), .ZN(n34591) );
  OAI222_X1 U33706 ( .A1(n31627), .A2(n39712), .B1(n31691), .B2(n39706), .C1(
        n31563), .C2(n39700), .ZN(n34596) );
  AOI221_X1 U33707 ( .B1(n39472), .B2(n29367), .C1(n39466), .C2(n29431), .A(
        n35870), .ZN(n35865) );
  OAI222_X1 U33708 ( .A1(n31627), .A2(n39460), .B1(n31691), .B2(n39454), .C1(
        n31563), .C2(n39448), .ZN(n35870) );
  AOI221_X1 U33709 ( .B1(n39724), .B2(n29366), .C1(n39718), .C2(n29430), .A(
        n34615), .ZN(n34610) );
  OAI222_X1 U33710 ( .A1(n31626), .A2(n39712), .B1(n31690), .B2(n39706), .C1(
        n31562), .C2(n39700), .ZN(n34615) );
  AOI221_X1 U33711 ( .B1(n39472), .B2(n29366), .C1(n39466), .C2(n29430), .A(
        n35889), .ZN(n35884) );
  OAI222_X1 U33712 ( .A1(n31626), .A2(n39460), .B1(n31690), .B2(n39454), .C1(
        n31562), .C2(n39448), .ZN(n35889) );
  AOI221_X1 U33713 ( .B1(n39724), .B2(n29365), .C1(n39718), .C2(n29429), .A(
        n34634), .ZN(n34629) );
  OAI222_X1 U33714 ( .A1(n31625), .A2(n39712), .B1(n31689), .B2(n39706), .C1(
        n31561), .C2(n39700), .ZN(n34634) );
  AOI221_X1 U33715 ( .B1(n39472), .B2(n29365), .C1(n39466), .C2(n29429), .A(
        n35908), .ZN(n35903) );
  OAI222_X1 U33716 ( .A1(n31625), .A2(n39460), .B1(n31689), .B2(n39454), .C1(
        n31561), .C2(n39448), .ZN(n35908) );
  AOI221_X1 U33717 ( .B1(n39724), .B2(n29364), .C1(n39718), .C2(n29428), .A(
        n34653), .ZN(n34648) );
  OAI222_X1 U33718 ( .A1(n31624), .A2(n39712), .B1(n31688), .B2(n39706), .C1(
        n31560), .C2(n39700), .ZN(n34653) );
  AOI221_X1 U33719 ( .B1(n39472), .B2(n29364), .C1(n39466), .C2(n29428), .A(
        n35927), .ZN(n35922) );
  OAI222_X1 U33720 ( .A1(n31624), .A2(n39460), .B1(n31688), .B2(n39454), .C1(
        n31560), .C2(n39448), .ZN(n35927) );
  AOI221_X1 U33721 ( .B1(n39724), .B2(n29363), .C1(n39718), .C2(n29427), .A(
        n34682), .ZN(n34667) );
  OAI222_X1 U33722 ( .A1(n31623), .A2(n39712), .B1(n31687), .B2(n39706), .C1(
        n31559), .C2(n39700), .ZN(n34682) );
  AOI221_X1 U33723 ( .B1(n39472), .B2(n29363), .C1(n39466), .C2(n29427), .A(
        n35956), .ZN(n35941) );
  OAI222_X1 U33724 ( .A1(n31623), .A2(n39460), .B1(n31687), .B2(n39454), .C1(
        n31559), .C2(n39448), .ZN(n35956) );
  AOI221_X1 U33725 ( .B1(n39072), .B2(n30469), .C1(n39066), .C2(n27996), .A(
        n37027), .ZN(n37020) );
  OAI222_X1 U33726 ( .A1(n30597), .A2(n39060), .B1(n30661), .B2(n39054), .C1(
        n30533), .C2(n39048), .ZN(n37027) );
  AOI221_X1 U33727 ( .B1(n39192), .B2(n29095), .C1(n39186), .C2(n29159), .A(
        n37019), .ZN(n37012) );
  OAI222_X1 U33728 ( .A1(n31483), .A2(n39180), .B1(n31547), .B2(n39174), .C1(
        n31419), .C2(n39168), .ZN(n37019) );
  AOI221_X1 U33729 ( .B1(n39073), .B2(n30468), .C1(n39067), .C2(n27995), .A(
        n37008), .ZN(n37001) );
  OAI222_X1 U33730 ( .A1(n30596), .A2(n39061), .B1(n30660), .B2(n39055), .C1(
        n30532), .C2(n39049), .ZN(n37008) );
  AOI221_X1 U33731 ( .B1(n39193), .B2(n29094), .C1(n39187), .C2(n29158), .A(
        n37000), .ZN(n36993) );
  OAI222_X1 U33732 ( .A1(n31482), .A2(n39181), .B1(n31546), .B2(n39175), .C1(
        n31418), .C2(n39169), .ZN(n37000) );
  AOI221_X1 U33733 ( .B1(n39073), .B2(n30467), .C1(n39067), .C2(n27994), .A(
        n36989), .ZN(n36982) );
  OAI222_X1 U33734 ( .A1(n30595), .A2(n39061), .B1(n30659), .B2(n39055), .C1(
        n30531), .C2(n39049), .ZN(n36989) );
  AOI221_X1 U33735 ( .B1(n39193), .B2(n29093), .C1(n39187), .C2(n29157), .A(
        n36981), .ZN(n36974) );
  OAI222_X1 U33736 ( .A1(n31481), .A2(n39181), .B1(n31545), .B2(n39175), .C1(
        n31417), .C2(n39169), .ZN(n36981) );
  AOI221_X1 U33737 ( .B1(n39073), .B2(n30466), .C1(n39067), .C2(n27993), .A(
        n36970), .ZN(n36963) );
  OAI222_X1 U33738 ( .A1(n30594), .A2(n39061), .B1(n30658), .B2(n39055), .C1(
        n30530), .C2(n39049), .ZN(n36970) );
  AOI221_X1 U33739 ( .B1(n39193), .B2(n29092), .C1(n39187), .C2(n29156), .A(
        n36962), .ZN(n36955) );
  OAI222_X1 U33740 ( .A1(n31480), .A2(n39181), .B1(n31544), .B2(n39175), .C1(
        n31416), .C2(n39169), .ZN(n36962) );
  AOI221_X1 U33741 ( .B1(n39073), .B2(n30465), .C1(n39067), .C2(n27992), .A(
        n36951), .ZN(n36944) );
  OAI222_X1 U33742 ( .A1(n30593), .A2(n39061), .B1(n30657), .B2(n39055), .C1(
        n30529), .C2(n39049), .ZN(n36951) );
  AOI221_X1 U33743 ( .B1(n39193), .B2(n29091), .C1(n39187), .C2(n29155), .A(
        n36943), .ZN(n36936) );
  OAI222_X1 U33744 ( .A1(n31479), .A2(n39181), .B1(n31543), .B2(n39175), .C1(
        n31415), .C2(n39169), .ZN(n36943) );
  AOI221_X1 U33745 ( .B1(n39073), .B2(n30464), .C1(n39067), .C2(n27991), .A(
        n36932), .ZN(n36925) );
  OAI222_X1 U33746 ( .A1(n30592), .A2(n39061), .B1(n30656), .B2(n39055), .C1(
        n30528), .C2(n39049), .ZN(n36932) );
  AOI221_X1 U33747 ( .B1(n39193), .B2(n29090), .C1(n39187), .C2(n29154), .A(
        n36924), .ZN(n36917) );
  OAI222_X1 U33748 ( .A1(n31478), .A2(n39181), .B1(n31542), .B2(n39175), .C1(
        n31414), .C2(n39169), .ZN(n36924) );
  AOI221_X1 U33749 ( .B1(n39073), .B2(n30463), .C1(n39067), .C2(n27990), .A(
        n36913), .ZN(n36906) );
  OAI222_X1 U33750 ( .A1(n30591), .A2(n39061), .B1(n30655), .B2(n39055), .C1(
        n30527), .C2(n39049), .ZN(n36913) );
  AOI221_X1 U33751 ( .B1(n39193), .B2(n29089), .C1(n39187), .C2(n29153), .A(
        n36905), .ZN(n36898) );
  OAI222_X1 U33752 ( .A1(n31477), .A2(n39181), .B1(n31541), .B2(n39175), .C1(
        n31413), .C2(n39169), .ZN(n36905) );
  AOI221_X1 U33753 ( .B1(n39073), .B2(n30462), .C1(n39067), .C2(n27989), .A(
        n36894), .ZN(n36887) );
  OAI222_X1 U33754 ( .A1(n30590), .A2(n39061), .B1(n30654), .B2(n39055), .C1(
        n30526), .C2(n39049), .ZN(n36894) );
  AOI221_X1 U33755 ( .B1(n39193), .B2(n29088), .C1(n39187), .C2(n29152), .A(
        n36886), .ZN(n36879) );
  OAI222_X1 U33756 ( .A1(n31476), .A2(n39181), .B1(n31540), .B2(n39175), .C1(
        n31412), .C2(n39169), .ZN(n36886) );
  AOI221_X1 U33757 ( .B1(n39073), .B2(n30461), .C1(n39067), .C2(n27988), .A(
        n36875), .ZN(n36868) );
  OAI222_X1 U33758 ( .A1(n30589), .A2(n39061), .B1(n30653), .B2(n39055), .C1(
        n30525), .C2(n39049), .ZN(n36875) );
  AOI221_X1 U33759 ( .B1(n39193), .B2(n29087), .C1(n39187), .C2(n29151), .A(
        n36867), .ZN(n36860) );
  OAI222_X1 U33760 ( .A1(n31475), .A2(n39181), .B1(n31539), .B2(n39175), .C1(
        n31411), .C2(n39169), .ZN(n36867) );
  AOI221_X1 U33761 ( .B1(n39073), .B2(n30460), .C1(n39067), .C2(n27987), .A(
        n36856), .ZN(n36849) );
  OAI222_X1 U33762 ( .A1(n30588), .A2(n39061), .B1(n30652), .B2(n39055), .C1(
        n30524), .C2(n39049), .ZN(n36856) );
  AOI221_X1 U33763 ( .B1(n39193), .B2(n29086), .C1(n39187), .C2(n29150), .A(
        n36848), .ZN(n36841) );
  OAI222_X1 U33764 ( .A1(n31474), .A2(n39181), .B1(n31538), .B2(n39175), .C1(
        n31410), .C2(n39169), .ZN(n36848) );
  AOI221_X1 U33765 ( .B1(n39073), .B2(n30459), .C1(n39067), .C2(n27986), .A(
        n36837), .ZN(n36830) );
  OAI222_X1 U33766 ( .A1(n30587), .A2(n39061), .B1(n30651), .B2(n39055), .C1(
        n30523), .C2(n39049), .ZN(n36837) );
  AOI221_X1 U33767 ( .B1(n39193), .B2(n29085), .C1(n39187), .C2(n29149), .A(
        n36829), .ZN(n36822) );
  OAI222_X1 U33768 ( .A1(n31473), .A2(n39181), .B1(n31537), .B2(n39175), .C1(
        n31409), .C2(n39169), .ZN(n36829) );
  AOI221_X1 U33769 ( .B1(n39073), .B2(n30458), .C1(n39067), .C2(n27985), .A(
        n36818), .ZN(n36811) );
  OAI222_X1 U33770 ( .A1(n30586), .A2(n39061), .B1(n30650), .B2(n39055), .C1(
        n30522), .C2(n39049), .ZN(n36818) );
  AOI221_X1 U33771 ( .B1(n39193), .B2(n29084), .C1(n39187), .C2(n29148), .A(
        n36810), .ZN(n36803) );
  OAI222_X1 U33772 ( .A1(n31472), .A2(n39181), .B1(n31536), .B2(n39175), .C1(
        n31408), .C2(n39169), .ZN(n36810) );
  AOI221_X1 U33773 ( .B1(n39073), .B2(n32546), .C1(n39067), .C2(n27984), .A(
        n36799), .ZN(n36792) );
  OAI222_X1 U33774 ( .A1(n30585), .A2(n39061), .B1(n30649), .B2(n39055), .C1(
        n30521), .C2(n39049), .ZN(n36799) );
  AOI221_X1 U33775 ( .B1(n39193), .B2(n29083), .C1(n39187), .C2(n29147), .A(
        n36791), .ZN(n36784) );
  OAI222_X1 U33776 ( .A1(n31471), .A2(n39181), .B1(n31535), .B2(n39175), .C1(
        n31407), .C2(n39169), .ZN(n36791) );
  AOI221_X1 U33777 ( .B1(n39074), .B2(n32545), .C1(n39068), .C2(n27983), .A(
        n36780), .ZN(n36773) );
  OAI222_X1 U33778 ( .A1(n30584), .A2(n39062), .B1(n30648), .B2(n39056), .C1(
        n30520), .C2(n39050), .ZN(n36780) );
  AOI221_X1 U33779 ( .B1(n39194), .B2(n29082), .C1(n39188), .C2(n29146), .A(
        n36772), .ZN(n36765) );
  OAI222_X1 U33780 ( .A1(n31470), .A2(n39182), .B1(n31534), .B2(n39176), .C1(
        n31406), .C2(n39170), .ZN(n36772) );
  AOI221_X1 U33781 ( .B1(n39074), .B2(n32544), .C1(n39068), .C2(n27982), .A(
        n36761), .ZN(n36754) );
  OAI222_X1 U33782 ( .A1(n30583), .A2(n39062), .B1(n30647), .B2(n39056), .C1(
        n30519), .C2(n39050), .ZN(n36761) );
  AOI221_X1 U33783 ( .B1(n39194), .B2(n29081), .C1(n39188), .C2(n29145), .A(
        n36753), .ZN(n36746) );
  OAI222_X1 U33784 ( .A1(n31469), .A2(n39182), .B1(n31533), .B2(n39176), .C1(
        n31405), .C2(n39170), .ZN(n36753) );
  AOI221_X1 U33785 ( .B1(n39074), .B2(n32543), .C1(n39068), .C2(n27981), .A(
        n36742), .ZN(n36735) );
  OAI222_X1 U33786 ( .A1(n30582), .A2(n39062), .B1(n30646), .B2(n39056), .C1(
        n30518), .C2(n39050), .ZN(n36742) );
  AOI221_X1 U33787 ( .B1(n39194), .B2(n29080), .C1(n39188), .C2(n29144), .A(
        n36734), .ZN(n36727) );
  OAI222_X1 U33788 ( .A1(n31468), .A2(n39182), .B1(n31532), .B2(n39176), .C1(
        n31404), .C2(n39170), .ZN(n36734) );
  AOI221_X1 U33789 ( .B1(n39074), .B2(n32542), .C1(n39068), .C2(n27980), .A(
        n36723), .ZN(n36716) );
  OAI222_X1 U33790 ( .A1(n30581), .A2(n39062), .B1(n30645), .B2(n39056), .C1(
        n30517), .C2(n39050), .ZN(n36723) );
  AOI221_X1 U33791 ( .B1(n39194), .B2(n29079), .C1(n39188), .C2(n29143), .A(
        n36715), .ZN(n36708) );
  OAI222_X1 U33792 ( .A1(n31467), .A2(n39182), .B1(n31531), .B2(n39176), .C1(
        n31403), .C2(n39170), .ZN(n36715) );
  AOI221_X1 U33793 ( .B1(n39074), .B2(n32541), .C1(n39068), .C2(n27979), .A(
        n36704), .ZN(n36697) );
  OAI222_X1 U33794 ( .A1(n30580), .A2(n39062), .B1(n30644), .B2(n39056), .C1(
        n30516), .C2(n39050), .ZN(n36704) );
  AOI221_X1 U33795 ( .B1(n39194), .B2(n29078), .C1(n39188), .C2(n29142), .A(
        n36696), .ZN(n36689) );
  OAI222_X1 U33796 ( .A1(n31466), .A2(n39182), .B1(n31530), .B2(n39176), .C1(
        n31402), .C2(n39170), .ZN(n36696) );
  AOI221_X1 U33797 ( .B1(n39074), .B2(n32540), .C1(n39068), .C2(n27978), .A(
        n36685), .ZN(n36678) );
  OAI222_X1 U33798 ( .A1(n30579), .A2(n39062), .B1(n30643), .B2(n39056), .C1(
        n30515), .C2(n39050), .ZN(n36685) );
  AOI221_X1 U33799 ( .B1(n39194), .B2(n29077), .C1(n39188), .C2(n29141), .A(
        n36677), .ZN(n36670) );
  OAI222_X1 U33800 ( .A1(n31465), .A2(n39182), .B1(n31529), .B2(n39176), .C1(
        n31401), .C2(n39170), .ZN(n36677) );
  AOI221_X1 U33801 ( .B1(n39074), .B2(n32539), .C1(n39068), .C2(n27977), .A(
        n36666), .ZN(n36659) );
  OAI222_X1 U33802 ( .A1(n30578), .A2(n39062), .B1(n30642), .B2(n39056), .C1(
        n30514), .C2(n39050), .ZN(n36666) );
  AOI221_X1 U33803 ( .B1(n39194), .B2(n29076), .C1(n39188), .C2(n29140), .A(
        n36658), .ZN(n36651) );
  OAI222_X1 U33804 ( .A1(n31464), .A2(n39182), .B1(n31528), .B2(n39176), .C1(
        n31400), .C2(n39170), .ZN(n36658) );
  AOI221_X1 U33805 ( .B1(n39074), .B2(n32538), .C1(n39068), .C2(n27976), .A(
        n36647), .ZN(n36640) );
  OAI222_X1 U33806 ( .A1(n30577), .A2(n39062), .B1(n30641), .B2(n39056), .C1(
        n30513), .C2(n39050), .ZN(n36647) );
  AOI221_X1 U33807 ( .B1(n39194), .B2(n29075), .C1(n39188), .C2(n29139), .A(
        n36639), .ZN(n36632) );
  OAI222_X1 U33808 ( .A1(n31463), .A2(n39182), .B1(n31527), .B2(n39176), .C1(
        n31399), .C2(n39170), .ZN(n36639) );
  AOI221_X1 U33809 ( .B1(n39074), .B2(n32537), .C1(n39068), .C2(n27975), .A(
        n36628), .ZN(n36621) );
  OAI222_X1 U33810 ( .A1(n30576), .A2(n39062), .B1(n30640), .B2(n39056), .C1(
        n30512), .C2(n39050), .ZN(n36628) );
  AOI221_X1 U33811 ( .B1(n39194), .B2(n29074), .C1(n39188), .C2(n29138), .A(
        n36620), .ZN(n36613) );
  OAI222_X1 U33812 ( .A1(n31462), .A2(n39182), .B1(n31526), .B2(n39176), .C1(
        n31398), .C2(n39170), .ZN(n36620) );
  AOI221_X1 U33813 ( .B1(n39074), .B2(n32536), .C1(n39068), .C2(n27974), .A(
        n36609), .ZN(n36602) );
  OAI222_X1 U33814 ( .A1(n30575), .A2(n39062), .B1(n30639), .B2(n39056), .C1(
        n30511), .C2(n39050), .ZN(n36609) );
  AOI221_X1 U33815 ( .B1(n39194), .B2(n29073), .C1(n39188), .C2(n29137), .A(
        n36601), .ZN(n36594) );
  OAI222_X1 U33816 ( .A1(n31461), .A2(n39182), .B1(n31525), .B2(n39176), .C1(
        n31397), .C2(n39170), .ZN(n36601) );
  AOI221_X1 U33817 ( .B1(n39074), .B2(n32535), .C1(n39068), .C2(n27973), .A(
        n36590), .ZN(n36583) );
  OAI222_X1 U33818 ( .A1(n30574), .A2(n39062), .B1(n30638), .B2(n39056), .C1(
        n30510), .C2(n39050), .ZN(n36590) );
  AOI221_X1 U33819 ( .B1(n39194), .B2(n29072), .C1(n39188), .C2(n29136), .A(
        n36582), .ZN(n36575) );
  OAI222_X1 U33820 ( .A1(n31460), .A2(n39182), .B1(n31524), .B2(n39176), .C1(
        n31396), .C2(n39170), .ZN(n36582) );
  AOI221_X1 U33821 ( .B1(n39074), .B2(n32534), .C1(n39068), .C2(n27972), .A(
        n36571), .ZN(n36564) );
  OAI222_X1 U33822 ( .A1(n30573), .A2(n39062), .B1(n30637), .B2(n39056), .C1(
        n30509), .C2(n39050), .ZN(n36571) );
  AOI221_X1 U33823 ( .B1(n39194), .B2(n29071), .C1(n39188), .C2(n29135), .A(
        n36563), .ZN(n36556) );
  OAI222_X1 U33824 ( .A1(n31459), .A2(n39182), .B1(n31523), .B2(n39176), .C1(
        n31395), .C2(n39170), .ZN(n36563) );
  AOI221_X1 U33825 ( .B1(n39075), .B2(n32533), .C1(n39069), .C2(n27971), .A(
        n36552), .ZN(n36545) );
  OAI222_X1 U33826 ( .A1(n30572), .A2(n39063), .B1(n30636), .B2(n39057), .C1(
        n30508), .C2(n39051), .ZN(n36552) );
  AOI221_X1 U33827 ( .B1(n39195), .B2(n29070), .C1(n39189), .C2(n29134), .A(
        n36544), .ZN(n36537) );
  OAI222_X1 U33828 ( .A1(n31458), .A2(n39183), .B1(n31522), .B2(n39177), .C1(
        n31394), .C2(n39171), .ZN(n36544) );
  AOI221_X1 U33829 ( .B1(n39075), .B2(n32532), .C1(n39069), .C2(n27970), .A(
        n36533), .ZN(n36526) );
  OAI222_X1 U33830 ( .A1(n30571), .A2(n39063), .B1(n30635), .B2(n39057), .C1(
        n30507), .C2(n39051), .ZN(n36533) );
  AOI221_X1 U33831 ( .B1(n39195), .B2(n29069), .C1(n39189), .C2(n29133), .A(
        n36525), .ZN(n36518) );
  OAI222_X1 U33832 ( .A1(n31457), .A2(n39183), .B1(n31521), .B2(n39177), .C1(
        n31393), .C2(n39171), .ZN(n36525) );
  AOI221_X1 U33833 ( .B1(n39075), .B2(n32531), .C1(n39069), .C2(n27969), .A(
        n36514), .ZN(n36507) );
  OAI222_X1 U33834 ( .A1(n30570), .A2(n39063), .B1(n30634), .B2(n39057), .C1(
        n30506), .C2(n39051), .ZN(n36514) );
  AOI221_X1 U33835 ( .B1(n39195), .B2(n29068), .C1(n39189), .C2(n29132), .A(
        n36506), .ZN(n36499) );
  OAI222_X1 U33836 ( .A1(n31456), .A2(n39183), .B1(n31520), .B2(n39177), .C1(
        n31392), .C2(n39171), .ZN(n36506) );
  AOI221_X1 U33837 ( .B1(n39075), .B2(n32530), .C1(n39069), .C2(n27968), .A(
        n36495), .ZN(n36488) );
  OAI222_X1 U33838 ( .A1(n30569), .A2(n39063), .B1(n30633), .B2(n39057), .C1(
        n30505), .C2(n39051), .ZN(n36495) );
  AOI221_X1 U33839 ( .B1(n39195), .B2(n29067), .C1(n39189), .C2(n29131), .A(
        n36487), .ZN(n36480) );
  OAI222_X1 U33840 ( .A1(n31455), .A2(n39183), .B1(n31519), .B2(n39177), .C1(
        n31391), .C2(n39171), .ZN(n36487) );
  AOI221_X1 U33841 ( .B1(n39075), .B2(n32529), .C1(n39069), .C2(n27967), .A(
        n36476), .ZN(n36469) );
  OAI222_X1 U33842 ( .A1(n30568), .A2(n39063), .B1(n30632), .B2(n39057), .C1(
        n30504), .C2(n39051), .ZN(n36476) );
  AOI221_X1 U33843 ( .B1(n39195), .B2(n29066), .C1(n39189), .C2(n29130), .A(
        n36468), .ZN(n36461) );
  OAI222_X1 U33844 ( .A1(n31454), .A2(n39183), .B1(n31518), .B2(n39177), .C1(
        n31390), .C2(n39171), .ZN(n36468) );
  AOI221_X1 U33845 ( .B1(n39075), .B2(n32528), .C1(n39069), .C2(n27966), .A(
        n36457), .ZN(n36450) );
  OAI222_X1 U33846 ( .A1(n30567), .A2(n39063), .B1(n30631), .B2(n39057), .C1(
        n30503), .C2(n39051), .ZN(n36457) );
  AOI221_X1 U33847 ( .B1(n39195), .B2(n29065), .C1(n39189), .C2(n29129), .A(
        n36449), .ZN(n36442) );
  OAI222_X1 U33848 ( .A1(n31453), .A2(n39183), .B1(n31517), .B2(n39177), .C1(
        n31389), .C2(n39171), .ZN(n36449) );
  AOI221_X1 U33849 ( .B1(n39075), .B2(n32527), .C1(n39069), .C2(n27965), .A(
        n36438), .ZN(n36431) );
  OAI222_X1 U33850 ( .A1(n30566), .A2(n39063), .B1(n30630), .B2(n39057), .C1(
        n30502), .C2(n39051), .ZN(n36438) );
  AOI221_X1 U33851 ( .B1(n39195), .B2(n29064), .C1(n39189), .C2(n29128), .A(
        n36430), .ZN(n36423) );
  OAI222_X1 U33852 ( .A1(n31452), .A2(n39183), .B1(n31516), .B2(n39177), .C1(
        n31388), .C2(n39171), .ZN(n36430) );
  AOI221_X1 U33853 ( .B1(n39075), .B2(n32526), .C1(n39069), .C2(n27964), .A(
        n36419), .ZN(n36412) );
  OAI222_X1 U33854 ( .A1(n30565), .A2(n39063), .B1(n30629), .B2(n39057), .C1(
        n30501), .C2(n39051), .ZN(n36419) );
  AOI221_X1 U33855 ( .B1(n39195), .B2(n29063), .C1(n39189), .C2(n29127), .A(
        n36411), .ZN(n36404) );
  OAI222_X1 U33856 ( .A1(n31451), .A2(n39183), .B1(n31515), .B2(n39177), .C1(
        n31387), .C2(n39171), .ZN(n36411) );
  AOI221_X1 U33857 ( .B1(n39075), .B2(n32525), .C1(n39069), .C2(n27963), .A(
        n36400), .ZN(n36393) );
  OAI222_X1 U33858 ( .A1(n30564), .A2(n39063), .B1(n30628), .B2(n39057), .C1(
        n30500), .C2(n39051), .ZN(n36400) );
  AOI221_X1 U33859 ( .B1(n39195), .B2(n29062), .C1(n39189), .C2(n29126), .A(
        n36392), .ZN(n36385) );
  OAI222_X1 U33860 ( .A1(n31450), .A2(n39183), .B1(n31514), .B2(n39177), .C1(
        n31386), .C2(n39171), .ZN(n36392) );
  AOI221_X1 U33861 ( .B1(n39075), .B2(n32524), .C1(n39069), .C2(n27962), .A(
        n36381), .ZN(n36374) );
  OAI222_X1 U33862 ( .A1(n30563), .A2(n39063), .B1(n30627), .B2(n39057), .C1(
        n30499), .C2(n39051), .ZN(n36381) );
  AOI221_X1 U33863 ( .B1(n39195), .B2(n29061), .C1(n39189), .C2(n29125), .A(
        n36373), .ZN(n36366) );
  OAI222_X1 U33864 ( .A1(n31449), .A2(n39183), .B1(n31513), .B2(n39177), .C1(
        n31385), .C2(n39171), .ZN(n36373) );
  AOI221_X1 U33865 ( .B1(n39075), .B2(n32523), .C1(n39069), .C2(n27961), .A(
        n36362), .ZN(n36355) );
  OAI222_X1 U33866 ( .A1(n30562), .A2(n39063), .B1(n30626), .B2(n39057), .C1(
        n30498), .C2(n39051), .ZN(n36362) );
  AOI221_X1 U33867 ( .B1(n39195), .B2(n29060), .C1(n39189), .C2(n29124), .A(
        n36354), .ZN(n36347) );
  OAI222_X1 U33868 ( .A1(n31448), .A2(n39183), .B1(n31512), .B2(n39177), .C1(
        n31384), .C2(n39171), .ZN(n36354) );
  AOI221_X1 U33869 ( .B1(n39075), .B2(n32522), .C1(n39069), .C2(n27960), .A(
        n36343), .ZN(n36336) );
  OAI222_X1 U33870 ( .A1(n30561), .A2(n39063), .B1(n30625), .B2(n39057), .C1(
        n30497), .C2(n39051), .ZN(n36343) );
  AOI221_X1 U33871 ( .B1(n39195), .B2(n29059), .C1(n39189), .C2(n29123), .A(
        n36335), .ZN(n36328) );
  OAI222_X1 U33872 ( .A1(n31447), .A2(n39183), .B1(n31511), .B2(n39177), .C1(
        n31383), .C2(n39171), .ZN(n36335) );
  AOI221_X1 U33873 ( .B1(n39076), .B2(n32521), .C1(n39070), .C2(n27959), .A(
        n36324), .ZN(n36317) );
  OAI222_X1 U33874 ( .A1(n30560), .A2(n39064), .B1(n30624), .B2(n39058), .C1(
        n30496), .C2(n39052), .ZN(n36324) );
  AOI221_X1 U33875 ( .B1(n39196), .B2(n29058), .C1(n39190), .C2(n29122), .A(
        n36316), .ZN(n36309) );
  OAI222_X1 U33876 ( .A1(n31446), .A2(n39184), .B1(n31510), .B2(n39178), .C1(
        n31382), .C2(n39172), .ZN(n36316) );
  AOI221_X1 U33877 ( .B1(n39076), .B2(n32520), .C1(n39070), .C2(n27958), .A(
        n36305), .ZN(n36298) );
  OAI222_X1 U33878 ( .A1(n30559), .A2(n39064), .B1(n30623), .B2(n39058), .C1(
        n30495), .C2(n39052), .ZN(n36305) );
  AOI221_X1 U33879 ( .B1(n39196), .B2(n29057), .C1(n39190), .C2(n29121), .A(
        n36297), .ZN(n36290) );
  OAI222_X1 U33880 ( .A1(n31445), .A2(n39184), .B1(n31509), .B2(n39178), .C1(
        n31381), .C2(n39172), .ZN(n36297) );
  AOI221_X1 U33881 ( .B1(n39076), .B2(n32519), .C1(n39070), .C2(n27957), .A(
        n36286), .ZN(n36279) );
  OAI222_X1 U33882 ( .A1(n30558), .A2(n39064), .B1(n30622), .B2(n39058), .C1(
        n30494), .C2(n39052), .ZN(n36286) );
  AOI221_X1 U33883 ( .B1(n39196), .B2(n29056), .C1(n39190), .C2(n29120), .A(
        n36278), .ZN(n36271) );
  OAI222_X1 U33884 ( .A1(n31444), .A2(n39184), .B1(n31508), .B2(n39178), .C1(
        n31380), .C2(n39172), .ZN(n36278) );
  AOI221_X1 U33885 ( .B1(n39076), .B2(n32518), .C1(n39070), .C2(n27956), .A(
        n36267), .ZN(n36260) );
  OAI222_X1 U33886 ( .A1(n30557), .A2(n39064), .B1(n30621), .B2(n39058), .C1(
        n30493), .C2(n39052), .ZN(n36267) );
  AOI221_X1 U33887 ( .B1(n39196), .B2(n29055), .C1(n39190), .C2(n29119), .A(
        n36259), .ZN(n36252) );
  OAI222_X1 U33888 ( .A1(n31443), .A2(n39184), .B1(n31507), .B2(n39178), .C1(
        n31379), .C2(n39172), .ZN(n36259) );
  AOI221_X1 U33889 ( .B1(n39076), .B2(n32517), .C1(n39070), .C2(n27955), .A(
        n36248), .ZN(n36241) );
  OAI222_X1 U33890 ( .A1(n30556), .A2(n39064), .B1(n30620), .B2(n39058), .C1(
        n30492), .C2(n39052), .ZN(n36248) );
  AOI221_X1 U33891 ( .B1(n39196), .B2(n29054), .C1(n39190), .C2(n29118), .A(
        n36240), .ZN(n36233) );
  OAI222_X1 U33892 ( .A1(n31442), .A2(n39184), .B1(n31506), .B2(n39178), .C1(
        n31378), .C2(n39172), .ZN(n36240) );
  AOI221_X1 U33893 ( .B1(n39076), .B2(n32516), .C1(n39070), .C2(n27954), .A(
        n36229), .ZN(n36222) );
  OAI222_X1 U33894 ( .A1(n30555), .A2(n39064), .B1(n30619), .B2(n39058), .C1(
        n30491), .C2(n39052), .ZN(n36229) );
  AOI221_X1 U33895 ( .B1(n39196), .B2(n29053), .C1(n39190), .C2(n29117), .A(
        n36221), .ZN(n36214) );
  OAI222_X1 U33896 ( .A1(n31441), .A2(n39184), .B1(n31505), .B2(n39178), .C1(
        n31377), .C2(n39172), .ZN(n36221) );
  AOI221_X1 U33897 ( .B1(n39072), .B2(n30479), .C1(n39066), .C2(n28006), .A(
        n37217), .ZN(n37210) );
  OAI222_X1 U33898 ( .A1(n30607), .A2(n39060), .B1(n30671), .B2(n39054), .C1(
        n30543), .C2(n39048), .ZN(n37217) );
  AOI221_X1 U33899 ( .B1(n39192), .B2(n29105), .C1(n39186), .C2(n29169), .A(
        n37209), .ZN(n37202) );
  OAI222_X1 U33900 ( .A1(n31493), .A2(n39180), .B1(n31557), .B2(n39174), .C1(
        n31429), .C2(n39168), .ZN(n37209) );
  AOI221_X1 U33901 ( .B1(n39072), .B2(n30478), .C1(n39066), .C2(n28005), .A(
        n37198), .ZN(n37191) );
  OAI222_X1 U33902 ( .A1(n30606), .A2(n39060), .B1(n30670), .B2(n39054), .C1(
        n30542), .C2(n39048), .ZN(n37198) );
  AOI221_X1 U33903 ( .B1(n39192), .B2(n29104), .C1(n39186), .C2(n29168), .A(
        n37190), .ZN(n37183) );
  OAI222_X1 U33904 ( .A1(n31492), .A2(n39180), .B1(n31556), .B2(n39174), .C1(
        n31428), .C2(n39168), .ZN(n37190) );
  AOI221_X1 U33905 ( .B1(n39072), .B2(n30477), .C1(n39066), .C2(n28004), .A(
        n37179), .ZN(n37172) );
  OAI222_X1 U33906 ( .A1(n30605), .A2(n39060), .B1(n30669), .B2(n39054), .C1(
        n30541), .C2(n39048), .ZN(n37179) );
  AOI221_X1 U33907 ( .B1(n39192), .B2(n29103), .C1(n39186), .C2(n29167), .A(
        n37171), .ZN(n37164) );
  OAI222_X1 U33908 ( .A1(n31491), .A2(n39180), .B1(n31555), .B2(n39174), .C1(
        n31427), .C2(n39168), .ZN(n37171) );
  AOI221_X1 U33909 ( .B1(n39072), .B2(n30476), .C1(n39066), .C2(n28003), .A(
        n37160), .ZN(n37153) );
  OAI222_X1 U33910 ( .A1(n30604), .A2(n39060), .B1(n30668), .B2(n39054), .C1(
        n30540), .C2(n39048), .ZN(n37160) );
  AOI221_X1 U33911 ( .B1(n39192), .B2(n29102), .C1(n39186), .C2(n29166), .A(
        n37152), .ZN(n37145) );
  OAI222_X1 U33912 ( .A1(n31490), .A2(n39180), .B1(n31554), .B2(n39174), .C1(
        n31426), .C2(n39168), .ZN(n37152) );
  AOI221_X1 U33913 ( .B1(n39072), .B2(n30475), .C1(n39066), .C2(n28002), .A(
        n37141), .ZN(n37134) );
  OAI222_X1 U33914 ( .A1(n30603), .A2(n39060), .B1(n30667), .B2(n39054), .C1(
        n30539), .C2(n39048), .ZN(n37141) );
  AOI221_X1 U33915 ( .B1(n39192), .B2(n29101), .C1(n39186), .C2(n29165), .A(
        n37133), .ZN(n37126) );
  OAI222_X1 U33916 ( .A1(n31489), .A2(n39180), .B1(n31553), .B2(n39174), .C1(
        n31425), .C2(n39168), .ZN(n37133) );
  AOI221_X1 U33917 ( .B1(n39077), .B2(n32507), .C1(n39071), .C2(n27947), .A(
        n36096), .ZN(n36089) );
  OAI222_X1 U33918 ( .A1(n30548), .A2(n39065), .B1(n30612), .B2(n39059), .C1(
        n30484), .C2(n39053), .ZN(n36096) );
  AOI221_X1 U33919 ( .B1(n39197), .B2(n29046), .C1(n39191), .C2(n29110), .A(
        n36088), .ZN(n36081) );
  OAI222_X1 U33920 ( .A1(n31434), .A2(n39185), .B1(n31498), .B2(n39179), .C1(
        n31370), .C2(n39173), .ZN(n36088) );
  AOI221_X1 U33921 ( .B1(n39077), .B2(n32506), .C1(n39071), .C2(n27946), .A(
        n36077), .ZN(n36070) );
  OAI222_X1 U33922 ( .A1(n30547), .A2(n39065), .B1(n30611), .B2(n39059), .C1(
        n30483), .C2(n39053), .ZN(n36077) );
  AOI221_X1 U33923 ( .B1(n39197), .B2(n29045), .C1(n39191), .C2(n29109), .A(
        n36069), .ZN(n36062) );
  OAI222_X1 U33924 ( .A1(n31433), .A2(n39185), .B1(n31497), .B2(n39179), .C1(
        n31369), .C2(n39173), .ZN(n36069) );
  AOI221_X1 U33925 ( .B1(n39077), .B2(n32509), .C1(n39071), .C2(n27945), .A(
        n36058), .ZN(n36051) );
  OAI222_X1 U33926 ( .A1(n30546), .A2(n39065), .B1(n30610), .B2(n39059), .C1(
        n30482), .C2(n39053), .ZN(n36058) );
  AOI221_X1 U33927 ( .B1(n39197), .B2(n29044), .C1(n39191), .C2(n29108), .A(
        n36050), .ZN(n36043) );
  OAI222_X1 U33928 ( .A1(n31432), .A2(n39185), .B1(n31496), .B2(n39179), .C1(
        n31368), .C2(n39173), .ZN(n36050) );
  AOI221_X1 U33929 ( .B1(n39077), .B2(n32508), .C1(n39071), .C2(n27944), .A(
        n36036), .ZN(n36012) );
  OAI222_X1 U33930 ( .A1(n30545), .A2(n39065), .B1(n30609), .B2(n39059), .C1(
        n30481), .C2(n39053), .ZN(n36036) );
  AOI221_X1 U33931 ( .B1(n39197), .B2(n29043), .C1(n39191), .C2(n29107), .A(
        n36008), .ZN(n35984) );
  OAI222_X1 U33932 ( .A1(n31431), .A2(n39185), .B1(n31495), .B2(n39179), .C1(
        n31367), .C2(n39173), .ZN(n36008) );
  AOI221_X1 U33933 ( .B1(n39072), .B2(n30480), .C1(n39066), .C2(n28007), .A(
        n37250), .ZN(n37241) );
  OAI222_X1 U33934 ( .A1(n30608), .A2(n39060), .B1(n30672), .B2(n39054), .C1(
        n30544), .C2(n39048), .ZN(n37250) );
  AOI221_X1 U33935 ( .B1(n39192), .B2(n29106), .C1(n39186), .C2(n29170), .A(
        n37238), .ZN(n37221) );
  OAI222_X1 U33936 ( .A1(n31494), .A2(n39180), .B1(n31558), .B2(n39174), .C1(
        n31430), .C2(n39168), .ZN(n37238) );
  AOI221_X1 U33937 ( .B1(n39072), .B2(n30474), .C1(n39066), .C2(n28001), .A(
        n37122), .ZN(n37115) );
  OAI222_X1 U33938 ( .A1(n30602), .A2(n39060), .B1(n30666), .B2(n39054), .C1(
        n30538), .C2(n39048), .ZN(n37122) );
  AOI221_X1 U33939 ( .B1(n39192), .B2(n29100), .C1(n39186), .C2(n29164), .A(
        n37114), .ZN(n37107) );
  OAI222_X1 U33940 ( .A1(n31488), .A2(n39180), .B1(n31552), .B2(n39174), .C1(
        n31424), .C2(n39168), .ZN(n37114) );
  AOI221_X1 U33941 ( .B1(n39072), .B2(n30473), .C1(n39066), .C2(n28000), .A(
        n37103), .ZN(n37096) );
  OAI222_X1 U33942 ( .A1(n30601), .A2(n39060), .B1(n30665), .B2(n39054), .C1(
        n30537), .C2(n39048), .ZN(n37103) );
  AOI221_X1 U33943 ( .B1(n39192), .B2(n29099), .C1(n39186), .C2(n29163), .A(
        n37095), .ZN(n37088) );
  OAI222_X1 U33944 ( .A1(n31487), .A2(n39180), .B1(n31551), .B2(n39174), .C1(
        n31423), .C2(n39168), .ZN(n37095) );
  AOI221_X1 U33945 ( .B1(n39072), .B2(n30472), .C1(n39066), .C2(n27999), .A(
        n37084), .ZN(n37077) );
  OAI222_X1 U33946 ( .A1(n30600), .A2(n39060), .B1(n30664), .B2(n39054), .C1(
        n30536), .C2(n39048), .ZN(n37084) );
  AOI221_X1 U33947 ( .B1(n39192), .B2(n29098), .C1(n39186), .C2(n29162), .A(
        n37076), .ZN(n37069) );
  OAI222_X1 U33948 ( .A1(n31486), .A2(n39180), .B1(n31550), .B2(n39174), .C1(
        n31422), .C2(n39168), .ZN(n37076) );
  AOI221_X1 U33949 ( .B1(n39072), .B2(n30471), .C1(n39066), .C2(n27998), .A(
        n37065), .ZN(n37058) );
  OAI222_X1 U33950 ( .A1(n30599), .A2(n39060), .B1(n30663), .B2(n39054), .C1(
        n30535), .C2(n39048), .ZN(n37065) );
  AOI221_X1 U33951 ( .B1(n39192), .B2(n29097), .C1(n39186), .C2(n29161), .A(
        n37057), .ZN(n37050) );
  OAI222_X1 U33952 ( .A1(n31485), .A2(n39180), .B1(n31549), .B2(n39174), .C1(
        n31421), .C2(n39168), .ZN(n37057) );
  AOI221_X1 U33953 ( .B1(n39072), .B2(n30470), .C1(n39066), .C2(n27997), .A(
        n37046), .ZN(n37039) );
  OAI222_X1 U33954 ( .A1(n30598), .A2(n39060), .B1(n30662), .B2(n39054), .C1(
        n30534), .C2(n39048), .ZN(n37046) );
  AOI221_X1 U33955 ( .B1(n39192), .B2(n29096), .C1(n39186), .C2(n29160), .A(
        n37038), .ZN(n37031) );
  OAI222_X1 U33956 ( .A1(n31484), .A2(n39180), .B1(n31548), .B2(n39174), .C1(
        n31420), .C2(n39168), .ZN(n37038) );
  AOI221_X1 U33957 ( .B1(n39076), .B2(n32515), .C1(n39070), .C2(n27953), .A(
        n36210), .ZN(n36203) );
  OAI222_X1 U33958 ( .A1(n30554), .A2(n39064), .B1(n30618), .B2(n39058), .C1(
        n30490), .C2(n39052), .ZN(n36210) );
  AOI221_X1 U33959 ( .B1(n39196), .B2(n29052), .C1(n39190), .C2(n29116), .A(
        n36202), .ZN(n36195) );
  OAI222_X1 U33960 ( .A1(n31440), .A2(n39184), .B1(n31504), .B2(n39178), .C1(
        n31376), .C2(n39172), .ZN(n36202) );
  AOI221_X1 U33961 ( .B1(n39076), .B2(n32514), .C1(n39070), .C2(n27952), .A(
        n36191), .ZN(n36184) );
  OAI222_X1 U33962 ( .A1(n30553), .A2(n39064), .B1(n30617), .B2(n39058), .C1(
        n30489), .C2(n39052), .ZN(n36191) );
  AOI221_X1 U33963 ( .B1(n39196), .B2(n29051), .C1(n39190), .C2(n29115), .A(
        n36183), .ZN(n36176) );
  OAI222_X1 U33964 ( .A1(n31439), .A2(n39184), .B1(n31503), .B2(n39178), .C1(
        n31375), .C2(n39172), .ZN(n36183) );
  AOI221_X1 U33965 ( .B1(n39076), .B2(n32513), .C1(n39070), .C2(n27951), .A(
        n36172), .ZN(n36165) );
  OAI222_X1 U33966 ( .A1(n30552), .A2(n39064), .B1(n30616), .B2(n39058), .C1(
        n30488), .C2(n39052), .ZN(n36172) );
  AOI221_X1 U33967 ( .B1(n39196), .B2(n29050), .C1(n39190), .C2(n29114), .A(
        n36164), .ZN(n36157) );
  OAI222_X1 U33968 ( .A1(n31438), .A2(n39184), .B1(n31502), .B2(n39178), .C1(
        n31374), .C2(n39172), .ZN(n36164) );
  AOI221_X1 U33969 ( .B1(n39076), .B2(n32512), .C1(n39070), .C2(n27950), .A(
        n36153), .ZN(n36146) );
  OAI222_X1 U33970 ( .A1(n30551), .A2(n39064), .B1(n30615), .B2(n39058), .C1(
        n30487), .C2(n39052), .ZN(n36153) );
  AOI221_X1 U33971 ( .B1(n39196), .B2(n29049), .C1(n39190), .C2(n29113), .A(
        n36145), .ZN(n36138) );
  OAI222_X1 U33972 ( .A1(n31437), .A2(n39184), .B1(n31501), .B2(n39178), .C1(
        n31373), .C2(n39172), .ZN(n36145) );
  AOI221_X1 U33973 ( .B1(n39076), .B2(n32511), .C1(n39070), .C2(n27949), .A(
        n36134), .ZN(n36127) );
  OAI222_X1 U33974 ( .A1(n30550), .A2(n39064), .B1(n30614), .B2(n39058), .C1(
        n30486), .C2(n39052), .ZN(n36134) );
  AOI221_X1 U33975 ( .B1(n39196), .B2(n29048), .C1(n39190), .C2(n29112), .A(
        n36126), .ZN(n36119) );
  OAI222_X1 U33976 ( .A1(n31436), .A2(n39184), .B1(n31500), .B2(n39178), .C1(
        n31372), .C2(n39172), .ZN(n36126) );
  AOI221_X1 U33977 ( .B1(n39076), .B2(n32510), .C1(n39070), .C2(n27948), .A(
        n36115), .ZN(n36108) );
  OAI222_X1 U33978 ( .A1(n30549), .A2(n39064), .B1(n30613), .B2(n39058), .C1(
        n30485), .C2(n39052), .ZN(n36115) );
  AOI221_X1 U33979 ( .B1(n39196), .B2(n29047), .C1(n39190), .C2(n29111), .A(
        n36107), .ZN(n36100) );
  OAI222_X1 U33980 ( .A1(n31435), .A2(n39184), .B1(n31499), .B2(n39178), .C1(
        n31371), .C2(n39172), .ZN(n36107) );
  AOI221_X1 U33981 ( .B1(n39579), .B2(n30480), .C1(n39573), .C2(n28007), .A(
        n33481), .ZN(n33457) );
  OAI222_X1 U33982 ( .A1(n30608), .A2(n39567), .B1(n30672), .B2(n39561), .C1(
        n30544), .C2(n39555), .ZN(n33481) );
  AOI221_X1 U33983 ( .B1(n39699), .B2(n29106), .C1(n39693), .C2(n29170), .A(
        n33453), .ZN(n33429) );
  OAI222_X1 U33984 ( .A1(n31494), .A2(n39687), .B1(n31558), .B2(n39681), .C1(
        n31430), .C2(n39675), .ZN(n33453) );
  AOI221_X1 U33985 ( .B1(n39327), .B2(n30480), .C1(n39321), .C2(n28007), .A(
        n34755), .ZN(n34731) );
  OAI222_X1 U33986 ( .A1(n30608), .A2(n39315), .B1(n30672), .B2(n39309), .C1(
        n30544), .C2(n39303), .ZN(n34755) );
  AOI221_X1 U33987 ( .B1(n39447), .B2(n29106), .C1(n39441), .C2(n29170), .A(
        n34727), .ZN(n34703) );
  OAI222_X1 U33988 ( .A1(n31494), .A2(n39435), .B1(n31558), .B2(n39429), .C1(
        n31430), .C2(n39423), .ZN(n34727) );
  AOI221_X1 U33989 ( .B1(n39579), .B2(n30479), .C1(n39573), .C2(n28006), .A(
        n33503), .ZN(n33496) );
  OAI222_X1 U33990 ( .A1(n30607), .A2(n39567), .B1(n30671), .B2(n39561), .C1(
        n30543), .C2(n39555), .ZN(n33503) );
  AOI221_X1 U33991 ( .B1(n39699), .B2(n29105), .C1(n39693), .C2(n29169), .A(
        n33495), .ZN(n33488) );
  OAI222_X1 U33992 ( .A1(n31493), .A2(n39687), .B1(n31557), .B2(n39681), .C1(
        n31429), .C2(n39675), .ZN(n33495) );
  AOI221_X1 U33993 ( .B1(n39327), .B2(n30479), .C1(n39321), .C2(n28006), .A(
        n34777), .ZN(n34770) );
  OAI222_X1 U33994 ( .A1(n30607), .A2(n39315), .B1(n30671), .B2(n39309), .C1(
        n30543), .C2(n39303), .ZN(n34777) );
  AOI221_X1 U33995 ( .B1(n39447), .B2(n29105), .C1(n39441), .C2(n29169), .A(
        n34769), .ZN(n34762) );
  OAI222_X1 U33996 ( .A1(n31493), .A2(n39435), .B1(n31557), .B2(n39429), .C1(
        n31429), .C2(n39423), .ZN(n34769) );
  AOI221_X1 U33997 ( .B1(n39579), .B2(n30478), .C1(n39573), .C2(n28005), .A(
        n33522), .ZN(n33515) );
  OAI222_X1 U33998 ( .A1(n30606), .A2(n39567), .B1(n30670), .B2(n39561), .C1(
        n30542), .C2(n39555), .ZN(n33522) );
  AOI221_X1 U33999 ( .B1(n39699), .B2(n29104), .C1(n39693), .C2(n29168), .A(
        n33514), .ZN(n33507) );
  OAI222_X1 U34000 ( .A1(n31492), .A2(n39687), .B1(n31556), .B2(n39681), .C1(
        n31428), .C2(n39675), .ZN(n33514) );
  AOI221_X1 U34001 ( .B1(n39327), .B2(n30478), .C1(n39321), .C2(n28005), .A(
        n34796), .ZN(n34789) );
  OAI222_X1 U34002 ( .A1(n30606), .A2(n39315), .B1(n30670), .B2(n39309), .C1(
        n30542), .C2(n39303), .ZN(n34796) );
  AOI221_X1 U34003 ( .B1(n39447), .B2(n29104), .C1(n39441), .C2(n29168), .A(
        n34788), .ZN(n34781) );
  OAI222_X1 U34004 ( .A1(n31492), .A2(n39435), .B1(n31556), .B2(n39429), .C1(
        n31428), .C2(n39423), .ZN(n34788) );
  AOI221_X1 U34005 ( .B1(n39579), .B2(n30477), .C1(n39573), .C2(n28004), .A(
        n33541), .ZN(n33534) );
  OAI222_X1 U34006 ( .A1(n30605), .A2(n39567), .B1(n30669), .B2(n39561), .C1(
        n30541), .C2(n39555), .ZN(n33541) );
  AOI221_X1 U34007 ( .B1(n39699), .B2(n29103), .C1(n39693), .C2(n29167), .A(
        n33533), .ZN(n33526) );
  OAI222_X1 U34008 ( .A1(n31491), .A2(n39687), .B1(n31555), .B2(n39681), .C1(
        n31427), .C2(n39675), .ZN(n33533) );
  AOI221_X1 U34009 ( .B1(n39327), .B2(n30477), .C1(n39321), .C2(n28004), .A(
        n34815), .ZN(n34808) );
  OAI222_X1 U34010 ( .A1(n30605), .A2(n39315), .B1(n30669), .B2(n39309), .C1(
        n30541), .C2(n39303), .ZN(n34815) );
  AOI221_X1 U34011 ( .B1(n39447), .B2(n29103), .C1(n39441), .C2(n29167), .A(
        n34807), .ZN(n34800) );
  OAI222_X1 U34012 ( .A1(n31491), .A2(n39435), .B1(n31555), .B2(n39429), .C1(
        n31427), .C2(n39423), .ZN(n34807) );
  AOI221_X1 U34013 ( .B1(n39578), .B2(n30476), .C1(n39572), .C2(n28003), .A(
        n33560), .ZN(n33553) );
  OAI222_X1 U34014 ( .A1(n30604), .A2(n39566), .B1(n30668), .B2(n39560), .C1(
        n30540), .C2(n39554), .ZN(n33560) );
  AOI221_X1 U34015 ( .B1(n39698), .B2(n29102), .C1(n39692), .C2(n29166), .A(
        n33552), .ZN(n33545) );
  OAI222_X1 U34016 ( .A1(n31490), .A2(n39686), .B1(n31554), .B2(n39680), .C1(
        n31426), .C2(n39674), .ZN(n33552) );
  AOI221_X1 U34017 ( .B1(n39326), .B2(n30476), .C1(n39320), .C2(n28003), .A(
        n34834), .ZN(n34827) );
  OAI222_X1 U34018 ( .A1(n30604), .A2(n39314), .B1(n30668), .B2(n39308), .C1(
        n30540), .C2(n39302), .ZN(n34834) );
  AOI221_X1 U34019 ( .B1(n39446), .B2(n29102), .C1(n39440), .C2(n29166), .A(
        n34826), .ZN(n34819) );
  OAI222_X1 U34020 ( .A1(n31490), .A2(n39434), .B1(n31554), .B2(n39428), .C1(
        n31426), .C2(n39422), .ZN(n34826) );
  AOI221_X1 U34021 ( .B1(n39578), .B2(n30475), .C1(n39572), .C2(n28002), .A(
        n33579), .ZN(n33572) );
  OAI222_X1 U34022 ( .A1(n30603), .A2(n39566), .B1(n30667), .B2(n39560), .C1(
        n30539), .C2(n39554), .ZN(n33579) );
  AOI221_X1 U34023 ( .B1(n39698), .B2(n29101), .C1(n39692), .C2(n29165), .A(
        n33571), .ZN(n33564) );
  OAI222_X1 U34024 ( .A1(n31489), .A2(n39686), .B1(n31553), .B2(n39680), .C1(
        n31425), .C2(n39674), .ZN(n33571) );
  AOI221_X1 U34025 ( .B1(n39326), .B2(n30475), .C1(n39320), .C2(n28002), .A(
        n34853), .ZN(n34846) );
  OAI222_X1 U34026 ( .A1(n30603), .A2(n39314), .B1(n30667), .B2(n39308), .C1(
        n30539), .C2(n39302), .ZN(n34853) );
  AOI221_X1 U34027 ( .B1(n39446), .B2(n29101), .C1(n39440), .C2(n29165), .A(
        n34845), .ZN(n34838) );
  OAI222_X1 U34028 ( .A1(n31489), .A2(n39434), .B1(n31553), .B2(n39428), .C1(
        n31425), .C2(n39422), .ZN(n34845) );
  AOI221_X1 U34029 ( .B1(n39578), .B2(n30474), .C1(n39572), .C2(n28001), .A(
        n33598), .ZN(n33591) );
  OAI222_X1 U34030 ( .A1(n30602), .A2(n39566), .B1(n30666), .B2(n39560), .C1(
        n30538), .C2(n39554), .ZN(n33598) );
  AOI221_X1 U34031 ( .B1(n39698), .B2(n29100), .C1(n39692), .C2(n29164), .A(
        n33590), .ZN(n33583) );
  OAI222_X1 U34032 ( .A1(n31488), .A2(n39686), .B1(n31552), .B2(n39680), .C1(
        n31424), .C2(n39674), .ZN(n33590) );
  AOI221_X1 U34033 ( .B1(n39326), .B2(n30474), .C1(n39320), .C2(n28001), .A(
        n34872), .ZN(n34865) );
  OAI222_X1 U34034 ( .A1(n30602), .A2(n39314), .B1(n30666), .B2(n39308), .C1(
        n30538), .C2(n39302), .ZN(n34872) );
  AOI221_X1 U34035 ( .B1(n39446), .B2(n29100), .C1(n39440), .C2(n29164), .A(
        n34864), .ZN(n34857) );
  OAI222_X1 U34036 ( .A1(n31488), .A2(n39434), .B1(n31552), .B2(n39428), .C1(
        n31424), .C2(n39422), .ZN(n34864) );
  AOI221_X1 U34037 ( .B1(n39578), .B2(n30473), .C1(n39572), .C2(n28000), .A(
        n33617), .ZN(n33610) );
  OAI222_X1 U34038 ( .A1(n30601), .A2(n39566), .B1(n30665), .B2(n39560), .C1(
        n30537), .C2(n39554), .ZN(n33617) );
  AOI221_X1 U34039 ( .B1(n39698), .B2(n29099), .C1(n39692), .C2(n29163), .A(
        n33609), .ZN(n33602) );
  OAI222_X1 U34040 ( .A1(n31487), .A2(n39686), .B1(n31551), .B2(n39680), .C1(
        n31423), .C2(n39674), .ZN(n33609) );
  AOI221_X1 U34041 ( .B1(n39326), .B2(n30473), .C1(n39320), .C2(n28000), .A(
        n34891), .ZN(n34884) );
  OAI222_X1 U34042 ( .A1(n30601), .A2(n39314), .B1(n30665), .B2(n39308), .C1(
        n30537), .C2(n39302), .ZN(n34891) );
  AOI221_X1 U34043 ( .B1(n39446), .B2(n29099), .C1(n39440), .C2(n29163), .A(
        n34883), .ZN(n34876) );
  OAI222_X1 U34044 ( .A1(n31487), .A2(n39434), .B1(n31551), .B2(n39428), .C1(
        n31423), .C2(n39422), .ZN(n34883) );
  AOI221_X1 U34045 ( .B1(n39578), .B2(n30472), .C1(n39572), .C2(n27999), .A(
        n33636), .ZN(n33629) );
  OAI222_X1 U34046 ( .A1(n30600), .A2(n39566), .B1(n30664), .B2(n39560), .C1(
        n30536), .C2(n39554), .ZN(n33636) );
  AOI221_X1 U34047 ( .B1(n39698), .B2(n29098), .C1(n39692), .C2(n29162), .A(
        n33628), .ZN(n33621) );
  OAI222_X1 U34048 ( .A1(n31486), .A2(n39686), .B1(n31550), .B2(n39680), .C1(
        n31422), .C2(n39674), .ZN(n33628) );
  AOI221_X1 U34049 ( .B1(n39326), .B2(n30472), .C1(n39320), .C2(n27999), .A(
        n34910), .ZN(n34903) );
  OAI222_X1 U34050 ( .A1(n30600), .A2(n39314), .B1(n30664), .B2(n39308), .C1(
        n30536), .C2(n39302), .ZN(n34910) );
  AOI221_X1 U34051 ( .B1(n39446), .B2(n29098), .C1(n39440), .C2(n29162), .A(
        n34902), .ZN(n34895) );
  OAI222_X1 U34052 ( .A1(n31486), .A2(n39434), .B1(n31550), .B2(n39428), .C1(
        n31422), .C2(n39422), .ZN(n34902) );
  AOI221_X1 U34053 ( .B1(n39578), .B2(n30471), .C1(n39572), .C2(n27998), .A(
        n33655), .ZN(n33648) );
  OAI222_X1 U34054 ( .A1(n30599), .A2(n39566), .B1(n30663), .B2(n39560), .C1(
        n30535), .C2(n39554), .ZN(n33655) );
  AOI221_X1 U34055 ( .B1(n39698), .B2(n29097), .C1(n39692), .C2(n29161), .A(
        n33647), .ZN(n33640) );
  OAI222_X1 U34056 ( .A1(n31485), .A2(n39686), .B1(n31549), .B2(n39680), .C1(
        n31421), .C2(n39674), .ZN(n33647) );
  AOI221_X1 U34057 ( .B1(n39326), .B2(n30471), .C1(n39320), .C2(n27998), .A(
        n34929), .ZN(n34922) );
  OAI222_X1 U34058 ( .A1(n30599), .A2(n39314), .B1(n30663), .B2(n39308), .C1(
        n30535), .C2(n39302), .ZN(n34929) );
  AOI221_X1 U34059 ( .B1(n39446), .B2(n29097), .C1(n39440), .C2(n29161), .A(
        n34921), .ZN(n34914) );
  OAI222_X1 U34060 ( .A1(n31485), .A2(n39434), .B1(n31549), .B2(n39428), .C1(
        n31421), .C2(n39422), .ZN(n34921) );
  AOI221_X1 U34061 ( .B1(n39578), .B2(n30470), .C1(n39572), .C2(n27997), .A(
        n33674), .ZN(n33667) );
  OAI222_X1 U34062 ( .A1(n30598), .A2(n39566), .B1(n30662), .B2(n39560), .C1(
        n30534), .C2(n39554), .ZN(n33674) );
  AOI221_X1 U34063 ( .B1(n39698), .B2(n29096), .C1(n39692), .C2(n29160), .A(
        n33666), .ZN(n33659) );
  OAI222_X1 U34064 ( .A1(n31484), .A2(n39686), .B1(n31548), .B2(n39680), .C1(
        n31420), .C2(n39674), .ZN(n33666) );
  AOI221_X1 U34065 ( .B1(n39326), .B2(n30470), .C1(n39320), .C2(n27997), .A(
        n34948), .ZN(n34941) );
  OAI222_X1 U34066 ( .A1(n30598), .A2(n39314), .B1(n30662), .B2(n39308), .C1(
        n30534), .C2(n39302), .ZN(n34948) );
  AOI221_X1 U34067 ( .B1(n39446), .B2(n29096), .C1(n39440), .C2(n29160), .A(
        n34940), .ZN(n34933) );
  OAI222_X1 U34068 ( .A1(n31484), .A2(n39434), .B1(n31548), .B2(n39428), .C1(
        n31420), .C2(n39422), .ZN(n34940) );
  AOI221_X1 U34069 ( .B1(n39578), .B2(n30469), .C1(n39572), .C2(n27996), .A(
        n33693), .ZN(n33686) );
  OAI222_X1 U34070 ( .A1(n30597), .A2(n39566), .B1(n30661), .B2(n39560), .C1(
        n30533), .C2(n39554), .ZN(n33693) );
  AOI221_X1 U34071 ( .B1(n39698), .B2(n29095), .C1(n39692), .C2(n29159), .A(
        n33685), .ZN(n33678) );
  OAI222_X1 U34072 ( .A1(n31483), .A2(n39686), .B1(n31547), .B2(n39680), .C1(
        n31419), .C2(n39674), .ZN(n33685) );
  AOI221_X1 U34073 ( .B1(n39326), .B2(n30469), .C1(n39320), .C2(n27996), .A(
        n34967), .ZN(n34960) );
  OAI222_X1 U34074 ( .A1(n30597), .A2(n39314), .B1(n30661), .B2(n39308), .C1(
        n30533), .C2(n39302), .ZN(n34967) );
  AOI221_X1 U34075 ( .B1(n39446), .B2(n29095), .C1(n39440), .C2(n29159), .A(
        n34959), .ZN(n34952) );
  OAI222_X1 U34076 ( .A1(n31483), .A2(n39434), .B1(n31547), .B2(n39428), .C1(
        n31419), .C2(n39422), .ZN(n34959) );
  AOI221_X1 U34077 ( .B1(n39578), .B2(n30468), .C1(n39572), .C2(n27995), .A(
        n33712), .ZN(n33705) );
  OAI222_X1 U34078 ( .A1(n30596), .A2(n39566), .B1(n30660), .B2(n39560), .C1(
        n30532), .C2(n39554), .ZN(n33712) );
  AOI221_X1 U34079 ( .B1(n39698), .B2(n29094), .C1(n39692), .C2(n29158), .A(
        n33704), .ZN(n33697) );
  OAI222_X1 U34080 ( .A1(n31482), .A2(n39686), .B1(n31546), .B2(n39680), .C1(
        n31418), .C2(n39674), .ZN(n33704) );
  AOI221_X1 U34081 ( .B1(n39326), .B2(n30468), .C1(n39320), .C2(n27995), .A(
        n34986), .ZN(n34979) );
  OAI222_X1 U34082 ( .A1(n30596), .A2(n39314), .B1(n30660), .B2(n39308), .C1(
        n30532), .C2(n39302), .ZN(n34986) );
  AOI221_X1 U34083 ( .B1(n39446), .B2(n29094), .C1(n39440), .C2(n29158), .A(
        n34978), .ZN(n34971) );
  OAI222_X1 U34084 ( .A1(n31482), .A2(n39434), .B1(n31546), .B2(n39428), .C1(
        n31418), .C2(n39422), .ZN(n34978) );
  AOI221_X1 U34085 ( .B1(n39578), .B2(n30467), .C1(n39572), .C2(n27994), .A(
        n33731), .ZN(n33724) );
  OAI222_X1 U34086 ( .A1(n30595), .A2(n39566), .B1(n30659), .B2(n39560), .C1(
        n30531), .C2(n39554), .ZN(n33731) );
  AOI221_X1 U34087 ( .B1(n39698), .B2(n29093), .C1(n39692), .C2(n29157), .A(
        n33723), .ZN(n33716) );
  OAI222_X1 U34088 ( .A1(n31481), .A2(n39686), .B1(n31545), .B2(n39680), .C1(
        n31417), .C2(n39674), .ZN(n33723) );
  AOI221_X1 U34089 ( .B1(n39326), .B2(n30467), .C1(n39320), .C2(n27994), .A(
        n35005), .ZN(n34998) );
  OAI222_X1 U34090 ( .A1(n30595), .A2(n39314), .B1(n30659), .B2(n39308), .C1(
        n30531), .C2(n39302), .ZN(n35005) );
  AOI221_X1 U34091 ( .B1(n39446), .B2(n29093), .C1(n39440), .C2(n29157), .A(
        n34997), .ZN(n34990) );
  OAI222_X1 U34092 ( .A1(n31481), .A2(n39434), .B1(n31545), .B2(n39428), .C1(
        n31417), .C2(n39422), .ZN(n34997) );
  AOI221_X1 U34093 ( .B1(n39578), .B2(n30466), .C1(n39572), .C2(n27993), .A(
        n33750), .ZN(n33743) );
  OAI222_X1 U34094 ( .A1(n30594), .A2(n39566), .B1(n30658), .B2(n39560), .C1(
        n30530), .C2(n39554), .ZN(n33750) );
  AOI221_X1 U34095 ( .B1(n39698), .B2(n29092), .C1(n39692), .C2(n29156), .A(
        n33742), .ZN(n33735) );
  OAI222_X1 U34096 ( .A1(n31480), .A2(n39686), .B1(n31544), .B2(n39680), .C1(
        n31416), .C2(n39674), .ZN(n33742) );
  AOI221_X1 U34097 ( .B1(n39326), .B2(n30466), .C1(n39320), .C2(n27993), .A(
        n35024), .ZN(n35017) );
  OAI222_X1 U34098 ( .A1(n30594), .A2(n39314), .B1(n30658), .B2(n39308), .C1(
        n30530), .C2(n39302), .ZN(n35024) );
  AOI221_X1 U34099 ( .B1(n39446), .B2(n29092), .C1(n39440), .C2(n29156), .A(
        n35016), .ZN(n35009) );
  OAI222_X1 U34100 ( .A1(n31480), .A2(n39434), .B1(n31544), .B2(n39428), .C1(
        n31416), .C2(n39422), .ZN(n35016) );
  AOI221_X1 U34101 ( .B1(n39578), .B2(n30465), .C1(n39572), .C2(n27992), .A(
        n33769), .ZN(n33762) );
  OAI222_X1 U34102 ( .A1(n30593), .A2(n39566), .B1(n30657), .B2(n39560), .C1(
        n30529), .C2(n39554), .ZN(n33769) );
  AOI221_X1 U34103 ( .B1(n39698), .B2(n29091), .C1(n39692), .C2(n29155), .A(
        n33761), .ZN(n33754) );
  OAI222_X1 U34104 ( .A1(n31479), .A2(n39686), .B1(n31543), .B2(n39680), .C1(
        n31415), .C2(n39674), .ZN(n33761) );
  AOI221_X1 U34105 ( .B1(n39326), .B2(n30465), .C1(n39320), .C2(n27992), .A(
        n35043), .ZN(n35036) );
  OAI222_X1 U34106 ( .A1(n30593), .A2(n39314), .B1(n30657), .B2(n39308), .C1(
        n30529), .C2(n39302), .ZN(n35043) );
  AOI221_X1 U34107 ( .B1(n39446), .B2(n29091), .C1(n39440), .C2(n29155), .A(
        n35035), .ZN(n35028) );
  OAI222_X1 U34108 ( .A1(n31479), .A2(n39434), .B1(n31543), .B2(n39428), .C1(
        n31415), .C2(n39422), .ZN(n35035) );
  AOI221_X1 U34109 ( .B1(n39577), .B2(n30464), .C1(n39571), .C2(n27991), .A(
        n33788), .ZN(n33781) );
  OAI222_X1 U34110 ( .A1(n30592), .A2(n39565), .B1(n30656), .B2(n39559), .C1(
        n30528), .C2(n39553), .ZN(n33788) );
  AOI221_X1 U34111 ( .B1(n39697), .B2(n29090), .C1(n39691), .C2(n29154), .A(
        n33780), .ZN(n33773) );
  OAI222_X1 U34112 ( .A1(n31478), .A2(n39685), .B1(n31542), .B2(n39679), .C1(
        n31414), .C2(n39673), .ZN(n33780) );
  AOI221_X1 U34113 ( .B1(n39325), .B2(n30464), .C1(n39319), .C2(n27991), .A(
        n35062), .ZN(n35055) );
  OAI222_X1 U34114 ( .A1(n30592), .A2(n39313), .B1(n30656), .B2(n39307), .C1(
        n30528), .C2(n39301), .ZN(n35062) );
  AOI221_X1 U34115 ( .B1(n39445), .B2(n29090), .C1(n39439), .C2(n29154), .A(
        n35054), .ZN(n35047) );
  OAI222_X1 U34116 ( .A1(n31478), .A2(n39433), .B1(n31542), .B2(n39427), .C1(
        n31414), .C2(n39421), .ZN(n35054) );
  AOI221_X1 U34117 ( .B1(n39577), .B2(n30463), .C1(n39571), .C2(n27990), .A(
        n33807), .ZN(n33800) );
  OAI222_X1 U34118 ( .A1(n30591), .A2(n39565), .B1(n30655), .B2(n39559), .C1(
        n30527), .C2(n39553), .ZN(n33807) );
  AOI221_X1 U34119 ( .B1(n39697), .B2(n29089), .C1(n39691), .C2(n29153), .A(
        n33799), .ZN(n33792) );
  OAI222_X1 U34120 ( .A1(n31477), .A2(n39685), .B1(n31541), .B2(n39679), .C1(
        n31413), .C2(n39673), .ZN(n33799) );
  AOI221_X1 U34121 ( .B1(n39325), .B2(n30463), .C1(n39319), .C2(n27990), .A(
        n35081), .ZN(n35074) );
  OAI222_X1 U34122 ( .A1(n30591), .A2(n39313), .B1(n30655), .B2(n39307), .C1(
        n30527), .C2(n39301), .ZN(n35081) );
  AOI221_X1 U34123 ( .B1(n39445), .B2(n29089), .C1(n39439), .C2(n29153), .A(
        n35073), .ZN(n35066) );
  OAI222_X1 U34124 ( .A1(n31477), .A2(n39433), .B1(n31541), .B2(n39427), .C1(
        n31413), .C2(n39421), .ZN(n35073) );
  AOI221_X1 U34125 ( .B1(n39577), .B2(n30462), .C1(n39571), .C2(n27989), .A(
        n33826), .ZN(n33819) );
  OAI222_X1 U34126 ( .A1(n30590), .A2(n39565), .B1(n30654), .B2(n39559), .C1(
        n30526), .C2(n39553), .ZN(n33826) );
  AOI221_X1 U34127 ( .B1(n39697), .B2(n29088), .C1(n39691), .C2(n29152), .A(
        n33818), .ZN(n33811) );
  OAI222_X1 U34128 ( .A1(n31476), .A2(n39685), .B1(n31540), .B2(n39679), .C1(
        n31412), .C2(n39673), .ZN(n33818) );
  AOI221_X1 U34129 ( .B1(n39325), .B2(n30462), .C1(n39319), .C2(n27989), .A(
        n35100), .ZN(n35093) );
  OAI222_X1 U34130 ( .A1(n30590), .A2(n39313), .B1(n30654), .B2(n39307), .C1(
        n30526), .C2(n39301), .ZN(n35100) );
  AOI221_X1 U34131 ( .B1(n39445), .B2(n29088), .C1(n39439), .C2(n29152), .A(
        n35092), .ZN(n35085) );
  OAI222_X1 U34132 ( .A1(n31476), .A2(n39433), .B1(n31540), .B2(n39427), .C1(
        n31412), .C2(n39421), .ZN(n35092) );
  AOI221_X1 U34133 ( .B1(n39577), .B2(n30461), .C1(n39571), .C2(n27988), .A(
        n33845), .ZN(n33838) );
  OAI222_X1 U34134 ( .A1(n30589), .A2(n39565), .B1(n30653), .B2(n39559), .C1(
        n30525), .C2(n39553), .ZN(n33845) );
  AOI221_X1 U34135 ( .B1(n39697), .B2(n29087), .C1(n39691), .C2(n29151), .A(
        n33837), .ZN(n33830) );
  OAI222_X1 U34136 ( .A1(n31475), .A2(n39685), .B1(n31539), .B2(n39679), .C1(
        n31411), .C2(n39673), .ZN(n33837) );
  AOI221_X1 U34137 ( .B1(n39325), .B2(n30461), .C1(n39319), .C2(n27988), .A(
        n35119), .ZN(n35112) );
  OAI222_X1 U34138 ( .A1(n30589), .A2(n39313), .B1(n30653), .B2(n39307), .C1(
        n30525), .C2(n39301), .ZN(n35119) );
  AOI221_X1 U34139 ( .B1(n39445), .B2(n29087), .C1(n39439), .C2(n29151), .A(
        n35111), .ZN(n35104) );
  OAI222_X1 U34140 ( .A1(n31475), .A2(n39433), .B1(n31539), .B2(n39427), .C1(
        n31411), .C2(n39421), .ZN(n35111) );
  AOI221_X1 U34141 ( .B1(n39577), .B2(n30460), .C1(n39571), .C2(n27987), .A(
        n33864), .ZN(n33857) );
  OAI222_X1 U34142 ( .A1(n30588), .A2(n39565), .B1(n30652), .B2(n39559), .C1(
        n30524), .C2(n39553), .ZN(n33864) );
  AOI221_X1 U34143 ( .B1(n39697), .B2(n29086), .C1(n39691), .C2(n29150), .A(
        n33856), .ZN(n33849) );
  OAI222_X1 U34144 ( .A1(n31474), .A2(n39685), .B1(n31538), .B2(n39679), .C1(
        n31410), .C2(n39673), .ZN(n33856) );
  AOI221_X1 U34145 ( .B1(n39325), .B2(n30460), .C1(n39319), .C2(n27987), .A(
        n35138), .ZN(n35131) );
  OAI222_X1 U34146 ( .A1(n30588), .A2(n39313), .B1(n30652), .B2(n39307), .C1(
        n30524), .C2(n39301), .ZN(n35138) );
  AOI221_X1 U34147 ( .B1(n39445), .B2(n29086), .C1(n39439), .C2(n29150), .A(
        n35130), .ZN(n35123) );
  OAI222_X1 U34148 ( .A1(n31474), .A2(n39433), .B1(n31538), .B2(n39427), .C1(
        n31410), .C2(n39421), .ZN(n35130) );
  AOI221_X1 U34149 ( .B1(n39577), .B2(n30459), .C1(n39571), .C2(n27986), .A(
        n33883), .ZN(n33876) );
  OAI222_X1 U34150 ( .A1(n30587), .A2(n39565), .B1(n30651), .B2(n39559), .C1(
        n30523), .C2(n39553), .ZN(n33883) );
  AOI221_X1 U34151 ( .B1(n39697), .B2(n29085), .C1(n39691), .C2(n29149), .A(
        n33875), .ZN(n33868) );
  OAI222_X1 U34152 ( .A1(n31473), .A2(n39685), .B1(n31537), .B2(n39679), .C1(
        n31409), .C2(n39673), .ZN(n33875) );
  AOI221_X1 U34153 ( .B1(n39325), .B2(n30459), .C1(n39319), .C2(n27986), .A(
        n35157), .ZN(n35150) );
  OAI222_X1 U34154 ( .A1(n30587), .A2(n39313), .B1(n30651), .B2(n39307), .C1(
        n30523), .C2(n39301), .ZN(n35157) );
  AOI221_X1 U34155 ( .B1(n39445), .B2(n29085), .C1(n39439), .C2(n29149), .A(
        n35149), .ZN(n35142) );
  OAI222_X1 U34156 ( .A1(n31473), .A2(n39433), .B1(n31537), .B2(n39427), .C1(
        n31409), .C2(n39421), .ZN(n35149) );
  AOI221_X1 U34157 ( .B1(n39577), .B2(n30458), .C1(n39571), .C2(n27985), .A(
        n33902), .ZN(n33895) );
  OAI222_X1 U34158 ( .A1(n30586), .A2(n39565), .B1(n30650), .B2(n39559), .C1(
        n30522), .C2(n39553), .ZN(n33902) );
  AOI221_X1 U34159 ( .B1(n39697), .B2(n29084), .C1(n39691), .C2(n29148), .A(
        n33894), .ZN(n33887) );
  OAI222_X1 U34160 ( .A1(n31472), .A2(n39685), .B1(n31536), .B2(n39679), .C1(
        n31408), .C2(n39673), .ZN(n33894) );
  AOI221_X1 U34161 ( .B1(n39325), .B2(n30458), .C1(n39319), .C2(n27985), .A(
        n35176), .ZN(n35169) );
  OAI222_X1 U34162 ( .A1(n30586), .A2(n39313), .B1(n30650), .B2(n39307), .C1(
        n30522), .C2(n39301), .ZN(n35176) );
  AOI221_X1 U34163 ( .B1(n39445), .B2(n29084), .C1(n39439), .C2(n29148), .A(
        n35168), .ZN(n35161) );
  OAI222_X1 U34164 ( .A1(n31472), .A2(n39433), .B1(n31536), .B2(n39427), .C1(
        n31408), .C2(n39421), .ZN(n35168) );
  AOI221_X1 U34165 ( .B1(n39577), .B2(n32546), .C1(n39571), .C2(n27984), .A(
        n33921), .ZN(n33914) );
  OAI222_X1 U34166 ( .A1(n30585), .A2(n39565), .B1(n30649), .B2(n39559), .C1(
        n30521), .C2(n39553), .ZN(n33921) );
  AOI221_X1 U34167 ( .B1(n39697), .B2(n29083), .C1(n39691), .C2(n29147), .A(
        n33913), .ZN(n33906) );
  OAI222_X1 U34168 ( .A1(n31471), .A2(n39685), .B1(n31535), .B2(n39679), .C1(
        n31407), .C2(n39673), .ZN(n33913) );
  AOI221_X1 U34169 ( .B1(n39325), .B2(n32546), .C1(n39319), .C2(n27984), .A(
        n35195), .ZN(n35188) );
  OAI222_X1 U34170 ( .A1(n30585), .A2(n39313), .B1(n30649), .B2(n39307), .C1(
        n30521), .C2(n39301), .ZN(n35195) );
  AOI221_X1 U34171 ( .B1(n39445), .B2(n29083), .C1(n39439), .C2(n29147), .A(
        n35187), .ZN(n35180) );
  OAI222_X1 U34172 ( .A1(n31471), .A2(n39433), .B1(n31535), .B2(n39427), .C1(
        n31407), .C2(n39421), .ZN(n35187) );
  AOI221_X1 U34173 ( .B1(n39577), .B2(n32545), .C1(n39571), .C2(n27983), .A(
        n33940), .ZN(n33933) );
  OAI222_X1 U34174 ( .A1(n30584), .A2(n39565), .B1(n30648), .B2(n39559), .C1(
        n30520), .C2(n39553), .ZN(n33940) );
  AOI221_X1 U34175 ( .B1(n39697), .B2(n29082), .C1(n39691), .C2(n29146), .A(
        n33932), .ZN(n33925) );
  OAI222_X1 U34176 ( .A1(n31470), .A2(n39685), .B1(n31534), .B2(n39679), .C1(
        n31406), .C2(n39673), .ZN(n33932) );
  AOI221_X1 U34177 ( .B1(n39325), .B2(n32545), .C1(n39319), .C2(n27983), .A(
        n35214), .ZN(n35207) );
  OAI222_X1 U34178 ( .A1(n30584), .A2(n39313), .B1(n30648), .B2(n39307), .C1(
        n30520), .C2(n39301), .ZN(n35214) );
  AOI221_X1 U34179 ( .B1(n39445), .B2(n29082), .C1(n39439), .C2(n29146), .A(
        n35206), .ZN(n35199) );
  OAI222_X1 U34180 ( .A1(n31470), .A2(n39433), .B1(n31534), .B2(n39427), .C1(
        n31406), .C2(n39421), .ZN(n35206) );
  AOI221_X1 U34181 ( .B1(n39577), .B2(n32544), .C1(n39571), .C2(n27982), .A(
        n33959), .ZN(n33952) );
  OAI222_X1 U34182 ( .A1(n30583), .A2(n39565), .B1(n30647), .B2(n39559), .C1(
        n30519), .C2(n39553), .ZN(n33959) );
  AOI221_X1 U34183 ( .B1(n39697), .B2(n29081), .C1(n39691), .C2(n29145), .A(
        n33951), .ZN(n33944) );
  OAI222_X1 U34184 ( .A1(n31469), .A2(n39685), .B1(n31533), .B2(n39679), .C1(
        n31405), .C2(n39673), .ZN(n33951) );
  AOI221_X1 U34185 ( .B1(n39325), .B2(n32544), .C1(n39319), .C2(n27982), .A(
        n35233), .ZN(n35226) );
  OAI222_X1 U34186 ( .A1(n30583), .A2(n39313), .B1(n30647), .B2(n39307), .C1(
        n30519), .C2(n39301), .ZN(n35233) );
  AOI221_X1 U34187 ( .B1(n39445), .B2(n29081), .C1(n39439), .C2(n29145), .A(
        n35225), .ZN(n35218) );
  OAI222_X1 U34188 ( .A1(n31469), .A2(n39433), .B1(n31533), .B2(n39427), .C1(
        n31405), .C2(n39421), .ZN(n35225) );
  AOI221_X1 U34189 ( .B1(n39577), .B2(n32543), .C1(n39571), .C2(n27981), .A(
        n33978), .ZN(n33971) );
  OAI222_X1 U34190 ( .A1(n30582), .A2(n39565), .B1(n30646), .B2(n39559), .C1(
        n30518), .C2(n39553), .ZN(n33978) );
  AOI221_X1 U34191 ( .B1(n39697), .B2(n29080), .C1(n39691), .C2(n29144), .A(
        n33970), .ZN(n33963) );
  OAI222_X1 U34192 ( .A1(n31468), .A2(n39685), .B1(n31532), .B2(n39679), .C1(
        n31404), .C2(n39673), .ZN(n33970) );
  AOI221_X1 U34193 ( .B1(n39325), .B2(n32543), .C1(n39319), .C2(n27981), .A(
        n35252), .ZN(n35245) );
  OAI222_X1 U34194 ( .A1(n30582), .A2(n39313), .B1(n30646), .B2(n39307), .C1(
        n30518), .C2(n39301), .ZN(n35252) );
  AOI221_X1 U34195 ( .B1(n39445), .B2(n29080), .C1(n39439), .C2(n29144), .A(
        n35244), .ZN(n35237) );
  OAI222_X1 U34196 ( .A1(n31468), .A2(n39433), .B1(n31532), .B2(n39427), .C1(
        n31404), .C2(n39421), .ZN(n35244) );
  AOI221_X1 U34197 ( .B1(n39577), .B2(n32542), .C1(n39571), .C2(n27980), .A(
        n33997), .ZN(n33990) );
  OAI222_X1 U34198 ( .A1(n30581), .A2(n39565), .B1(n30645), .B2(n39559), .C1(
        n30517), .C2(n39553), .ZN(n33997) );
  AOI221_X1 U34199 ( .B1(n39697), .B2(n29079), .C1(n39691), .C2(n29143), .A(
        n33989), .ZN(n33982) );
  OAI222_X1 U34200 ( .A1(n31467), .A2(n39685), .B1(n31531), .B2(n39679), .C1(
        n31403), .C2(n39673), .ZN(n33989) );
  AOI221_X1 U34201 ( .B1(n39325), .B2(n32542), .C1(n39319), .C2(n27980), .A(
        n35271), .ZN(n35264) );
  OAI222_X1 U34202 ( .A1(n30581), .A2(n39313), .B1(n30645), .B2(n39307), .C1(
        n30517), .C2(n39301), .ZN(n35271) );
  AOI221_X1 U34203 ( .B1(n39445), .B2(n29079), .C1(n39439), .C2(n29143), .A(
        n35263), .ZN(n35256) );
  OAI222_X1 U34204 ( .A1(n31467), .A2(n39433), .B1(n31531), .B2(n39427), .C1(
        n31403), .C2(n39421), .ZN(n35263) );
  AOI221_X1 U34205 ( .B1(n39576), .B2(n32541), .C1(n39570), .C2(n27979), .A(
        n34016), .ZN(n34009) );
  OAI222_X1 U34206 ( .A1(n30580), .A2(n39564), .B1(n30644), .B2(n39558), .C1(
        n30516), .C2(n39552), .ZN(n34016) );
  AOI221_X1 U34207 ( .B1(n39696), .B2(n29078), .C1(n39690), .C2(n29142), .A(
        n34008), .ZN(n34001) );
  OAI222_X1 U34208 ( .A1(n31466), .A2(n39684), .B1(n31530), .B2(n39678), .C1(
        n31402), .C2(n39672), .ZN(n34008) );
  AOI221_X1 U34209 ( .B1(n39324), .B2(n32541), .C1(n39318), .C2(n27979), .A(
        n35290), .ZN(n35283) );
  OAI222_X1 U34210 ( .A1(n30580), .A2(n39312), .B1(n30644), .B2(n39306), .C1(
        n30516), .C2(n39300), .ZN(n35290) );
  AOI221_X1 U34211 ( .B1(n39444), .B2(n29078), .C1(n39438), .C2(n29142), .A(
        n35282), .ZN(n35275) );
  OAI222_X1 U34212 ( .A1(n31466), .A2(n39432), .B1(n31530), .B2(n39426), .C1(
        n31402), .C2(n39420), .ZN(n35282) );
  AOI221_X1 U34213 ( .B1(n39576), .B2(n32540), .C1(n39570), .C2(n27978), .A(
        n34035), .ZN(n34028) );
  OAI222_X1 U34214 ( .A1(n30579), .A2(n39564), .B1(n30643), .B2(n39558), .C1(
        n30515), .C2(n39552), .ZN(n34035) );
  AOI221_X1 U34215 ( .B1(n39696), .B2(n29077), .C1(n39690), .C2(n29141), .A(
        n34027), .ZN(n34020) );
  OAI222_X1 U34216 ( .A1(n31465), .A2(n39684), .B1(n31529), .B2(n39678), .C1(
        n31401), .C2(n39672), .ZN(n34027) );
  AOI221_X1 U34217 ( .B1(n39324), .B2(n32540), .C1(n39318), .C2(n27978), .A(
        n35309), .ZN(n35302) );
  OAI222_X1 U34218 ( .A1(n30579), .A2(n39312), .B1(n30643), .B2(n39306), .C1(
        n30515), .C2(n39300), .ZN(n35309) );
  AOI221_X1 U34219 ( .B1(n39444), .B2(n29077), .C1(n39438), .C2(n29141), .A(
        n35301), .ZN(n35294) );
  OAI222_X1 U34220 ( .A1(n31465), .A2(n39432), .B1(n31529), .B2(n39426), .C1(
        n31401), .C2(n39420), .ZN(n35301) );
  AOI221_X1 U34221 ( .B1(n39576), .B2(n32539), .C1(n39570), .C2(n27977), .A(
        n34054), .ZN(n34047) );
  OAI222_X1 U34222 ( .A1(n30578), .A2(n39564), .B1(n30642), .B2(n39558), .C1(
        n30514), .C2(n39552), .ZN(n34054) );
  AOI221_X1 U34223 ( .B1(n39696), .B2(n29076), .C1(n39690), .C2(n29140), .A(
        n34046), .ZN(n34039) );
  OAI222_X1 U34224 ( .A1(n31464), .A2(n39684), .B1(n31528), .B2(n39678), .C1(
        n31400), .C2(n39672), .ZN(n34046) );
  AOI221_X1 U34225 ( .B1(n39324), .B2(n32539), .C1(n39318), .C2(n27977), .A(
        n35328), .ZN(n35321) );
  OAI222_X1 U34226 ( .A1(n30578), .A2(n39312), .B1(n30642), .B2(n39306), .C1(
        n30514), .C2(n39300), .ZN(n35328) );
  AOI221_X1 U34227 ( .B1(n39444), .B2(n29076), .C1(n39438), .C2(n29140), .A(
        n35320), .ZN(n35313) );
  OAI222_X1 U34228 ( .A1(n31464), .A2(n39432), .B1(n31528), .B2(n39426), .C1(
        n31400), .C2(n39420), .ZN(n35320) );
  AOI221_X1 U34229 ( .B1(n39576), .B2(n32538), .C1(n39570), .C2(n27976), .A(
        n34073), .ZN(n34066) );
  OAI222_X1 U34230 ( .A1(n30577), .A2(n39564), .B1(n30641), .B2(n39558), .C1(
        n30513), .C2(n39552), .ZN(n34073) );
  AOI221_X1 U34231 ( .B1(n39696), .B2(n29075), .C1(n39690), .C2(n29139), .A(
        n34065), .ZN(n34058) );
  OAI222_X1 U34232 ( .A1(n31463), .A2(n39684), .B1(n31527), .B2(n39678), .C1(
        n31399), .C2(n39672), .ZN(n34065) );
  AOI221_X1 U34233 ( .B1(n39324), .B2(n32538), .C1(n39318), .C2(n27976), .A(
        n35347), .ZN(n35340) );
  OAI222_X1 U34234 ( .A1(n30577), .A2(n39312), .B1(n30641), .B2(n39306), .C1(
        n30513), .C2(n39300), .ZN(n35347) );
  AOI221_X1 U34235 ( .B1(n39444), .B2(n29075), .C1(n39438), .C2(n29139), .A(
        n35339), .ZN(n35332) );
  OAI222_X1 U34236 ( .A1(n31463), .A2(n39432), .B1(n31527), .B2(n39426), .C1(
        n31399), .C2(n39420), .ZN(n35339) );
  AOI221_X1 U34237 ( .B1(n39576), .B2(n32537), .C1(n39570), .C2(n27975), .A(
        n34092), .ZN(n34085) );
  OAI222_X1 U34238 ( .A1(n30576), .A2(n39564), .B1(n30640), .B2(n39558), .C1(
        n30512), .C2(n39552), .ZN(n34092) );
  AOI221_X1 U34239 ( .B1(n39696), .B2(n29074), .C1(n39690), .C2(n29138), .A(
        n34084), .ZN(n34077) );
  OAI222_X1 U34240 ( .A1(n31462), .A2(n39684), .B1(n31526), .B2(n39678), .C1(
        n31398), .C2(n39672), .ZN(n34084) );
  AOI221_X1 U34241 ( .B1(n39324), .B2(n32537), .C1(n39318), .C2(n27975), .A(
        n35366), .ZN(n35359) );
  OAI222_X1 U34242 ( .A1(n30576), .A2(n39312), .B1(n30640), .B2(n39306), .C1(
        n30512), .C2(n39300), .ZN(n35366) );
  AOI221_X1 U34243 ( .B1(n39444), .B2(n29074), .C1(n39438), .C2(n29138), .A(
        n35358), .ZN(n35351) );
  OAI222_X1 U34244 ( .A1(n31462), .A2(n39432), .B1(n31526), .B2(n39426), .C1(
        n31398), .C2(n39420), .ZN(n35358) );
  AOI221_X1 U34245 ( .B1(n39576), .B2(n32536), .C1(n39570), .C2(n27974), .A(
        n34111), .ZN(n34104) );
  OAI222_X1 U34246 ( .A1(n30575), .A2(n39564), .B1(n30639), .B2(n39558), .C1(
        n30511), .C2(n39552), .ZN(n34111) );
  AOI221_X1 U34247 ( .B1(n39696), .B2(n29073), .C1(n39690), .C2(n29137), .A(
        n34103), .ZN(n34096) );
  OAI222_X1 U34248 ( .A1(n31461), .A2(n39684), .B1(n31525), .B2(n39678), .C1(
        n31397), .C2(n39672), .ZN(n34103) );
  AOI221_X1 U34249 ( .B1(n39324), .B2(n32536), .C1(n39318), .C2(n27974), .A(
        n35385), .ZN(n35378) );
  OAI222_X1 U34250 ( .A1(n30575), .A2(n39312), .B1(n30639), .B2(n39306), .C1(
        n30511), .C2(n39300), .ZN(n35385) );
  AOI221_X1 U34251 ( .B1(n39444), .B2(n29073), .C1(n39438), .C2(n29137), .A(
        n35377), .ZN(n35370) );
  OAI222_X1 U34252 ( .A1(n31461), .A2(n39432), .B1(n31525), .B2(n39426), .C1(
        n31397), .C2(n39420), .ZN(n35377) );
  AOI221_X1 U34253 ( .B1(n39576), .B2(n32535), .C1(n39570), .C2(n27973), .A(
        n34130), .ZN(n34123) );
  OAI222_X1 U34254 ( .A1(n30574), .A2(n39564), .B1(n30638), .B2(n39558), .C1(
        n30510), .C2(n39552), .ZN(n34130) );
  AOI221_X1 U34255 ( .B1(n39696), .B2(n29072), .C1(n39690), .C2(n29136), .A(
        n34122), .ZN(n34115) );
  OAI222_X1 U34256 ( .A1(n31460), .A2(n39684), .B1(n31524), .B2(n39678), .C1(
        n31396), .C2(n39672), .ZN(n34122) );
  AOI221_X1 U34257 ( .B1(n39324), .B2(n32535), .C1(n39318), .C2(n27973), .A(
        n35404), .ZN(n35397) );
  OAI222_X1 U34258 ( .A1(n30574), .A2(n39312), .B1(n30638), .B2(n39306), .C1(
        n30510), .C2(n39300), .ZN(n35404) );
  AOI221_X1 U34259 ( .B1(n39444), .B2(n29072), .C1(n39438), .C2(n29136), .A(
        n35396), .ZN(n35389) );
  OAI222_X1 U34260 ( .A1(n31460), .A2(n39432), .B1(n31524), .B2(n39426), .C1(
        n31396), .C2(n39420), .ZN(n35396) );
  AOI221_X1 U34261 ( .B1(n39576), .B2(n32534), .C1(n39570), .C2(n27972), .A(
        n34149), .ZN(n34142) );
  OAI222_X1 U34262 ( .A1(n30573), .A2(n39564), .B1(n30637), .B2(n39558), .C1(
        n30509), .C2(n39552), .ZN(n34149) );
  AOI221_X1 U34263 ( .B1(n39696), .B2(n29071), .C1(n39690), .C2(n29135), .A(
        n34141), .ZN(n34134) );
  OAI222_X1 U34264 ( .A1(n31459), .A2(n39684), .B1(n31523), .B2(n39678), .C1(
        n31395), .C2(n39672), .ZN(n34141) );
  AOI221_X1 U34265 ( .B1(n39324), .B2(n32534), .C1(n39318), .C2(n27972), .A(
        n35423), .ZN(n35416) );
  OAI222_X1 U34266 ( .A1(n30573), .A2(n39312), .B1(n30637), .B2(n39306), .C1(
        n30509), .C2(n39300), .ZN(n35423) );
  AOI221_X1 U34267 ( .B1(n39444), .B2(n29071), .C1(n39438), .C2(n29135), .A(
        n35415), .ZN(n35408) );
  OAI222_X1 U34268 ( .A1(n31459), .A2(n39432), .B1(n31523), .B2(n39426), .C1(
        n31395), .C2(n39420), .ZN(n35415) );
  AOI221_X1 U34269 ( .B1(n39576), .B2(n32533), .C1(n39570), .C2(n27971), .A(
        n34168), .ZN(n34161) );
  OAI222_X1 U34270 ( .A1(n30572), .A2(n39564), .B1(n30636), .B2(n39558), .C1(
        n30508), .C2(n39552), .ZN(n34168) );
  AOI221_X1 U34271 ( .B1(n39696), .B2(n29070), .C1(n39690), .C2(n29134), .A(
        n34160), .ZN(n34153) );
  OAI222_X1 U34272 ( .A1(n31458), .A2(n39684), .B1(n31522), .B2(n39678), .C1(
        n31394), .C2(n39672), .ZN(n34160) );
  AOI221_X1 U34273 ( .B1(n39324), .B2(n32533), .C1(n39318), .C2(n27971), .A(
        n35442), .ZN(n35435) );
  OAI222_X1 U34274 ( .A1(n30572), .A2(n39312), .B1(n30636), .B2(n39306), .C1(
        n30508), .C2(n39300), .ZN(n35442) );
  AOI221_X1 U34275 ( .B1(n39444), .B2(n29070), .C1(n39438), .C2(n29134), .A(
        n35434), .ZN(n35427) );
  OAI222_X1 U34276 ( .A1(n31458), .A2(n39432), .B1(n31522), .B2(n39426), .C1(
        n31394), .C2(n39420), .ZN(n35434) );
  AOI221_X1 U34277 ( .B1(n39576), .B2(n32532), .C1(n39570), .C2(n27970), .A(
        n34187), .ZN(n34180) );
  OAI222_X1 U34278 ( .A1(n30571), .A2(n39564), .B1(n30635), .B2(n39558), .C1(
        n30507), .C2(n39552), .ZN(n34187) );
  AOI221_X1 U34279 ( .B1(n39696), .B2(n29069), .C1(n39690), .C2(n29133), .A(
        n34179), .ZN(n34172) );
  OAI222_X1 U34280 ( .A1(n31457), .A2(n39684), .B1(n31521), .B2(n39678), .C1(
        n31393), .C2(n39672), .ZN(n34179) );
  AOI221_X1 U34281 ( .B1(n39324), .B2(n32532), .C1(n39318), .C2(n27970), .A(
        n35461), .ZN(n35454) );
  OAI222_X1 U34282 ( .A1(n30571), .A2(n39312), .B1(n30635), .B2(n39306), .C1(
        n30507), .C2(n39300), .ZN(n35461) );
  AOI221_X1 U34283 ( .B1(n39444), .B2(n29069), .C1(n39438), .C2(n29133), .A(
        n35453), .ZN(n35446) );
  OAI222_X1 U34284 ( .A1(n31457), .A2(n39432), .B1(n31521), .B2(n39426), .C1(
        n31393), .C2(n39420), .ZN(n35453) );
  AOI221_X1 U34285 ( .B1(n39576), .B2(n32531), .C1(n39570), .C2(n27969), .A(
        n34206), .ZN(n34199) );
  OAI222_X1 U34286 ( .A1(n30570), .A2(n39564), .B1(n30634), .B2(n39558), .C1(
        n30506), .C2(n39552), .ZN(n34206) );
  AOI221_X1 U34287 ( .B1(n39696), .B2(n29068), .C1(n39690), .C2(n29132), .A(
        n34198), .ZN(n34191) );
  OAI222_X1 U34288 ( .A1(n31456), .A2(n39684), .B1(n31520), .B2(n39678), .C1(
        n31392), .C2(n39672), .ZN(n34198) );
  AOI221_X1 U34289 ( .B1(n39324), .B2(n32531), .C1(n39318), .C2(n27969), .A(
        n35480), .ZN(n35473) );
  OAI222_X1 U34290 ( .A1(n30570), .A2(n39312), .B1(n30634), .B2(n39306), .C1(
        n30506), .C2(n39300), .ZN(n35480) );
  AOI221_X1 U34291 ( .B1(n39444), .B2(n29068), .C1(n39438), .C2(n29132), .A(
        n35472), .ZN(n35465) );
  OAI222_X1 U34292 ( .A1(n31456), .A2(n39432), .B1(n31520), .B2(n39426), .C1(
        n31392), .C2(n39420), .ZN(n35472) );
  AOI221_X1 U34293 ( .B1(n39576), .B2(n32530), .C1(n39570), .C2(n27968), .A(
        n34225), .ZN(n34218) );
  OAI222_X1 U34294 ( .A1(n30569), .A2(n39564), .B1(n30633), .B2(n39558), .C1(
        n30505), .C2(n39552), .ZN(n34225) );
  AOI221_X1 U34295 ( .B1(n39696), .B2(n29067), .C1(n39690), .C2(n29131), .A(
        n34217), .ZN(n34210) );
  OAI222_X1 U34296 ( .A1(n31455), .A2(n39684), .B1(n31519), .B2(n39678), .C1(
        n31391), .C2(n39672), .ZN(n34217) );
  AOI221_X1 U34297 ( .B1(n39324), .B2(n32530), .C1(n39318), .C2(n27968), .A(
        n35499), .ZN(n35492) );
  OAI222_X1 U34298 ( .A1(n30569), .A2(n39312), .B1(n30633), .B2(n39306), .C1(
        n30505), .C2(n39300), .ZN(n35499) );
  AOI221_X1 U34299 ( .B1(n39444), .B2(n29067), .C1(n39438), .C2(n29131), .A(
        n35491), .ZN(n35484) );
  OAI222_X1 U34300 ( .A1(n31455), .A2(n39432), .B1(n31519), .B2(n39426), .C1(
        n31391), .C2(n39420), .ZN(n35491) );
  AOI221_X1 U34301 ( .B1(n39575), .B2(n32529), .C1(n39569), .C2(n27967), .A(
        n34244), .ZN(n34237) );
  OAI222_X1 U34302 ( .A1(n30568), .A2(n39563), .B1(n30632), .B2(n39557), .C1(
        n30504), .C2(n39551), .ZN(n34244) );
  AOI221_X1 U34303 ( .B1(n39695), .B2(n29066), .C1(n39689), .C2(n29130), .A(
        n34236), .ZN(n34229) );
  OAI222_X1 U34304 ( .A1(n31454), .A2(n39683), .B1(n31518), .B2(n39677), .C1(
        n31390), .C2(n39671), .ZN(n34236) );
  AOI221_X1 U34305 ( .B1(n39323), .B2(n32529), .C1(n39317), .C2(n27967), .A(
        n35518), .ZN(n35511) );
  OAI222_X1 U34306 ( .A1(n30568), .A2(n39311), .B1(n30632), .B2(n39305), .C1(
        n30504), .C2(n39299), .ZN(n35518) );
  AOI221_X1 U34307 ( .B1(n39443), .B2(n29066), .C1(n39437), .C2(n29130), .A(
        n35510), .ZN(n35503) );
  OAI222_X1 U34308 ( .A1(n31454), .A2(n39431), .B1(n31518), .B2(n39425), .C1(
        n31390), .C2(n39419), .ZN(n35510) );
  AOI221_X1 U34309 ( .B1(n39575), .B2(n32528), .C1(n39569), .C2(n27966), .A(
        n34263), .ZN(n34256) );
  OAI222_X1 U34310 ( .A1(n30567), .A2(n39563), .B1(n30631), .B2(n39557), .C1(
        n30503), .C2(n39551), .ZN(n34263) );
  AOI221_X1 U34311 ( .B1(n39695), .B2(n29065), .C1(n39689), .C2(n29129), .A(
        n34255), .ZN(n34248) );
  OAI222_X1 U34312 ( .A1(n31453), .A2(n39683), .B1(n31517), .B2(n39677), .C1(
        n31389), .C2(n39671), .ZN(n34255) );
  AOI221_X1 U34313 ( .B1(n39323), .B2(n32528), .C1(n39317), .C2(n27966), .A(
        n35537), .ZN(n35530) );
  OAI222_X1 U34314 ( .A1(n30567), .A2(n39311), .B1(n30631), .B2(n39305), .C1(
        n30503), .C2(n39299), .ZN(n35537) );
  AOI221_X1 U34315 ( .B1(n39443), .B2(n29065), .C1(n39437), .C2(n29129), .A(
        n35529), .ZN(n35522) );
  OAI222_X1 U34316 ( .A1(n31453), .A2(n39431), .B1(n31517), .B2(n39425), .C1(
        n31389), .C2(n39419), .ZN(n35529) );
  AOI221_X1 U34317 ( .B1(n39575), .B2(n32527), .C1(n39569), .C2(n27965), .A(
        n34282), .ZN(n34275) );
  OAI222_X1 U34318 ( .A1(n30566), .A2(n39563), .B1(n30630), .B2(n39557), .C1(
        n30502), .C2(n39551), .ZN(n34282) );
  AOI221_X1 U34319 ( .B1(n39695), .B2(n29064), .C1(n39689), .C2(n29128), .A(
        n34274), .ZN(n34267) );
  OAI222_X1 U34320 ( .A1(n31452), .A2(n39683), .B1(n31516), .B2(n39677), .C1(
        n31388), .C2(n39671), .ZN(n34274) );
  AOI221_X1 U34321 ( .B1(n39323), .B2(n32527), .C1(n39317), .C2(n27965), .A(
        n35556), .ZN(n35549) );
  OAI222_X1 U34322 ( .A1(n30566), .A2(n39311), .B1(n30630), .B2(n39305), .C1(
        n30502), .C2(n39299), .ZN(n35556) );
  AOI221_X1 U34323 ( .B1(n39443), .B2(n29064), .C1(n39437), .C2(n29128), .A(
        n35548), .ZN(n35541) );
  OAI222_X1 U34324 ( .A1(n31452), .A2(n39431), .B1(n31516), .B2(n39425), .C1(
        n31388), .C2(n39419), .ZN(n35548) );
  AOI221_X1 U34325 ( .B1(n39575), .B2(n32526), .C1(n39569), .C2(n27964), .A(
        n34301), .ZN(n34294) );
  OAI222_X1 U34326 ( .A1(n30565), .A2(n39563), .B1(n30629), .B2(n39557), .C1(
        n30501), .C2(n39551), .ZN(n34301) );
  AOI221_X1 U34327 ( .B1(n39695), .B2(n29063), .C1(n39689), .C2(n29127), .A(
        n34293), .ZN(n34286) );
  OAI222_X1 U34328 ( .A1(n31451), .A2(n39683), .B1(n31515), .B2(n39677), .C1(
        n31387), .C2(n39671), .ZN(n34293) );
  AOI221_X1 U34329 ( .B1(n39323), .B2(n32526), .C1(n39317), .C2(n27964), .A(
        n35575), .ZN(n35568) );
  OAI222_X1 U34330 ( .A1(n30565), .A2(n39311), .B1(n30629), .B2(n39305), .C1(
        n30501), .C2(n39299), .ZN(n35575) );
  AOI221_X1 U34331 ( .B1(n39443), .B2(n29063), .C1(n39437), .C2(n29127), .A(
        n35567), .ZN(n35560) );
  OAI222_X1 U34332 ( .A1(n31451), .A2(n39431), .B1(n31515), .B2(n39425), .C1(
        n31387), .C2(n39419), .ZN(n35567) );
  AOI221_X1 U34333 ( .B1(n39575), .B2(n32525), .C1(n39569), .C2(n27963), .A(
        n34320), .ZN(n34313) );
  OAI222_X1 U34334 ( .A1(n30564), .A2(n39563), .B1(n30628), .B2(n39557), .C1(
        n30500), .C2(n39551), .ZN(n34320) );
  AOI221_X1 U34335 ( .B1(n39695), .B2(n29062), .C1(n39689), .C2(n29126), .A(
        n34312), .ZN(n34305) );
  OAI222_X1 U34336 ( .A1(n31450), .A2(n39683), .B1(n31514), .B2(n39677), .C1(
        n31386), .C2(n39671), .ZN(n34312) );
  AOI221_X1 U34337 ( .B1(n39323), .B2(n32525), .C1(n39317), .C2(n27963), .A(
        n35594), .ZN(n35587) );
  OAI222_X1 U34338 ( .A1(n30564), .A2(n39311), .B1(n30628), .B2(n39305), .C1(
        n30500), .C2(n39299), .ZN(n35594) );
  AOI221_X1 U34339 ( .B1(n39443), .B2(n29062), .C1(n39437), .C2(n29126), .A(
        n35586), .ZN(n35579) );
  OAI222_X1 U34340 ( .A1(n31450), .A2(n39431), .B1(n31514), .B2(n39425), .C1(
        n31386), .C2(n39419), .ZN(n35586) );
  AOI221_X1 U34341 ( .B1(n39575), .B2(n32524), .C1(n39569), .C2(n27962), .A(
        n34339), .ZN(n34332) );
  OAI222_X1 U34342 ( .A1(n30563), .A2(n39563), .B1(n30627), .B2(n39557), .C1(
        n30499), .C2(n39551), .ZN(n34339) );
  AOI221_X1 U34343 ( .B1(n39695), .B2(n29061), .C1(n39689), .C2(n29125), .A(
        n34331), .ZN(n34324) );
  OAI222_X1 U34344 ( .A1(n31449), .A2(n39683), .B1(n31513), .B2(n39677), .C1(
        n31385), .C2(n39671), .ZN(n34331) );
  AOI221_X1 U34345 ( .B1(n39323), .B2(n32524), .C1(n39317), .C2(n27962), .A(
        n35613), .ZN(n35606) );
  OAI222_X1 U34346 ( .A1(n30563), .A2(n39311), .B1(n30627), .B2(n39305), .C1(
        n30499), .C2(n39299), .ZN(n35613) );
  AOI221_X1 U34347 ( .B1(n39443), .B2(n29061), .C1(n39437), .C2(n29125), .A(
        n35605), .ZN(n35598) );
  OAI222_X1 U34348 ( .A1(n31449), .A2(n39431), .B1(n31513), .B2(n39425), .C1(
        n31385), .C2(n39419), .ZN(n35605) );
  AOI221_X1 U34349 ( .B1(n39575), .B2(n32523), .C1(n39569), .C2(n27961), .A(
        n34358), .ZN(n34351) );
  OAI222_X1 U34350 ( .A1(n30562), .A2(n39563), .B1(n30626), .B2(n39557), .C1(
        n30498), .C2(n39551), .ZN(n34358) );
  AOI221_X1 U34351 ( .B1(n39695), .B2(n29060), .C1(n39689), .C2(n29124), .A(
        n34350), .ZN(n34343) );
  OAI222_X1 U34352 ( .A1(n31448), .A2(n39683), .B1(n31512), .B2(n39677), .C1(
        n31384), .C2(n39671), .ZN(n34350) );
  AOI221_X1 U34353 ( .B1(n39323), .B2(n32523), .C1(n39317), .C2(n27961), .A(
        n35632), .ZN(n35625) );
  OAI222_X1 U34354 ( .A1(n30562), .A2(n39311), .B1(n30626), .B2(n39305), .C1(
        n30498), .C2(n39299), .ZN(n35632) );
  AOI221_X1 U34355 ( .B1(n39443), .B2(n29060), .C1(n39437), .C2(n29124), .A(
        n35624), .ZN(n35617) );
  OAI222_X1 U34356 ( .A1(n31448), .A2(n39431), .B1(n31512), .B2(n39425), .C1(
        n31384), .C2(n39419), .ZN(n35624) );
  AOI221_X1 U34357 ( .B1(n39575), .B2(n32522), .C1(n39569), .C2(n27960), .A(
        n34377), .ZN(n34370) );
  OAI222_X1 U34358 ( .A1(n30561), .A2(n39563), .B1(n30625), .B2(n39557), .C1(
        n30497), .C2(n39551), .ZN(n34377) );
  AOI221_X1 U34359 ( .B1(n39695), .B2(n29059), .C1(n39689), .C2(n29123), .A(
        n34369), .ZN(n34362) );
  OAI222_X1 U34360 ( .A1(n31447), .A2(n39683), .B1(n31511), .B2(n39677), .C1(
        n31383), .C2(n39671), .ZN(n34369) );
  AOI221_X1 U34361 ( .B1(n39323), .B2(n32522), .C1(n39317), .C2(n27960), .A(
        n35651), .ZN(n35644) );
  OAI222_X1 U34362 ( .A1(n30561), .A2(n39311), .B1(n30625), .B2(n39305), .C1(
        n30497), .C2(n39299), .ZN(n35651) );
  AOI221_X1 U34363 ( .B1(n39443), .B2(n29059), .C1(n39437), .C2(n29123), .A(
        n35643), .ZN(n35636) );
  OAI222_X1 U34364 ( .A1(n31447), .A2(n39431), .B1(n31511), .B2(n39425), .C1(
        n31383), .C2(n39419), .ZN(n35643) );
  AOI221_X1 U34365 ( .B1(n39575), .B2(n32521), .C1(n39569), .C2(n27959), .A(
        n34396), .ZN(n34389) );
  OAI222_X1 U34366 ( .A1(n30560), .A2(n39563), .B1(n30624), .B2(n39557), .C1(
        n30496), .C2(n39551), .ZN(n34396) );
  AOI221_X1 U34367 ( .B1(n39695), .B2(n29058), .C1(n39689), .C2(n29122), .A(
        n34388), .ZN(n34381) );
  OAI222_X1 U34368 ( .A1(n31446), .A2(n39683), .B1(n31510), .B2(n39677), .C1(
        n31382), .C2(n39671), .ZN(n34388) );
  AOI221_X1 U34369 ( .B1(n39323), .B2(n32521), .C1(n39317), .C2(n27959), .A(
        n35670), .ZN(n35663) );
  OAI222_X1 U34370 ( .A1(n30560), .A2(n39311), .B1(n30624), .B2(n39305), .C1(
        n30496), .C2(n39299), .ZN(n35670) );
  AOI221_X1 U34371 ( .B1(n39443), .B2(n29058), .C1(n39437), .C2(n29122), .A(
        n35662), .ZN(n35655) );
  OAI222_X1 U34372 ( .A1(n31446), .A2(n39431), .B1(n31510), .B2(n39425), .C1(
        n31382), .C2(n39419), .ZN(n35662) );
  AOI221_X1 U34373 ( .B1(n39575), .B2(n32520), .C1(n39569), .C2(n27958), .A(
        n34415), .ZN(n34408) );
  OAI222_X1 U34374 ( .A1(n30559), .A2(n39563), .B1(n30623), .B2(n39557), .C1(
        n30495), .C2(n39551), .ZN(n34415) );
  AOI221_X1 U34375 ( .B1(n39695), .B2(n29057), .C1(n39689), .C2(n29121), .A(
        n34407), .ZN(n34400) );
  OAI222_X1 U34376 ( .A1(n31445), .A2(n39683), .B1(n31509), .B2(n39677), .C1(
        n31381), .C2(n39671), .ZN(n34407) );
  AOI221_X1 U34377 ( .B1(n39323), .B2(n32520), .C1(n39317), .C2(n27958), .A(
        n35689), .ZN(n35682) );
  OAI222_X1 U34378 ( .A1(n30559), .A2(n39311), .B1(n30623), .B2(n39305), .C1(
        n30495), .C2(n39299), .ZN(n35689) );
  AOI221_X1 U34379 ( .B1(n39443), .B2(n29057), .C1(n39437), .C2(n29121), .A(
        n35681), .ZN(n35674) );
  OAI222_X1 U34380 ( .A1(n31445), .A2(n39431), .B1(n31509), .B2(n39425), .C1(
        n31381), .C2(n39419), .ZN(n35681) );
  AOI221_X1 U34381 ( .B1(n39575), .B2(n32519), .C1(n39569), .C2(n27957), .A(
        n34434), .ZN(n34427) );
  OAI222_X1 U34382 ( .A1(n30558), .A2(n39563), .B1(n30622), .B2(n39557), .C1(
        n30494), .C2(n39551), .ZN(n34434) );
  AOI221_X1 U34383 ( .B1(n39695), .B2(n29056), .C1(n39689), .C2(n29120), .A(
        n34426), .ZN(n34419) );
  OAI222_X1 U34384 ( .A1(n31444), .A2(n39683), .B1(n31508), .B2(n39677), .C1(
        n31380), .C2(n39671), .ZN(n34426) );
  AOI221_X1 U34385 ( .B1(n39323), .B2(n32519), .C1(n39317), .C2(n27957), .A(
        n35708), .ZN(n35701) );
  OAI222_X1 U34386 ( .A1(n30558), .A2(n39311), .B1(n30622), .B2(n39305), .C1(
        n30494), .C2(n39299), .ZN(n35708) );
  AOI221_X1 U34387 ( .B1(n39443), .B2(n29056), .C1(n39437), .C2(n29120), .A(
        n35700), .ZN(n35693) );
  OAI222_X1 U34388 ( .A1(n31444), .A2(n39431), .B1(n31508), .B2(n39425), .C1(
        n31380), .C2(n39419), .ZN(n35700) );
  AOI221_X1 U34389 ( .B1(n39575), .B2(n32518), .C1(n39569), .C2(n27956), .A(
        n34453), .ZN(n34446) );
  OAI222_X1 U34390 ( .A1(n30557), .A2(n39563), .B1(n30621), .B2(n39557), .C1(
        n30493), .C2(n39551), .ZN(n34453) );
  AOI221_X1 U34391 ( .B1(n39695), .B2(n29055), .C1(n39689), .C2(n29119), .A(
        n34445), .ZN(n34438) );
  OAI222_X1 U34392 ( .A1(n31443), .A2(n39683), .B1(n31507), .B2(n39677), .C1(
        n31379), .C2(n39671), .ZN(n34445) );
  AOI221_X1 U34393 ( .B1(n39323), .B2(n32518), .C1(n39317), .C2(n27956), .A(
        n35727), .ZN(n35720) );
  OAI222_X1 U34394 ( .A1(n30557), .A2(n39311), .B1(n30621), .B2(n39305), .C1(
        n30493), .C2(n39299), .ZN(n35727) );
  AOI221_X1 U34395 ( .B1(n39443), .B2(n29055), .C1(n39437), .C2(n29119), .A(
        n35719), .ZN(n35712) );
  OAI222_X1 U34396 ( .A1(n31443), .A2(n39431), .B1(n31507), .B2(n39425), .C1(
        n31379), .C2(n39419), .ZN(n35719) );
  AOI221_X1 U34397 ( .B1(n39574), .B2(n32517), .C1(n39568), .C2(n27955), .A(
        n34472), .ZN(n34465) );
  OAI222_X1 U34398 ( .A1(n30556), .A2(n39562), .B1(n30620), .B2(n39556), .C1(
        n30492), .C2(n39550), .ZN(n34472) );
  AOI221_X1 U34399 ( .B1(n39694), .B2(n29054), .C1(n39688), .C2(n29118), .A(
        n34464), .ZN(n34457) );
  OAI222_X1 U34400 ( .A1(n31442), .A2(n39682), .B1(n31506), .B2(n39676), .C1(
        n31378), .C2(n39670), .ZN(n34464) );
  AOI221_X1 U34401 ( .B1(n39322), .B2(n32517), .C1(n39316), .C2(n27955), .A(
        n35746), .ZN(n35739) );
  OAI222_X1 U34402 ( .A1(n30556), .A2(n39310), .B1(n30620), .B2(n39304), .C1(
        n30492), .C2(n39298), .ZN(n35746) );
  AOI221_X1 U34403 ( .B1(n39442), .B2(n29054), .C1(n39436), .C2(n29118), .A(
        n35738), .ZN(n35731) );
  OAI222_X1 U34404 ( .A1(n31442), .A2(n39430), .B1(n31506), .B2(n39424), .C1(
        n31378), .C2(n39418), .ZN(n35738) );
  AOI221_X1 U34405 ( .B1(n39574), .B2(n32516), .C1(n39568), .C2(n27954), .A(
        n34491), .ZN(n34484) );
  OAI222_X1 U34406 ( .A1(n30555), .A2(n39562), .B1(n30619), .B2(n39556), .C1(
        n30491), .C2(n39550), .ZN(n34491) );
  AOI221_X1 U34407 ( .B1(n39694), .B2(n29053), .C1(n39688), .C2(n29117), .A(
        n34483), .ZN(n34476) );
  OAI222_X1 U34408 ( .A1(n31441), .A2(n39682), .B1(n31505), .B2(n39676), .C1(
        n31377), .C2(n39670), .ZN(n34483) );
  AOI221_X1 U34409 ( .B1(n39322), .B2(n32516), .C1(n39316), .C2(n27954), .A(
        n35765), .ZN(n35758) );
  OAI222_X1 U34410 ( .A1(n30555), .A2(n39310), .B1(n30619), .B2(n39304), .C1(
        n30491), .C2(n39298), .ZN(n35765) );
  AOI221_X1 U34411 ( .B1(n39442), .B2(n29053), .C1(n39436), .C2(n29117), .A(
        n35757), .ZN(n35750) );
  OAI222_X1 U34412 ( .A1(n31441), .A2(n39430), .B1(n31505), .B2(n39424), .C1(
        n31377), .C2(n39418), .ZN(n35757) );
  AOI221_X1 U34413 ( .B1(n39574), .B2(n32515), .C1(n39568), .C2(n27953), .A(
        n34510), .ZN(n34503) );
  OAI222_X1 U34414 ( .A1(n30554), .A2(n39562), .B1(n30618), .B2(n39556), .C1(
        n30490), .C2(n39550), .ZN(n34510) );
  AOI221_X1 U34415 ( .B1(n39694), .B2(n29052), .C1(n39688), .C2(n29116), .A(
        n34502), .ZN(n34495) );
  OAI222_X1 U34416 ( .A1(n31440), .A2(n39682), .B1(n31504), .B2(n39676), .C1(
        n31376), .C2(n39670), .ZN(n34502) );
  AOI221_X1 U34417 ( .B1(n39322), .B2(n32515), .C1(n39316), .C2(n27953), .A(
        n35784), .ZN(n35777) );
  OAI222_X1 U34418 ( .A1(n30554), .A2(n39310), .B1(n30618), .B2(n39304), .C1(
        n30490), .C2(n39298), .ZN(n35784) );
  AOI221_X1 U34419 ( .B1(n39442), .B2(n29052), .C1(n39436), .C2(n29116), .A(
        n35776), .ZN(n35769) );
  OAI222_X1 U34420 ( .A1(n31440), .A2(n39430), .B1(n31504), .B2(n39424), .C1(
        n31376), .C2(n39418), .ZN(n35776) );
  AOI221_X1 U34421 ( .B1(n39574), .B2(n32514), .C1(n39568), .C2(n27952), .A(
        n34529), .ZN(n34522) );
  OAI222_X1 U34422 ( .A1(n30553), .A2(n39562), .B1(n30617), .B2(n39556), .C1(
        n30489), .C2(n39550), .ZN(n34529) );
  AOI221_X1 U34423 ( .B1(n39694), .B2(n29051), .C1(n39688), .C2(n29115), .A(
        n34521), .ZN(n34514) );
  OAI222_X1 U34424 ( .A1(n31439), .A2(n39682), .B1(n31503), .B2(n39676), .C1(
        n31375), .C2(n39670), .ZN(n34521) );
  AOI221_X1 U34425 ( .B1(n39322), .B2(n32514), .C1(n39316), .C2(n27952), .A(
        n35803), .ZN(n35796) );
  OAI222_X1 U34426 ( .A1(n30553), .A2(n39310), .B1(n30617), .B2(n39304), .C1(
        n30489), .C2(n39298), .ZN(n35803) );
  AOI221_X1 U34427 ( .B1(n39442), .B2(n29051), .C1(n39436), .C2(n29115), .A(
        n35795), .ZN(n35788) );
  OAI222_X1 U34428 ( .A1(n31439), .A2(n39430), .B1(n31503), .B2(n39424), .C1(
        n31375), .C2(n39418), .ZN(n35795) );
  AOI221_X1 U34429 ( .B1(n39574), .B2(n32513), .C1(n39568), .C2(n27951), .A(
        n34548), .ZN(n34541) );
  OAI222_X1 U34430 ( .A1(n30552), .A2(n39562), .B1(n30616), .B2(n39556), .C1(
        n30488), .C2(n39550), .ZN(n34548) );
  AOI221_X1 U34431 ( .B1(n39694), .B2(n29050), .C1(n39688), .C2(n29114), .A(
        n34540), .ZN(n34533) );
  OAI222_X1 U34432 ( .A1(n31438), .A2(n39682), .B1(n31502), .B2(n39676), .C1(
        n31374), .C2(n39670), .ZN(n34540) );
  AOI221_X1 U34433 ( .B1(n39322), .B2(n32513), .C1(n39316), .C2(n27951), .A(
        n35822), .ZN(n35815) );
  OAI222_X1 U34434 ( .A1(n30552), .A2(n39310), .B1(n30616), .B2(n39304), .C1(
        n30488), .C2(n39298), .ZN(n35822) );
  AOI221_X1 U34435 ( .B1(n39442), .B2(n29050), .C1(n39436), .C2(n29114), .A(
        n35814), .ZN(n35807) );
  OAI222_X1 U34436 ( .A1(n31438), .A2(n39430), .B1(n31502), .B2(n39424), .C1(
        n31374), .C2(n39418), .ZN(n35814) );
  AOI221_X1 U34437 ( .B1(n39574), .B2(n32512), .C1(n39568), .C2(n27950), .A(
        n34567), .ZN(n34560) );
  OAI222_X1 U34438 ( .A1(n30551), .A2(n39562), .B1(n30615), .B2(n39556), .C1(
        n30487), .C2(n39550), .ZN(n34567) );
  AOI221_X1 U34439 ( .B1(n39694), .B2(n29049), .C1(n39688), .C2(n29113), .A(
        n34559), .ZN(n34552) );
  OAI222_X1 U34440 ( .A1(n31437), .A2(n39682), .B1(n31501), .B2(n39676), .C1(
        n31373), .C2(n39670), .ZN(n34559) );
  AOI221_X1 U34441 ( .B1(n39322), .B2(n32512), .C1(n39316), .C2(n27950), .A(
        n35841), .ZN(n35834) );
  OAI222_X1 U34442 ( .A1(n30551), .A2(n39310), .B1(n30615), .B2(n39304), .C1(
        n30487), .C2(n39298), .ZN(n35841) );
  AOI221_X1 U34443 ( .B1(n39442), .B2(n29049), .C1(n39436), .C2(n29113), .A(
        n35833), .ZN(n35826) );
  OAI222_X1 U34444 ( .A1(n31437), .A2(n39430), .B1(n31501), .B2(n39424), .C1(
        n31373), .C2(n39418), .ZN(n35833) );
  AOI221_X1 U34445 ( .B1(n39574), .B2(n32511), .C1(n39568), .C2(n27949), .A(
        n34586), .ZN(n34579) );
  OAI222_X1 U34446 ( .A1(n30550), .A2(n39562), .B1(n30614), .B2(n39556), .C1(
        n30486), .C2(n39550), .ZN(n34586) );
  AOI221_X1 U34447 ( .B1(n39694), .B2(n29048), .C1(n39688), .C2(n29112), .A(
        n34578), .ZN(n34571) );
  OAI222_X1 U34448 ( .A1(n31436), .A2(n39682), .B1(n31500), .B2(n39676), .C1(
        n31372), .C2(n39670), .ZN(n34578) );
  AOI221_X1 U34449 ( .B1(n39322), .B2(n32511), .C1(n39316), .C2(n27949), .A(
        n35860), .ZN(n35853) );
  OAI222_X1 U34450 ( .A1(n30550), .A2(n39310), .B1(n30614), .B2(n39304), .C1(
        n30486), .C2(n39298), .ZN(n35860) );
  AOI221_X1 U34451 ( .B1(n39442), .B2(n29048), .C1(n39436), .C2(n29112), .A(
        n35852), .ZN(n35845) );
  OAI222_X1 U34452 ( .A1(n31436), .A2(n39430), .B1(n31500), .B2(n39424), .C1(
        n31372), .C2(n39418), .ZN(n35852) );
  AOI221_X1 U34453 ( .B1(n39574), .B2(n32510), .C1(n39568), .C2(n27948), .A(
        n34605), .ZN(n34598) );
  OAI222_X1 U34454 ( .A1(n30549), .A2(n39562), .B1(n30613), .B2(n39556), .C1(
        n30485), .C2(n39550), .ZN(n34605) );
  AOI221_X1 U34455 ( .B1(n39694), .B2(n29047), .C1(n39688), .C2(n29111), .A(
        n34597), .ZN(n34590) );
  OAI222_X1 U34456 ( .A1(n31435), .A2(n39682), .B1(n31499), .B2(n39676), .C1(
        n31371), .C2(n39670), .ZN(n34597) );
  AOI221_X1 U34457 ( .B1(n39322), .B2(n32510), .C1(n39316), .C2(n27948), .A(
        n35879), .ZN(n35872) );
  OAI222_X1 U34458 ( .A1(n30549), .A2(n39310), .B1(n30613), .B2(n39304), .C1(
        n30485), .C2(n39298), .ZN(n35879) );
  AOI221_X1 U34459 ( .B1(n39442), .B2(n29047), .C1(n39436), .C2(n29111), .A(
        n35871), .ZN(n35864) );
  OAI222_X1 U34460 ( .A1(n31435), .A2(n39430), .B1(n31499), .B2(n39424), .C1(
        n31371), .C2(n39418), .ZN(n35871) );
  AOI221_X1 U34461 ( .B1(n39574), .B2(n32507), .C1(n39568), .C2(n27947), .A(
        n34624), .ZN(n34617) );
  OAI222_X1 U34462 ( .A1(n30548), .A2(n39562), .B1(n30612), .B2(n39556), .C1(
        n30484), .C2(n39550), .ZN(n34624) );
  AOI221_X1 U34463 ( .B1(n39694), .B2(n29046), .C1(n39688), .C2(n29110), .A(
        n34616), .ZN(n34609) );
  OAI222_X1 U34464 ( .A1(n31434), .A2(n39682), .B1(n31498), .B2(n39676), .C1(
        n31370), .C2(n39670), .ZN(n34616) );
  AOI221_X1 U34465 ( .B1(n39322), .B2(n32507), .C1(n39316), .C2(n27947), .A(
        n35898), .ZN(n35891) );
  OAI222_X1 U34466 ( .A1(n30548), .A2(n39310), .B1(n30612), .B2(n39304), .C1(
        n30484), .C2(n39298), .ZN(n35898) );
  AOI221_X1 U34467 ( .B1(n39442), .B2(n29046), .C1(n39436), .C2(n29110), .A(
        n35890), .ZN(n35883) );
  OAI222_X1 U34468 ( .A1(n31434), .A2(n39430), .B1(n31498), .B2(n39424), .C1(
        n31370), .C2(n39418), .ZN(n35890) );
  AOI221_X1 U34469 ( .B1(n39574), .B2(n32506), .C1(n39568), .C2(n27946), .A(
        n34643), .ZN(n34636) );
  OAI222_X1 U34470 ( .A1(n30547), .A2(n39562), .B1(n30611), .B2(n39556), .C1(
        n30483), .C2(n39550), .ZN(n34643) );
  AOI221_X1 U34471 ( .B1(n39694), .B2(n29045), .C1(n39688), .C2(n29109), .A(
        n34635), .ZN(n34628) );
  OAI222_X1 U34472 ( .A1(n31433), .A2(n39682), .B1(n31497), .B2(n39676), .C1(
        n31369), .C2(n39670), .ZN(n34635) );
  AOI221_X1 U34473 ( .B1(n39322), .B2(n32506), .C1(n39316), .C2(n27946), .A(
        n35917), .ZN(n35910) );
  OAI222_X1 U34474 ( .A1(n30547), .A2(n39310), .B1(n30611), .B2(n39304), .C1(
        n30483), .C2(n39298), .ZN(n35917) );
  AOI221_X1 U34475 ( .B1(n39442), .B2(n29045), .C1(n39436), .C2(n29109), .A(
        n35909), .ZN(n35902) );
  OAI222_X1 U34476 ( .A1(n31433), .A2(n39430), .B1(n31497), .B2(n39424), .C1(
        n31369), .C2(n39418), .ZN(n35909) );
  AOI221_X1 U34477 ( .B1(n39574), .B2(n32509), .C1(n39568), .C2(n27945), .A(
        n34662), .ZN(n34655) );
  OAI222_X1 U34478 ( .A1(n30546), .A2(n39562), .B1(n30610), .B2(n39556), .C1(
        n30482), .C2(n39550), .ZN(n34662) );
  AOI221_X1 U34479 ( .B1(n39694), .B2(n29044), .C1(n39688), .C2(n29108), .A(
        n34654), .ZN(n34647) );
  OAI222_X1 U34480 ( .A1(n31432), .A2(n39682), .B1(n31496), .B2(n39676), .C1(
        n31368), .C2(n39670), .ZN(n34654) );
  AOI221_X1 U34481 ( .B1(n39322), .B2(n32509), .C1(n39316), .C2(n27945), .A(
        n35936), .ZN(n35929) );
  OAI222_X1 U34482 ( .A1(n30546), .A2(n39310), .B1(n30610), .B2(n39304), .C1(
        n30482), .C2(n39298), .ZN(n35936) );
  AOI221_X1 U34483 ( .B1(n39442), .B2(n29044), .C1(n39436), .C2(n29108), .A(
        n35928), .ZN(n35921) );
  OAI222_X1 U34484 ( .A1(n31432), .A2(n39430), .B1(n31496), .B2(n39424), .C1(
        n31368), .C2(n39418), .ZN(n35928) );
  AOI221_X1 U34485 ( .B1(n39574), .B2(n32508), .C1(n39568), .C2(n27944), .A(
        n34695), .ZN(n34685) );
  OAI222_X1 U34486 ( .A1(n30545), .A2(n39562), .B1(n30609), .B2(n39556), .C1(
        n30481), .C2(n39550), .ZN(n34695) );
  AOI221_X1 U34487 ( .B1(n39694), .B2(n29043), .C1(n39688), .C2(n29107), .A(
        n34683), .ZN(n34666) );
  OAI222_X1 U34488 ( .A1(n31431), .A2(n39682), .B1(n31495), .B2(n39676), .C1(
        n31367), .C2(n39670), .ZN(n34683) );
  AOI221_X1 U34489 ( .B1(n39322), .B2(n32508), .C1(n39316), .C2(n27944), .A(
        n35969), .ZN(n35959) );
  OAI222_X1 U34490 ( .A1(n30545), .A2(n39310), .B1(n30609), .B2(n39304), .C1(
        n30481), .C2(n39298), .ZN(n35969) );
  AOI221_X1 U34491 ( .B1(n39442), .B2(n29043), .C1(n39436), .C2(n29107), .A(
        n35957), .ZN(n35940) );
  OAI222_X1 U34492 ( .A1(n31431), .A2(n39430), .B1(n31495), .B2(n39424), .C1(
        n31367), .C2(n39418), .ZN(n35957) );
  OAI22_X1 U34493 ( .A1(n16938), .A2(n39295), .B1(n36078), .B2(n39293), .ZN(
        n7198) );
  NOR2_X1 U34494 ( .A1(n36079), .A2(n36080), .ZN(n36078) );
  NAND4_X1 U34495 ( .A1(n36081), .A2(n36082), .A3(n36083), .A4(n36084), .ZN(
        n36080) );
  NAND4_X1 U34496 ( .A1(n36089), .A2(n36090), .A3(n36091), .A4(n36092), .ZN(
        n36079) );
  OAI22_X1 U34497 ( .A1(n16939), .A2(n39294), .B1(n36059), .B2(n39293), .ZN(
        n7199) );
  NOR2_X1 U34498 ( .A1(n36060), .A2(n36061), .ZN(n36059) );
  NAND4_X1 U34499 ( .A1(n36062), .A2(n36063), .A3(n36064), .A4(n36065), .ZN(
        n36061) );
  NAND4_X1 U34500 ( .A1(n36070), .A2(n36071), .A3(n36072), .A4(n36073), .ZN(
        n36060) );
  OAI22_X1 U34501 ( .A1(n16940), .A2(n39296), .B1(n36040), .B2(n39293), .ZN(
        n7200) );
  NOR2_X1 U34502 ( .A1(n36041), .A2(n36042), .ZN(n36040) );
  NAND4_X1 U34503 ( .A1(n36043), .A2(n36044), .A3(n36045), .A4(n36046), .ZN(
        n36042) );
  NAND4_X1 U34504 ( .A1(n36051), .A2(n36052), .A3(n36053), .A4(n36054), .ZN(
        n36041) );
  OAI22_X1 U34505 ( .A1(n16941), .A2(n39295), .B1(n35980), .B2(n39293), .ZN(
        n7201) );
  NOR2_X1 U34506 ( .A1(n35982), .A2(n35983), .ZN(n35980) );
  NAND4_X1 U34507 ( .A1(n35984), .A2(n35985), .A3(n35986), .A4(n35987), .ZN(
        n35983) );
  NAND4_X1 U34508 ( .A1(n36012), .A2(n36013), .A3(n36014), .A4(n36015), .ZN(
        n35982) );
  OAI22_X1 U34509 ( .A1(n17069), .A2(n39801), .B1(n33425), .B2(n39795), .ZN(
        n7330) );
  NOR2_X1 U34510 ( .A1(n33427), .A2(n33428), .ZN(n33425) );
  NAND4_X1 U34511 ( .A1(n33429), .A2(n33430), .A3(n33431), .A4(n33432), .ZN(
        n33428) );
  NAND4_X1 U34512 ( .A1(n33457), .A2(n33458), .A3(n33459), .A4(n33460), .ZN(
        n33427) );
  OAI22_X1 U34513 ( .A1(n17005), .A2(n39549), .B1(n34699), .B2(n39543), .ZN(
        n7266) );
  NOR2_X1 U34514 ( .A1(n34701), .A2(n34702), .ZN(n34699) );
  NAND4_X1 U34515 ( .A1(n34703), .A2(n34704), .A3(n34705), .A4(n34706), .ZN(
        n34702) );
  NAND4_X1 U34516 ( .A1(n34731), .A2(n34732), .A3(n34733), .A4(n34734), .ZN(
        n34701) );
  OAI22_X1 U34517 ( .A1(n17068), .A2(n39801), .B1(n33485), .B2(n39795), .ZN(
        n7329) );
  NOR2_X1 U34518 ( .A1(n33486), .A2(n33487), .ZN(n33485) );
  NAND4_X1 U34519 ( .A1(n33488), .A2(n33489), .A3(n33490), .A4(n33491), .ZN(
        n33487) );
  NAND4_X1 U34520 ( .A1(n33496), .A2(n33497), .A3(n33498), .A4(n33499), .ZN(
        n33486) );
  OAI22_X1 U34521 ( .A1(n17004), .A2(n39549), .B1(n34759), .B2(n39543), .ZN(
        n7265) );
  NOR2_X1 U34522 ( .A1(n34760), .A2(n34761), .ZN(n34759) );
  NAND4_X1 U34523 ( .A1(n34762), .A2(n34763), .A3(n34764), .A4(n34765), .ZN(
        n34761) );
  NAND4_X1 U34524 ( .A1(n34770), .A2(n34771), .A3(n34772), .A4(n34773), .ZN(
        n34760) );
  OAI22_X1 U34525 ( .A1(n17067), .A2(n39801), .B1(n33504), .B2(n39795), .ZN(
        n7328) );
  NOR2_X1 U34526 ( .A1(n33505), .A2(n33506), .ZN(n33504) );
  NAND4_X1 U34527 ( .A1(n33507), .A2(n33508), .A3(n33509), .A4(n33510), .ZN(
        n33506) );
  NAND4_X1 U34528 ( .A1(n33515), .A2(n33516), .A3(n33517), .A4(n33518), .ZN(
        n33505) );
  OAI22_X1 U34529 ( .A1(n17003), .A2(n39549), .B1(n34778), .B2(n39543), .ZN(
        n7264) );
  NOR2_X1 U34530 ( .A1(n34779), .A2(n34780), .ZN(n34778) );
  NAND4_X1 U34531 ( .A1(n34781), .A2(n34782), .A3(n34783), .A4(n34784), .ZN(
        n34780) );
  NAND4_X1 U34532 ( .A1(n34789), .A2(n34790), .A3(n34791), .A4(n34792), .ZN(
        n34779) );
  OAI22_X1 U34533 ( .A1(n17066), .A2(n39801), .B1(n33523), .B2(n39795), .ZN(
        n7327) );
  NOR2_X1 U34534 ( .A1(n33524), .A2(n33525), .ZN(n33523) );
  NAND4_X1 U34535 ( .A1(n33526), .A2(n33527), .A3(n33528), .A4(n33529), .ZN(
        n33525) );
  NAND4_X1 U34536 ( .A1(n33534), .A2(n33535), .A3(n33536), .A4(n33537), .ZN(
        n33524) );
  OAI22_X1 U34537 ( .A1(n17002), .A2(n39549), .B1(n34797), .B2(n39543), .ZN(
        n7263) );
  NOR2_X1 U34538 ( .A1(n34798), .A2(n34799), .ZN(n34797) );
  NAND4_X1 U34539 ( .A1(n34800), .A2(n34801), .A3(n34802), .A4(n34803), .ZN(
        n34799) );
  NAND4_X1 U34540 ( .A1(n34808), .A2(n34809), .A3(n34810), .A4(n34811), .ZN(
        n34798) );
  XOR2_X1 U34541 ( .A(n2683), .B(n39047), .Z(n33297) );
  NAND2_X1 U34542 ( .A1(n32242), .A2(\add_146/carry[4] ), .ZN(n39047) );
  OAI22_X1 U34543 ( .A1(n16878), .A2(n39296), .B1(n37218), .B2(n39288), .ZN(
        n7138) );
  NOR2_X1 U34544 ( .A1(n37219), .A2(n37220), .ZN(n37218) );
  NAND4_X1 U34545 ( .A1(n37221), .A2(n37222), .A3(n37223), .A4(n37224), .ZN(
        n37220) );
  NAND4_X1 U34546 ( .A1(n37241), .A2(n37242), .A3(n37243), .A4(n37244), .ZN(
        n37219) );
  OAI22_X1 U34547 ( .A1(n16932), .A2(n39295), .B1(n36192), .B2(n39292), .ZN(
        n7192) );
  NOR2_X1 U34548 ( .A1(n36193), .A2(n36194), .ZN(n36192) );
  NAND4_X1 U34549 ( .A1(n36195), .A2(n36196), .A3(n36197), .A4(n36198), .ZN(
        n36194) );
  NAND4_X1 U34550 ( .A1(n36203), .A2(n36204), .A3(n36205), .A4(n36206), .ZN(
        n36193) );
  OAI22_X1 U34551 ( .A1(n16933), .A2(n39294), .B1(n36173), .B2(n39292), .ZN(
        n7193) );
  NOR2_X1 U34552 ( .A1(n36174), .A2(n36175), .ZN(n36173) );
  NAND4_X1 U34553 ( .A1(n36176), .A2(n36177), .A3(n36178), .A4(n36179), .ZN(
        n36175) );
  NAND4_X1 U34554 ( .A1(n36184), .A2(n36185), .A3(n36186), .A4(n36187), .ZN(
        n36174) );
  OAI22_X1 U34555 ( .A1(n16934), .A2(n39296), .B1(n36154), .B2(n39292), .ZN(
        n7194) );
  NOR2_X1 U34556 ( .A1(n36155), .A2(n36156), .ZN(n36154) );
  NAND4_X1 U34557 ( .A1(n36157), .A2(n36158), .A3(n36159), .A4(n36160), .ZN(
        n36156) );
  NAND4_X1 U34558 ( .A1(n36165), .A2(n36166), .A3(n36167), .A4(n36168), .ZN(
        n36155) );
  OAI22_X1 U34559 ( .A1(n16935), .A2(n39295), .B1(n36135), .B2(n39292), .ZN(
        n7195) );
  NOR2_X1 U34560 ( .A1(n36136), .A2(n36137), .ZN(n36135) );
  NAND4_X1 U34561 ( .A1(n36138), .A2(n36139), .A3(n36140), .A4(n36141), .ZN(
        n36137) );
  NAND4_X1 U34562 ( .A1(n36146), .A2(n36147), .A3(n36148), .A4(n36149), .ZN(
        n36136) );
  OAI22_X1 U34563 ( .A1(n16936), .A2(n39294), .B1(n36116), .B2(n39292), .ZN(
        n7196) );
  NOR2_X1 U34564 ( .A1(n36117), .A2(n36118), .ZN(n36116) );
  NAND4_X1 U34565 ( .A1(n36119), .A2(n36120), .A3(n36121), .A4(n36122), .ZN(
        n36118) );
  NAND4_X1 U34566 ( .A1(n36127), .A2(n36128), .A3(n36129), .A4(n36130), .ZN(
        n36117) );
  OAI22_X1 U34567 ( .A1(n16937), .A2(n39296), .B1(n36097), .B2(n39292), .ZN(
        n7197) );
  NOR2_X1 U34568 ( .A1(n36098), .A2(n36099), .ZN(n36097) );
  NAND4_X1 U34569 ( .A1(n36100), .A2(n36101), .A3(n36102), .A4(n36103), .ZN(
        n36099) );
  NAND4_X1 U34570 ( .A1(n36108), .A2(n36109), .A3(n36110), .A4(n36111), .ZN(
        n36098) );
  OAI22_X1 U34571 ( .A1(n16889), .A2(n39296), .B1(n37009), .B2(n39288), .ZN(
        n7149) );
  NOR2_X1 U34572 ( .A1(n37010), .A2(n37011), .ZN(n37009) );
  NAND4_X1 U34573 ( .A1(n37012), .A2(n37013), .A3(n37014), .A4(n37015), .ZN(
        n37011) );
  NAND4_X1 U34574 ( .A1(n37020), .A2(n37021), .A3(n37022), .A4(n37023), .ZN(
        n37010) );
  OAI22_X1 U34575 ( .A1(n16890), .A2(n39296), .B1(n36990), .B2(n39289), .ZN(
        n7150) );
  NOR2_X1 U34576 ( .A1(n36991), .A2(n36992), .ZN(n36990) );
  NAND4_X1 U34577 ( .A1(n36993), .A2(n36994), .A3(n36995), .A4(n36996), .ZN(
        n36992) );
  NAND4_X1 U34578 ( .A1(n37001), .A2(n37002), .A3(n37003), .A4(n37004), .ZN(
        n36991) );
  OAI22_X1 U34579 ( .A1(n16891), .A2(n39296), .B1(n36971), .B2(n39289), .ZN(
        n7151) );
  NOR2_X1 U34580 ( .A1(n36972), .A2(n36973), .ZN(n36971) );
  NAND4_X1 U34581 ( .A1(n36974), .A2(n36975), .A3(n36976), .A4(n36977), .ZN(
        n36973) );
  NAND4_X1 U34582 ( .A1(n36982), .A2(n36983), .A3(n36984), .A4(n36985), .ZN(
        n36972) );
  OAI22_X1 U34583 ( .A1(n16892), .A2(n39296), .B1(n36952), .B2(n39289), .ZN(
        n7152) );
  NOR2_X1 U34584 ( .A1(n36953), .A2(n36954), .ZN(n36952) );
  NAND4_X1 U34585 ( .A1(n36955), .A2(n36956), .A3(n36957), .A4(n36958), .ZN(
        n36954) );
  NAND4_X1 U34586 ( .A1(n36963), .A2(n36964), .A3(n36965), .A4(n36966), .ZN(
        n36953) );
  OAI22_X1 U34587 ( .A1(n16893), .A2(n39296), .B1(n36933), .B2(n39289), .ZN(
        n7153) );
  NOR2_X1 U34588 ( .A1(n36934), .A2(n36935), .ZN(n36933) );
  NAND4_X1 U34589 ( .A1(n36936), .A2(n36937), .A3(n36938), .A4(n36939), .ZN(
        n36935) );
  NAND4_X1 U34590 ( .A1(n36944), .A2(n36945), .A3(n36946), .A4(n36947), .ZN(
        n36934) );
  OAI22_X1 U34591 ( .A1(n16894), .A2(n39296), .B1(n36914), .B2(n39289), .ZN(
        n7154) );
  NOR2_X1 U34592 ( .A1(n36915), .A2(n36916), .ZN(n36914) );
  NAND4_X1 U34593 ( .A1(n36917), .A2(n36918), .A3(n36919), .A4(n36920), .ZN(
        n36916) );
  NAND4_X1 U34594 ( .A1(n36925), .A2(n36926), .A3(n36927), .A4(n36928), .ZN(
        n36915) );
  OAI22_X1 U34595 ( .A1(n16895), .A2(n39296), .B1(n36895), .B2(n39289), .ZN(
        n7155) );
  NOR2_X1 U34596 ( .A1(n36896), .A2(n36897), .ZN(n36895) );
  NAND4_X1 U34597 ( .A1(n36898), .A2(n36899), .A3(n36900), .A4(n36901), .ZN(
        n36897) );
  NAND4_X1 U34598 ( .A1(n36906), .A2(n36907), .A3(n36908), .A4(n36909), .ZN(
        n36896) );
  OAI22_X1 U34599 ( .A1(n16896), .A2(n39296), .B1(n36876), .B2(n39289), .ZN(
        n7156) );
  NOR2_X1 U34600 ( .A1(n36877), .A2(n36878), .ZN(n36876) );
  NAND4_X1 U34601 ( .A1(n36879), .A2(n36880), .A3(n36881), .A4(n36882), .ZN(
        n36878) );
  NAND4_X1 U34602 ( .A1(n36887), .A2(n36888), .A3(n36889), .A4(n36890), .ZN(
        n36877) );
  OAI22_X1 U34603 ( .A1(n16897), .A2(n39295), .B1(n36857), .B2(n39289), .ZN(
        n7157) );
  NOR2_X1 U34604 ( .A1(n36858), .A2(n36859), .ZN(n36857) );
  NAND4_X1 U34605 ( .A1(n36860), .A2(n36861), .A3(n36862), .A4(n36863), .ZN(
        n36859) );
  NAND4_X1 U34606 ( .A1(n36868), .A2(n36869), .A3(n36870), .A4(n36871), .ZN(
        n36858) );
  OAI22_X1 U34607 ( .A1(n16898), .A2(n39296), .B1(n36838), .B2(n39289), .ZN(
        n7158) );
  NOR2_X1 U34608 ( .A1(n36839), .A2(n36840), .ZN(n36838) );
  NAND4_X1 U34609 ( .A1(n36841), .A2(n36842), .A3(n36843), .A4(n36844), .ZN(
        n36840) );
  NAND4_X1 U34610 ( .A1(n36849), .A2(n36850), .A3(n36851), .A4(n36852), .ZN(
        n36839) );
  OAI22_X1 U34611 ( .A1(n16899), .A2(n39295), .B1(n36819), .B2(n39289), .ZN(
        n7159) );
  NOR2_X1 U34612 ( .A1(n36820), .A2(n36821), .ZN(n36819) );
  NAND4_X1 U34613 ( .A1(n36822), .A2(n36823), .A3(n36824), .A4(n36825), .ZN(
        n36821) );
  NAND4_X1 U34614 ( .A1(n36830), .A2(n36831), .A3(n36832), .A4(n36833), .ZN(
        n36820) );
  OAI22_X1 U34615 ( .A1(n16900), .A2(n39296), .B1(n36800), .B2(n39289), .ZN(
        n7160) );
  NOR2_X1 U34616 ( .A1(n36801), .A2(n36802), .ZN(n36800) );
  NAND4_X1 U34617 ( .A1(n36803), .A2(n36804), .A3(n36805), .A4(n36806), .ZN(
        n36802) );
  NAND4_X1 U34618 ( .A1(n36811), .A2(n36812), .A3(n36813), .A4(n36814), .ZN(
        n36801) );
  OAI22_X1 U34619 ( .A1(n16901), .A2(n39295), .B1(n36781), .B2(n39289), .ZN(
        n7161) );
  NOR2_X1 U34620 ( .A1(n36782), .A2(n36783), .ZN(n36781) );
  NAND4_X1 U34621 ( .A1(n36784), .A2(n36785), .A3(n36786), .A4(n36787), .ZN(
        n36783) );
  NAND4_X1 U34622 ( .A1(n36792), .A2(n36793), .A3(n36794), .A4(n36795), .ZN(
        n36782) );
  OAI22_X1 U34623 ( .A1(n16902), .A2(n39296), .B1(n36762), .B2(n39290), .ZN(
        n7162) );
  NOR2_X1 U34624 ( .A1(n36763), .A2(n36764), .ZN(n36762) );
  NAND4_X1 U34625 ( .A1(n36765), .A2(n36766), .A3(n36767), .A4(n36768), .ZN(
        n36764) );
  NAND4_X1 U34626 ( .A1(n36773), .A2(n36774), .A3(n36775), .A4(n36776), .ZN(
        n36763) );
  OAI22_X1 U34627 ( .A1(n16903), .A2(n39295), .B1(n36743), .B2(n39290), .ZN(
        n7163) );
  NOR2_X1 U34628 ( .A1(n36744), .A2(n36745), .ZN(n36743) );
  NAND4_X1 U34629 ( .A1(n36746), .A2(n36747), .A3(n36748), .A4(n36749), .ZN(
        n36745) );
  NAND4_X1 U34630 ( .A1(n36754), .A2(n36755), .A3(n36756), .A4(n36757), .ZN(
        n36744) );
  OAI22_X1 U34631 ( .A1(n16904), .A2(n39296), .B1(n36724), .B2(n39290), .ZN(
        n7164) );
  NOR2_X1 U34632 ( .A1(n36725), .A2(n36726), .ZN(n36724) );
  NAND4_X1 U34633 ( .A1(n36727), .A2(n36728), .A3(n36729), .A4(n36730), .ZN(
        n36726) );
  NAND4_X1 U34634 ( .A1(n36735), .A2(n36736), .A3(n36737), .A4(n36738), .ZN(
        n36725) );
  OAI22_X1 U34635 ( .A1(n16905), .A2(n39295), .B1(n36705), .B2(n39290), .ZN(
        n7165) );
  NOR2_X1 U34636 ( .A1(n36706), .A2(n36707), .ZN(n36705) );
  NAND4_X1 U34637 ( .A1(n36708), .A2(n36709), .A3(n36710), .A4(n36711), .ZN(
        n36707) );
  NAND4_X1 U34638 ( .A1(n36716), .A2(n36717), .A3(n36718), .A4(n36719), .ZN(
        n36706) );
  OAI22_X1 U34639 ( .A1(n16906), .A2(n39296), .B1(n36686), .B2(n39290), .ZN(
        n7166) );
  NOR2_X1 U34640 ( .A1(n36687), .A2(n36688), .ZN(n36686) );
  NAND4_X1 U34641 ( .A1(n36689), .A2(n36690), .A3(n36691), .A4(n36692), .ZN(
        n36688) );
  NAND4_X1 U34642 ( .A1(n36697), .A2(n36698), .A3(n36699), .A4(n36700), .ZN(
        n36687) );
  OAI22_X1 U34643 ( .A1(n16907), .A2(n39295), .B1(n36667), .B2(n39290), .ZN(
        n7167) );
  NOR2_X1 U34644 ( .A1(n36668), .A2(n36669), .ZN(n36667) );
  NAND4_X1 U34645 ( .A1(n36670), .A2(n36671), .A3(n36672), .A4(n36673), .ZN(
        n36669) );
  NAND4_X1 U34646 ( .A1(n36678), .A2(n36679), .A3(n36680), .A4(n36681), .ZN(
        n36668) );
  OAI22_X1 U34647 ( .A1(n16908), .A2(n39295), .B1(n36648), .B2(n39290), .ZN(
        n7168) );
  NOR2_X1 U34648 ( .A1(n36649), .A2(n36650), .ZN(n36648) );
  NAND4_X1 U34649 ( .A1(n36651), .A2(n36652), .A3(n36653), .A4(n36654), .ZN(
        n36650) );
  NAND4_X1 U34650 ( .A1(n36659), .A2(n36660), .A3(n36661), .A4(n36662), .ZN(
        n36649) );
  OAI22_X1 U34651 ( .A1(n16909), .A2(n39295), .B1(n36629), .B2(n39290), .ZN(
        n7169) );
  NOR2_X1 U34652 ( .A1(n36630), .A2(n36631), .ZN(n36629) );
  NAND4_X1 U34653 ( .A1(n36632), .A2(n36633), .A3(n36634), .A4(n36635), .ZN(
        n36631) );
  NAND4_X1 U34654 ( .A1(n36640), .A2(n36641), .A3(n36642), .A4(n36643), .ZN(
        n36630) );
  OAI22_X1 U34655 ( .A1(n16910), .A2(n39295), .B1(n36610), .B2(n39290), .ZN(
        n7170) );
  NOR2_X1 U34656 ( .A1(n36611), .A2(n36612), .ZN(n36610) );
  NAND4_X1 U34657 ( .A1(n36613), .A2(n36614), .A3(n36615), .A4(n36616), .ZN(
        n36612) );
  NAND4_X1 U34658 ( .A1(n36621), .A2(n36622), .A3(n36623), .A4(n36624), .ZN(
        n36611) );
  OAI22_X1 U34659 ( .A1(n16911), .A2(n39295), .B1(n36591), .B2(n39290), .ZN(
        n7171) );
  NOR2_X1 U34660 ( .A1(n36592), .A2(n36593), .ZN(n36591) );
  NAND4_X1 U34661 ( .A1(n36594), .A2(n36595), .A3(n36596), .A4(n36597), .ZN(
        n36593) );
  NAND4_X1 U34662 ( .A1(n36602), .A2(n36603), .A3(n36604), .A4(n36605), .ZN(
        n36592) );
  OAI22_X1 U34663 ( .A1(n16912), .A2(n39295), .B1(n36572), .B2(n39290), .ZN(
        n7172) );
  NOR2_X1 U34664 ( .A1(n36573), .A2(n36574), .ZN(n36572) );
  NAND4_X1 U34665 ( .A1(n36575), .A2(n36576), .A3(n36577), .A4(n36578), .ZN(
        n36574) );
  NAND4_X1 U34666 ( .A1(n36583), .A2(n36584), .A3(n36585), .A4(n36586), .ZN(
        n36573) );
  OAI22_X1 U34667 ( .A1(n16913), .A2(n39295), .B1(n36553), .B2(n39290), .ZN(
        n7173) );
  NOR2_X1 U34668 ( .A1(n36554), .A2(n36555), .ZN(n36553) );
  NAND4_X1 U34669 ( .A1(n36556), .A2(n36557), .A3(n36558), .A4(n36559), .ZN(
        n36555) );
  NAND4_X1 U34670 ( .A1(n36564), .A2(n36565), .A3(n36566), .A4(n36567), .ZN(
        n36554) );
  OAI22_X1 U34671 ( .A1(n16914), .A2(n39295), .B1(n36534), .B2(n39291), .ZN(
        n7174) );
  NOR2_X1 U34672 ( .A1(n36535), .A2(n36536), .ZN(n36534) );
  NAND4_X1 U34673 ( .A1(n36537), .A2(n36538), .A3(n36539), .A4(n36540), .ZN(
        n36536) );
  NAND4_X1 U34674 ( .A1(n36545), .A2(n36546), .A3(n36547), .A4(n36548), .ZN(
        n36535) );
  OAI22_X1 U34675 ( .A1(n16915), .A2(n39295), .B1(n36515), .B2(n39291), .ZN(
        n7175) );
  NOR2_X1 U34676 ( .A1(n36516), .A2(n36517), .ZN(n36515) );
  NAND4_X1 U34677 ( .A1(n36518), .A2(n36519), .A3(n36520), .A4(n36521), .ZN(
        n36517) );
  NAND4_X1 U34678 ( .A1(n36526), .A2(n36527), .A3(n36528), .A4(n36529), .ZN(
        n36516) );
  OAI22_X1 U34679 ( .A1(n16916), .A2(n39295), .B1(n36496), .B2(n39291), .ZN(
        n7176) );
  NOR2_X1 U34680 ( .A1(n36497), .A2(n36498), .ZN(n36496) );
  NAND4_X1 U34681 ( .A1(n36499), .A2(n36500), .A3(n36501), .A4(n36502), .ZN(
        n36498) );
  NAND4_X1 U34682 ( .A1(n36507), .A2(n36508), .A3(n36509), .A4(n36510), .ZN(
        n36497) );
  OAI22_X1 U34683 ( .A1(n16917), .A2(n39295), .B1(n36477), .B2(n39291), .ZN(
        n7177) );
  NOR2_X1 U34684 ( .A1(n36478), .A2(n36479), .ZN(n36477) );
  NAND4_X1 U34685 ( .A1(n36480), .A2(n36481), .A3(n36482), .A4(n36483), .ZN(
        n36479) );
  NAND4_X1 U34686 ( .A1(n36488), .A2(n36489), .A3(n36490), .A4(n36491), .ZN(
        n36478) );
  OAI22_X1 U34687 ( .A1(n16918), .A2(n39295), .B1(n36458), .B2(n39291), .ZN(
        n7178) );
  NOR2_X1 U34688 ( .A1(n36459), .A2(n36460), .ZN(n36458) );
  NAND4_X1 U34689 ( .A1(n36461), .A2(n36462), .A3(n36463), .A4(n36464), .ZN(
        n36460) );
  NAND4_X1 U34690 ( .A1(n36469), .A2(n36470), .A3(n36471), .A4(n36472), .ZN(
        n36459) );
  OAI22_X1 U34691 ( .A1(n16919), .A2(n39294), .B1(n36439), .B2(n39291), .ZN(
        n7179) );
  NOR2_X1 U34692 ( .A1(n36440), .A2(n36441), .ZN(n36439) );
  NAND4_X1 U34693 ( .A1(n36442), .A2(n36443), .A3(n36444), .A4(n36445), .ZN(
        n36441) );
  NAND4_X1 U34694 ( .A1(n36450), .A2(n36451), .A3(n36452), .A4(n36453), .ZN(
        n36440) );
  OAI22_X1 U34695 ( .A1(n16920), .A2(n39294), .B1(n36420), .B2(n39291), .ZN(
        n7180) );
  NOR2_X1 U34696 ( .A1(n36421), .A2(n36422), .ZN(n36420) );
  NAND4_X1 U34697 ( .A1(n36423), .A2(n36424), .A3(n36425), .A4(n36426), .ZN(
        n36422) );
  NAND4_X1 U34698 ( .A1(n36431), .A2(n36432), .A3(n36433), .A4(n36434), .ZN(
        n36421) );
  OAI22_X1 U34699 ( .A1(n16921), .A2(n39294), .B1(n36401), .B2(n39291), .ZN(
        n7181) );
  NOR2_X1 U34700 ( .A1(n36402), .A2(n36403), .ZN(n36401) );
  NAND4_X1 U34701 ( .A1(n36404), .A2(n36405), .A3(n36406), .A4(n36407), .ZN(
        n36403) );
  NAND4_X1 U34702 ( .A1(n36412), .A2(n36413), .A3(n36414), .A4(n36415), .ZN(
        n36402) );
  OAI22_X1 U34703 ( .A1(n16922), .A2(n39294), .B1(n36382), .B2(n39291), .ZN(
        n7182) );
  NOR2_X1 U34704 ( .A1(n36383), .A2(n36384), .ZN(n36382) );
  NAND4_X1 U34705 ( .A1(n36385), .A2(n36386), .A3(n36387), .A4(n36388), .ZN(
        n36384) );
  NAND4_X1 U34706 ( .A1(n36393), .A2(n36394), .A3(n36395), .A4(n36396), .ZN(
        n36383) );
  OAI22_X1 U34707 ( .A1(n16923), .A2(n39294), .B1(n36363), .B2(n39291), .ZN(
        n7183) );
  NOR2_X1 U34708 ( .A1(n36364), .A2(n36365), .ZN(n36363) );
  NAND4_X1 U34709 ( .A1(n36366), .A2(n36367), .A3(n36368), .A4(n36369), .ZN(
        n36365) );
  NAND4_X1 U34710 ( .A1(n36374), .A2(n36375), .A3(n36376), .A4(n36377), .ZN(
        n36364) );
  OAI22_X1 U34711 ( .A1(n16924), .A2(n39294), .B1(n36344), .B2(n39291), .ZN(
        n7184) );
  NOR2_X1 U34712 ( .A1(n36345), .A2(n36346), .ZN(n36344) );
  NAND4_X1 U34713 ( .A1(n36347), .A2(n36348), .A3(n36349), .A4(n36350), .ZN(
        n36346) );
  NAND4_X1 U34714 ( .A1(n36355), .A2(n36356), .A3(n36357), .A4(n36358), .ZN(
        n36345) );
  OAI22_X1 U34715 ( .A1(n16925), .A2(n39294), .B1(n36325), .B2(n39291), .ZN(
        n7185) );
  NOR2_X1 U34716 ( .A1(n36326), .A2(n36327), .ZN(n36325) );
  NAND4_X1 U34717 ( .A1(n36328), .A2(n36329), .A3(n36330), .A4(n36331), .ZN(
        n36327) );
  NAND4_X1 U34718 ( .A1(n36336), .A2(n36337), .A3(n36338), .A4(n36339), .ZN(
        n36326) );
  OAI22_X1 U34719 ( .A1(n16926), .A2(n39294), .B1(n36306), .B2(n39292), .ZN(
        n7186) );
  NOR2_X1 U34720 ( .A1(n36307), .A2(n36308), .ZN(n36306) );
  NAND4_X1 U34721 ( .A1(n36309), .A2(n36310), .A3(n36311), .A4(n36312), .ZN(
        n36308) );
  NAND4_X1 U34722 ( .A1(n36317), .A2(n36318), .A3(n36319), .A4(n36320), .ZN(
        n36307) );
  OAI22_X1 U34723 ( .A1(n16927), .A2(n39295), .B1(n36287), .B2(n39292), .ZN(
        n7187) );
  NOR2_X1 U34724 ( .A1(n36288), .A2(n36289), .ZN(n36287) );
  NAND4_X1 U34725 ( .A1(n36290), .A2(n36291), .A3(n36292), .A4(n36293), .ZN(
        n36289) );
  NAND4_X1 U34726 ( .A1(n36298), .A2(n36299), .A3(n36300), .A4(n36301), .ZN(
        n36288) );
  OAI22_X1 U34727 ( .A1(n16928), .A2(n39294), .B1(n36268), .B2(n39292), .ZN(
        n7188) );
  NOR2_X1 U34728 ( .A1(n36269), .A2(n36270), .ZN(n36268) );
  NAND4_X1 U34729 ( .A1(n36271), .A2(n36272), .A3(n36273), .A4(n36274), .ZN(
        n36270) );
  NAND4_X1 U34730 ( .A1(n36279), .A2(n36280), .A3(n36281), .A4(n36282), .ZN(
        n36269) );
  OAI22_X1 U34731 ( .A1(n16929), .A2(n39294), .B1(n36249), .B2(n39292), .ZN(
        n7189) );
  NOR2_X1 U34732 ( .A1(n36250), .A2(n36251), .ZN(n36249) );
  NAND4_X1 U34733 ( .A1(n36252), .A2(n36253), .A3(n36254), .A4(n36255), .ZN(
        n36251) );
  NAND4_X1 U34734 ( .A1(n36260), .A2(n36261), .A3(n36262), .A4(n36263), .ZN(
        n36250) );
  OAI22_X1 U34735 ( .A1(n16930), .A2(n39294), .B1(n36230), .B2(n39292), .ZN(
        n7190) );
  NOR2_X1 U34736 ( .A1(n36231), .A2(n36232), .ZN(n36230) );
  NAND4_X1 U34737 ( .A1(n36233), .A2(n36234), .A3(n36235), .A4(n36236), .ZN(
        n36232) );
  NAND4_X1 U34738 ( .A1(n36241), .A2(n36242), .A3(n36243), .A4(n36244), .ZN(
        n36231) );
  OAI22_X1 U34739 ( .A1(n16931), .A2(n39294), .B1(n36211), .B2(n39292), .ZN(
        n7191) );
  NOR2_X1 U34740 ( .A1(n36212), .A2(n36213), .ZN(n36211) );
  NAND4_X1 U34741 ( .A1(n36214), .A2(n36215), .A3(n36216), .A4(n36217), .ZN(
        n36213) );
  NAND4_X1 U34742 ( .A1(n36222), .A2(n36223), .A3(n36224), .A4(n36225), .ZN(
        n36212) );
  OAI22_X1 U34743 ( .A1(n16879), .A2(n39295), .B1(n37199), .B2(n39288), .ZN(
        n7139) );
  NOR2_X1 U34744 ( .A1(n37200), .A2(n37201), .ZN(n37199) );
  NAND4_X1 U34745 ( .A1(n37202), .A2(n37203), .A3(n37204), .A4(n37205), .ZN(
        n37201) );
  NAND4_X1 U34746 ( .A1(n37210), .A2(n37211), .A3(n37212), .A4(n37213), .ZN(
        n37200) );
  OAI22_X1 U34747 ( .A1(n16880), .A2(n39294), .B1(n37180), .B2(n39288), .ZN(
        n7140) );
  NOR2_X1 U34748 ( .A1(n37181), .A2(n37182), .ZN(n37180) );
  NAND4_X1 U34749 ( .A1(n37183), .A2(n37184), .A3(n37185), .A4(n37186), .ZN(
        n37182) );
  NAND4_X1 U34750 ( .A1(n37191), .A2(n37192), .A3(n37193), .A4(n37194), .ZN(
        n37181) );
  OAI22_X1 U34751 ( .A1(n16881), .A2(n39296), .B1(n37161), .B2(n39288), .ZN(
        n7141) );
  NOR2_X1 U34752 ( .A1(n37162), .A2(n37163), .ZN(n37161) );
  NAND4_X1 U34753 ( .A1(n37164), .A2(n37165), .A3(n37166), .A4(n37167), .ZN(
        n37163) );
  NAND4_X1 U34754 ( .A1(n37172), .A2(n37173), .A3(n37174), .A4(n37175), .ZN(
        n37162) );
  OAI22_X1 U34755 ( .A1(n16882), .A2(n39295), .B1(n37142), .B2(n39288), .ZN(
        n7142) );
  NOR2_X1 U34756 ( .A1(n37143), .A2(n37144), .ZN(n37142) );
  NAND4_X1 U34757 ( .A1(n37145), .A2(n37146), .A3(n37147), .A4(n37148), .ZN(
        n37144) );
  NAND4_X1 U34758 ( .A1(n37153), .A2(n37154), .A3(n37155), .A4(n37156), .ZN(
        n37143) );
  OAI22_X1 U34759 ( .A1(n16883), .A2(n39294), .B1(n37123), .B2(n39288), .ZN(
        n7143) );
  NOR2_X1 U34760 ( .A1(n37124), .A2(n37125), .ZN(n37123) );
  NAND4_X1 U34761 ( .A1(n37126), .A2(n37127), .A3(n37128), .A4(n37129), .ZN(
        n37125) );
  NAND4_X1 U34762 ( .A1(n37134), .A2(n37135), .A3(n37136), .A4(n37137), .ZN(
        n37124) );
  OAI22_X1 U34763 ( .A1(n16884), .A2(n39296), .B1(n37104), .B2(n39288), .ZN(
        n7144) );
  NOR2_X1 U34764 ( .A1(n37105), .A2(n37106), .ZN(n37104) );
  NAND4_X1 U34765 ( .A1(n37107), .A2(n37108), .A3(n37109), .A4(n37110), .ZN(
        n37106) );
  NAND4_X1 U34766 ( .A1(n37115), .A2(n37116), .A3(n37117), .A4(n37118), .ZN(
        n37105) );
  OAI22_X1 U34767 ( .A1(n16885), .A2(n39296), .B1(n37085), .B2(n39288), .ZN(
        n7145) );
  NOR2_X1 U34768 ( .A1(n37086), .A2(n37087), .ZN(n37085) );
  NAND4_X1 U34769 ( .A1(n37088), .A2(n37089), .A3(n37090), .A4(n37091), .ZN(
        n37087) );
  NAND4_X1 U34770 ( .A1(n37096), .A2(n37097), .A3(n37098), .A4(n37099), .ZN(
        n37086) );
  OAI22_X1 U34771 ( .A1(n16886), .A2(n39296), .B1(n37066), .B2(n39288), .ZN(
        n7146) );
  NOR2_X1 U34772 ( .A1(n37067), .A2(n37068), .ZN(n37066) );
  NAND4_X1 U34773 ( .A1(n37069), .A2(n37070), .A3(n37071), .A4(n37072), .ZN(
        n37068) );
  NAND4_X1 U34774 ( .A1(n37077), .A2(n37078), .A3(n37079), .A4(n37080), .ZN(
        n37067) );
  OAI22_X1 U34775 ( .A1(n16887), .A2(n39296), .B1(n37047), .B2(n39288), .ZN(
        n7147) );
  NOR2_X1 U34776 ( .A1(n37048), .A2(n37049), .ZN(n37047) );
  NAND4_X1 U34777 ( .A1(n37050), .A2(n37051), .A3(n37052), .A4(n37053), .ZN(
        n37049) );
  NAND4_X1 U34778 ( .A1(n37058), .A2(n37059), .A3(n37060), .A4(n37061), .ZN(
        n37048) );
  OAI22_X1 U34779 ( .A1(n16888), .A2(n39296), .B1(n37028), .B2(n39288), .ZN(
        n7148) );
  NOR2_X1 U34780 ( .A1(n37029), .A2(n37030), .ZN(n37028) );
  NAND4_X1 U34781 ( .A1(n37031), .A2(n37032), .A3(n37033), .A4(n37034), .ZN(
        n37030) );
  NAND4_X1 U34782 ( .A1(n37039), .A2(n37040), .A3(n37041), .A4(n37042), .ZN(
        n37029) );
  OAI22_X1 U34783 ( .A1(n17065), .A2(n39801), .B1(n33542), .B2(n39794), .ZN(
        n7326) );
  NOR2_X1 U34784 ( .A1(n33543), .A2(n33544), .ZN(n33542) );
  NAND4_X1 U34785 ( .A1(n33545), .A2(n33546), .A3(n33547), .A4(n33548), .ZN(
        n33544) );
  NAND4_X1 U34786 ( .A1(n33553), .A2(n33554), .A3(n33555), .A4(n33556), .ZN(
        n33543) );
  OAI22_X1 U34787 ( .A1(n17001), .A2(n39549), .B1(n34816), .B2(n39542), .ZN(
        n7262) );
  NOR2_X1 U34788 ( .A1(n34817), .A2(n34818), .ZN(n34816) );
  NAND4_X1 U34789 ( .A1(n34819), .A2(n34820), .A3(n34821), .A4(n34822), .ZN(
        n34818) );
  NAND4_X1 U34790 ( .A1(n34827), .A2(n34828), .A3(n34829), .A4(n34830), .ZN(
        n34817) );
  OAI22_X1 U34791 ( .A1(n17064), .A2(n39800), .B1(n33561), .B2(n39794), .ZN(
        n7325) );
  NOR2_X1 U34792 ( .A1(n33562), .A2(n33563), .ZN(n33561) );
  NAND4_X1 U34793 ( .A1(n33564), .A2(n33565), .A3(n33566), .A4(n33567), .ZN(
        n33563) );
  NAND4_X1 U34794 ( .A1(n33572), .A2(n33573), .A3(n33574), .A4(n33575), .ZN(
        n33562) );
  OAI22_X1 U34795 ( .A1(n17000), .A2(n39548), .B1(n34835), .B2(n39542), .ZN(
        n7261) );
  NOR2_X1 U34796 ( .A1(n34836), .A2(n34837), .ZN(n34835) );
  NAND4_X1 U34797 ( .A1(n34838), .A2(n34839), .A3(n34840), .A4(n34841), .ZN(
        n34837) );
  NAND4_X1 U34798 ( .A1(n34846), .A2(n34847), .A3(n34848), .A4(n34849), .ZN(
        n34836) );
  OAI22_X1 U34799 ( .A1(n17063), .A2(n39800), .B1(n33580), .B2(n39794), .ZN(
        n7324) );
  NOR2_X1 U34800 ( .A1(n33581), .A2(n33582), .ZN(n33580) );
  NAND4_X1 U34801 ( .A1(n33583), .A2(n33584), .A3(n33585), .A4(n33586), .ZN(
        n33582) );
  NAND4_X1 U34802 ( .A1(n33591), .A2(n33592), .A3(n33593), .A4(n33594), .ZN(
        n33581) );
  OAI22_X1 U34803 ( .A1(n16999), .A2(n39548), .B1(n34854), .B2(n39542), .ZN(
        n7260) );
  NOR2_X1 U34804 ( .A1(n34855), .A2(n34856), .ZN(n34854) );
  NAND4_X1 U34805 ( .A1(n34857), .A2(n34858), .A3(n34859), .A4(n34860), .ZN(
        n34856) );
  NAND4_X1 U34806 ( .A1(n34865), .A2(n34866), .A3(n34867), .A4(n34868), .ZN(
        n34855) );
  OAI22_X1 U34807 ( .A1(n17062), .A2(n39800), .B1(n33599), .B2(n39794), .ZN(
        n7323) );
  NOR2_X1 U34808 ( .A1(n33600), .A2(n33601), .ZN(n33599) );
  NAND4_X1 U34809 ( .A1(n33602), .A2(n33603), .A3(n33604), .A4(n33605), .ZN(
        n33601) );
  NAND4_X1 U34810 ( .A1(n33610), .A2(n33611), .A3(n33612), .A4(n33613), .ZN(
        n33600) );
  OAI22_X1 U34811 ( .A1(n16998), .A2(n39548), .B1(n34873), .B2(n39542), .ZN(
        n7259) );
  NOR2_X1 U34812 ( .A1(n34874), .A2(n34875), .ZN(n34873) );
  NAND4_X1 U34813 ( .A1(n34876), .A2(n34877), .A3(n34878), .A4(n34879), .ZN(
        n34875) );
  NAND4_X1 U34814 ( .A1(n34884), .A2(n34885), .A3(n34886), .A4(n34887), .ZN(
        n34874) );
  OAI22_X1 U34815 ( .A1(n17061), .A2(n39800), .B1(n33618), .B2(n39794), .ZN(
        n7322) );
  NOR2_X1 U34816 ( .A1(n33619), .A2(n33620), .ZN(n33618) );
  NAND4_X1 U34817 ( .A1(n33621), .A2(n33622), .A3(n33623), .A4(n33624), .ZN(
        n33620) );
  NAND4_X1 U34818 ( .A1(n33629), .A2(n33630), .A3(n33631), .A4(n33632), .ZN(
        n33619) );
  OAI22_X1 U34819 ( .A1(n16997), .A2(n39548), .B1(n34892), .B2(n39542), .ZN(
        n7258) );
  NOR2_X1 U34820 ( .A1(n34893), .A2(n34894), .ZN(n34892) );
  NAND4_X1 U34821 ( .A1(n34895), .A2(n34896), .A3(n34897), .A4(n34898), .ZN(
        n34894) );
  NAND4_X1 U34822 ( .A1(n34903), .A2(n34904), .A3(n34905), .A4(n34906), .ZN(
        n34893) );
  OAI22_X1 U34823 ( .A1(n17060), .A2(n39800), .B1(n33637), .B2(n39794), .ZN(
        n7321) );
  NOR2_X1 U34824 ( .A1(n33638), .A2(n33639), .ZN(n33637) );
  NAND4_X1 U34825 ( .A1(n33640), .A2(n33641), .A3(n33642), .A4(n33643), .ZN(
        n33639) );
  NAND4_X1 U34826 ( .A1(n33648), .A2(n33649), .A3(n33650), .A4(n33651), .ZN(
        n33638) );
  OAI22_X1 U34827 ( .A1(n16996), .A2(n39548), .B1(n34911), .B2(n39542), .ZN(
        n7257) );
  NOR2_X1 U34828 ( .A1(n34912), .A2(n34913), .ZN(n34911) );
  NAND4_X1 U34829 ( .A1(n34914), .A2(n34915), .A3(n34916), .A4(n34917), .ZN(
        n34913) );
  NAND4_X1 U34830 ( .A1(n34922), .A2(n34923), .A3(n34924), .A4(n34925), .ZN(
        n34912) );
  OAI22_X1 U34831 ( .A1(n17059), .A2(n39800), .B1(n33656), .B2(n39794), .ZN(
        n7320) );
  NOR2_X1 U34832 ( .A1(n33657), .A2(n33658), .ZN(n33656) );
  NAND4_X1 U34833 ( .A1(n33659), .A2(n33660), .A3(n33661), .A4(n33662), .ZN(
        n33658) );
  NAND4_X1 U34834 ( .A1(n33667), .A2(n33668), .A3(n33669), .A4(n33670), .ZN(
        n33657) );
  OAI22_X1 U34835 ( .A1(n16995), .A2(n39548), .B1(n34930), .B2(n39542), .ZN(
        n7256) );
  NOR2_X1 U34836 ( .A1(n34931), .A2(n34932), .ZN(n34930) );
  NAND4_X1 U34837 ( .A1(n34933), .A2(n34934), .A3(n34935), .A4(n34936), .ZN(
        n34932) );
  NAND4_X1 U34838 ( .A1(n34941), .A2(n34942), .A3(n34943), .A4(n34944), .ZN(
        n34931) );
  OAI22_X1 U34839 ( .A1(n17058), .A2(n39800), .B1(n33675), .B2(n39794), .ZN(
        n7319) );
  NOR2_X1 U34840 ( .A1(n33676), .A2(n33677), .ZN(n33675) );
  NAND4_X1 U34841 ( .A1(n33678), .A2(n33679), .A3(n33680), .A4(n33681), .ZN(
        n33677) );
  NAND4_X1 U34842 ( .A1(n33686), .A2(n33687), .A3(n33688), .A4(n33689), .ZN(
        n33676) );
  OAI22_X1 U34843 ( .A1(n16994), .A2(n39548), .B1(n34949), .B2(n39542), .ZN(
        n7255) );
  NOR2_X1 U34844 ( .A1(n34950), .A2(n34951), .ZN(n34949) );
  NAND4_X1 U34845 ( .A1(n34952), .A2(n34953), .A3(n34954), .A4(n34955), .ZN(
        n34951) );
  NAND4_X1 U34846 ( .A1(n34960), .A2(n34961), .A3(n34962), .A4(n34963), .ZN(
        n34950) );
  OAI22_X1 U34847 ( .A1(n17057), .A2(n39800), .B1(n33694), .B2(n39794), .ZN(
        n7318) );
  NOR2_X1 U34848 ( .A1(n33695), .A2(n33696), .ZN(n33694) );
  NAND4_X1 U34849 ( .A1(n33697), .A2(n33698), .A3(n33699), .A4(n33700), .ZN(
        n33696) );
  NAND4_X1 U34850 ( .A1(n33705), .A2(n33706), .A3(n33707), .A4(n33708), .ZN(
        n33695) );
  OAI22_X1 U34851 ( .A1(n16993), .A2(n39548), .B1(n34968), .B2(n39542), .ZN(
        n7254) );
  NOR2_X1 U34852 ( .A1(n34969), .A2(n34970), .ZN(n34968) );
  NAND4_X1 U34853 ( .A1(n34971), .A2(n34972), .A3(n34973), .A4(n34974), .ZN(
        n34970) );
  NAND4_X1 U34854 ( .A1(n34979), .A2(n34980), .A3(n34981), .A4(n34982), .ZN(
        n34969) );
  OAI22_X1 U34855 ( .A1(n17056), .A2(n39800), .B1(n33713), .B2(n39794), .ZN(
        n7317) );
  NOR2_X1 U34856 ( .A1(n33714), .A2(n33715), .ZN(n33713) );
  NAND4_X1 U34857 ( .A1(n33716), .A2(n33717), .A3(n33718), .A4(n33719), .ZN(
        n33715) );
  NAND4_X1 U34858 ( .A1(n33724), .A2(n33725), .A3(n33726), .A4(n33727), .ZN(
        n33714) );
  OAI22_X1 U34859 ( .A1(n16992), .A2(n39548), .B1(n34987), .B2(n39542), .ZN(
        n7253) );
  NOR2_X1 U34860 ( .A1(n34988), .A2(n34989), .ZN(n34987) );
  NAND4_X1 U34861 ( .A1(n34990), .A2(n34991), .A3(n34992), .A4(n34993), .ZN(
        n34989) );
  NAND4_X1 U34862 ( .A1(n34998), .A2(n34999), .A3(n35000), .A4(n35001), .ZN(
        n34988) );
  OAI22_X1 U34863 ( .A1(n17055), .A2(n39800), .B1(n33732), .B2(n39794), .ZN(
        n7316) );
  NOR2_X1 U34864 ( .A1(n33733), .A2(n33734), .ZN(n33732) );
  NAND4_X1 U34865 ( .A1(n33735), .A2(n33736), .A3(n33737), .A4(n33738), .ZN(
        n33734) );
  NAND4_X1 U34866 ( .A1(n33743), .A2(n33744), .A3(n33745), .A4(n33746), .ZN(
        n33733) );
  OAI22_X1 U34867 ( .A1(n16991), .A2(n39548), .B1(n35006), .B2(n39542), .ZN(
        n7252) );
  NOR2_X1 U34868 ( .A1(n35007), .A2(n35008), .ZN(n35006) );
  NAND4_X1 U34869 ( .A1(n35009), .A2(n35010), .A3(n35011), .A4(n35012), .ZN(
        n35008) );
  NAND4_X1 U34870 ( .A1(n35017), .A2(n35018), .A3(n35019), .A4(n35020), .ZN(
        n35007) );
  OAI22_X1 U34871 ( .A1(n17054), .A2(n39800), .B1(n33751), .B2(n39794), .ZN(
        n7315) );
  NOR2_X1 U34872 ( .A1(n33752), .A2(n33753), .ZN(n33751) );
  NAND4_X1 U34873 ( .A1(n33754), .A2(n33755), .A3(n33756), .A4(n33757), .ZN(
        n33753) );
  NAND4_X1 U34874 ( .A1(n33762), .A2(n33763), .A3(n33764), .A4(n33765), .ZN(
        n33752) );
  OAI22_X1 U34875 ( .A1(n16990), .A2(n39548), .B1(n35025), .B2(n39542), .ZN(
        n7251) );
  NOR2_X1 U34876 ( .A1(n35026), .A2(n35027), .ZN(n35025) );
  NAND4_X1 U34877 ( .A1(n35028), .A2(n35029), .A3(n35030), .A4(n35031), .ZN(
        n35027) );
  NAND4_X1 U34878 ( .A1(n35036), .A2(n35037), .A3(n35038), .A4(n35039), .ZN(
        n35026) );
  OAI22_X1 U34879 ( .A1(n17053), .A2(n39800), .B1(n33770), .B2(n39793), .ZN(
        n7314) );
  NOR2_X1 U34880 ( .A1(n33771), .A2(n33772), .ZN(n33770) );
  NAND4_X1 U34881 ( .A1(n33773), .A2(n33774), .A3(n33775), .A4(n33776), .ZN(
        n33772) );
  NAND4_X1 U34882 ( .A1(n33781), .A2(n33782), .A3(n33783), .A4(n33784), .ZN(
        n33771) );
  OAI22_X1 U34883 ( .A1(n16989), .A2(n39548), .B1(n35044), .B2(n39541), .ZN(
        n7250) );
  NOR2_X1 U34884 ( .A1(n35045), .A2(n35046), .ZN(n35044) );
  NAND4_X1 U34885 ( .A1(n35047), .A2(n35048), .A3(n35049), .A4(n35050), .ZN(
        n35046) );
  NAND4_X1 U34886 ( .A1(n35055), .A2(n35056), .A3(n35057), .A4(n35058), .ZN(
        n35045) );
  OAI22_X1 U34887 ( .A1(n17052), .A2(n39799), .B1(n33789), .B2(n39793), .ZN(
        n7313) );
  NOR2_X1 U34888 ( .A1(n33790), .A2(n33791), .ZN(n33789) );
  NAND4_X1 U34889 ( .A1(n33792), .A2(n33793), .A3(n33794), .A4(n33795), .ZN(
        n33791) );
  NAND4_X1 U34890 ( .A1(n33800), .A2(n33801), .A3(n33802), .A4(n33803), .ZN(
        n33790) );
  OAI22_X1 U34891 ( .A1(n16988), .A2(n39547), .B1(n35063), .B2(n39541), .ZN(
        n7249) );
  NOR2_X1 U34892 ( .A1(n35064), .A2(n35065), .ZN(n35063) );
  NAND4_X1 U34893 ( .A1(n35066), .A2(n35067), .A3(n35068), .A4(n35069), .ZN(
        n35065) );
  NAND4_X1 U34894 ( .A1(n35074), .A2(n35075), .A3(n35076), .A4(n35077), .ZN(
        n35064) );
  OAI22_X1 U34895 ( .A1(n17051), .A2(n39799), .B1(n33808), .B2(n39793), .ZN(
        n7312) );
  NOR2_X1 U34896 ( .A1(n33809), .A2(n33810), .ZN(n33808) );
  NAND4_X1 U34897 ( .A1(n33811), .A2(n33812), .A3(n33813), .A4(n33814), .ZN(
        n33810) );
  NAND4_X1 U34898 ( .A1(n33819), .A2(n33820), .A3(n33821), .A4(n33822), .ZN(
        n33809) );
  OAI22_X1 U34899 ( .A1(n16987), .A2(n39547), .B1(n35082), .B2(n39541), .ZN(
        n7248) );
  NOR2_X1 U34900 ( .A1(n35083), .A2(n35084), .ZN(n35082) );
  NAND4_X1 U34901 ( .A1(n35085), .A2(n35086), .A3(n35087), .A4(n35088), .ZN(
        n35084) );
  NAND4_X1 U34902 ( .A1(n35093), .A2(n35094), .A3(n35095), .A4(n35096), .ZN(
        n35083) );
  OAI22_X1 U34903 ( .A1(n17050), .A2(n39799), .B1(n33827), .B2(n39793), .ZN(
        n7311) );
  NOR2_X1 U34904 ( .A1(n33828), .A2(n33829), .ZN(n33827) );
  NAND4_X1 U34905 ( .A1(n33830), .A2(n33831), .A3(n33832), .A4(n33833), .ZN(
        n33829) );
  NAND4_X1 U34906 ( .A1(n33838), .A2(n33839), .A3(n33840), .A4(n33841), .ZN(
        n33828) );
  OAI22_X1 U34907 ( .A1(n16986), .A2(n39547), .B1(n35101), .B2(n39541), .ZN(
        n7247) );
  NOR2_X1 U34908 ( .A1(n35102), .A2(n35103), .ZN(n35101) );
  NAND4_X1 U34909 ( .A1(n35104), .A2(n35105), .A3(n35106), .A4(n35107), .ZN(
        n35103) );
  NAND4_X1 U34910 ( .A1(n35112), .A2(n35113), .A3(n35114), .A4(n35115), .ZN(
        n35102) );
  OAI22_X1 U34911 ( .A1(n17049), .A2(n39799), .B1(n33846), .B2(n39793), .ZN(
        n7310) );
  NOR2_X1 U34912 ( .A1(n33847), .A2(n33848), .ZN(n33846) );
  NAND4_X1 U34913 ( .A1(n33849), .A2(n33850), .A3(n33851), .A4(n33852), .ZN(
        n33848) );
  NAND4_X1 U34914 ( .A1(n33857), .A2(n33858), .A3(n33859), .A4(n33860), .ZN(
        n33847) );
  OAI22_X1 U34915 ( .A1(n16985), .A2(n39547), .B1(n35120), .B2(n39541), .ZN(
        n7246) );
  NOR2_X1 U34916 ( .A1(n35121), .A2(n35122), .ZN(n35120) );
  NAND4_X1 U34917 ( .A1(n35123), .A2(n35124), .A3(n35125), .A4(n35126), .ZN(
        n35122) );
  NAND4_X1 U34918 ( .A1(n35131), .A2(n35132), .A3(n35133), .A4(n35134), .ZN(
        n35121) );
  OAI22_X1 U34919 ( .A1(n17048), .A2(n39799), .B1(n33865), .B2(n39793), .ZN(
        n7309) );
  NOR2_X1 U34920 ( .A1(n33866), .A2(n33867), .ZN(n33865) );
  NAND4_X1 U34921 ( .A1(n33868), .A2(n33869), .A3(n33870), .A4(n33871), .ZN(
        n33867) );
  NAND4_X1 U34922 ( .A1(n33876), .A2(n33877), .A3(n33878), .A4(n33879), .ZN(
        n33866) );
  OAI22_X1 U34923 ( .A1(n16984), .A2(n39547), .B1(n35139), .B2(n39541), .ZN(
        n7245) );
  NOR2_X1 U34924 ( .A1(n35140), .A2(n35141), .ZN(n35139) );
  NAND4_X1 U34925 ( .A1(n35142), .A2(n35143), .A3(n35144), .A4(n35145), .ZN(
        n35141) );
  NAND4_X1 U34926 ( .A1(n35150), .A2(n35151), .A3(n35152), .A4(n35153), .ZN(
        n35140) );
  OAI22_X1 U34927 ( .A1(n17047), .A2(n39799), .B1(n33884), .B2(n39793), .ZN(
        n7308) );
  NOR2_X1 U34928 ( .A1(n33885), .A2(n33886), .ZN(n33884) );
  NAND4_X1 U34929 ( .A1(n33887), .A2(n33888), .A3(n33889), .A4(n33890), .ZN(
        n33886) );
  NAND4_X1 U34930 ( .A1(n33895), .A2(n33896), .A3(n33897), .A4(n33898), .ZN(
        n33885) );
  OAI22_X1 U34931 ( .A1(n16983), .A2(n39547), .B1(n35158), .B2(n39541), .ZN(
        n7244) );
  NOR2_X1 U34932 ( .A1(n35159), .A2(n35160), .ZN(n35158) );
  NAND4_X1 U34933 ( .A1(n35161), .A2(n35162), .A3(n35163), .A4(n35164), .ZN(
        n35160) );
  NAND4_X1 U34934 ( .A1(n35169), .A2(n35170), .A3(n35171), .A4(n35172), .ZN(
        n35159) );
  OAI22_X1 U34935 ( .A1(n17046), .A2(n39799), .B1(n33903), .B2(n39793), .ZN(
        n7307) );
  NOR2_X1 U34936 ( .A1(n33904), .A2(n33905), .ZN(n33903) );
  NAND4_X1 U34937 ( .A1(n33906), .A2(n33907), .A3(n33908), .A4(n33909), .ZN(
        n33905) );
  NAND4_X1 U34938 ( .A1(n33914), .A2(n33915), .A3(n33916), .A4(n33917), .ZN(
        n33904) );
  OAI22_X1 U34939 ( .A1(n16982), .A2(n39547), .B1(n35177), .B2(n39541), .ZN(
        n7243) );
  NOR2_X1 U34940 ( .A1(n35178), .A2(n35179), .ZN(n35177) );
  NAND4_X1 U34941 ( .A1(n35180), .A2(n35181), .A3(n35182), .A4(n35183), .ZN(
        n35179) );
  NAND4_X1 U34942 ( .A1(n35188), .A2(n35189), .A3(n35190), .A4(n35191), .ZN(
        n35178) );
  OAI22_X1 U34943 ( .A1(n17045), .A2(n39799), .B1(n33922), .B2(n39793), .ZN(
        n7306) );
  NOR2_X1 U34944 ( .A1(n33923), .A2(n33924), .ZN(n33922) );
  NAND4_X1 U34945 ( .A1(n33925), .A2(n33926), .A3(n33927), .A4(n33928), .ZN(
        n33924) );
  NAND4_X1 U34946 ( .A1(n33933), .A2(n33934), .A3(n33935), .A4(n33936), .ZN(
        n33923) );
  OAI22_X1 U34947 ( .A1(n16981), .A2(n39547), .B1(n35196), .B2(n39541), .ZN(
        n7242) );
  NOR2_X1 U34948 ( .A1(n35197), .A2(n35198), .ZN(n35196) );
  NAND4_X1 U34949 ( .A1(n35199), .A2(n35200), .A3(n35201), .A4(n35202), .ZN(
        n35198) );
  NAND4_X1 U34950 ( .A1(n35207), .A2(n35208), .A3(n35209), .A4(n35210), .ZN(
        n35197) );
  OAI22_X1 U34951 ( .A1(n17044), .A2(n39799), .B1(n33941), .B2(n39793), .ZN(
        n7305) );
  NOR2_X1 U34952 ( .A1(n33942), .A2(n33943), .ZN(n33941) );
  NAND4_X1 U34953 ( .A1(n33944), .A2(n33945), .A3(n33946), .A4(n33947), .ZN(
        n33943) );
  NAND4_X1 U34954 ( .A1(n33952), .A2(n33953), .A3(n33954), .A4(n33955), .ZN(
        n33942) );
  OAI22_X1 U34955 ( .A1(n16980), .A2(n39547), .B1(n35215), .B2(n39541), .ZN(
        n7241) );
  NOR2_X1 U34956 ( .A1(n35216), .A2(n35217), .ZN(n35215) );
  NAND4_X1 U34957 ( .A1(n35218), .A2(n35219), .A3(n35220), .A4(n35221), .ZN(
        n35217) );
  NAND4_X1 U34958 ( .A1(n35226), .A2(n35227), .A3(n35228), .A4(n35229), .ZN(
        n35216) );
  OAI22_X1 U34959 ( .A1(n17043), .A2(n39799), .B1(n33960), .B2(n39793), .ZN(
        n7304) );
  NOR2_X1 U34960 ( .A1(n33961), .A2(n33962), .ZN(n33960) );
  NAND4_X1 U34961 ( .A1(n33963), .A2(n33964), .A3(n33965), .A4(n33966), .ZN(
        n33962) );
  NAND4_X1 U34962 ( .A1(n33971), .A2(n33972), .A3(n33973), .A4(n33974), .ZN(
        n33961) );
  OAI22_X1 U34963 ( .A1(n16979), .A2(n39547), .B1(n35234), .B2(n39541), .ZN(
        n7240) );
  NOR2_X1 U34964 ( .A1(n35235), .A2(n35236), .ZN(n35234) );
  NAND4_X1 U34965 ( .A1(n35237), .A2(n35238), .A3(n35239), .A4(n35240), .ZN(
        n35236) );
  NAND4_X1 U34966 ( .A1(n35245), .A2(n35246), .A3(n35247), .A4(n35248), .ZN(
        n35235) );
  OAI22_X1 U34967 ( .A1(n17042), .A2(n39799), .B1(n33979), .B2(n39793), .ZN(
        n7303) );
  NOR2_X1 U34968 ( .A1(n33980), .A2(n33981), .ZN(n33979) );
  NAND4_X1 U34969 ( .A1(n33982), .A2(n33983), .A3(n33984), .A4(n33985), .ZN(
        n33981) );
  NAND4_X1 U34970 ( .A1(n33990), .A2(n33991), .A3(n33992), .A4(n33993), .ZN(
        n33980) );
  OAI22_X1 U34971 ( .A1(n16978), .A2(n39547), .B1(n35253), .B2(n39541), .ZN(
        n7239) );
  NOR2_X1 U34972 ( .A1(n35254), .A2(n35255), .ZN(n35253) );
  NAND4_X1 U34973 ( .A1(n35256), .A2(n35257), .A3(n35258), .A4(n35259), .ZN(
        n35255) );
  NAND4_X1 U34974 ( .A1(n35264), .A2(n35265), .A3(n35266), .A4(n35267), .ZN(
        n35254) );
  OAI22_X1 U34975 ( .A1(n17041), .A2(n39799), .B1(n33998), .B2(n39792), .ZN(
        n7302) );
  NOR2_X1 U34976 ( .A1(n33999), .A2(n34000), .ZN(n33998) );
  NAND4_X1 U34977 ( .A1(n34001), .A2(n34002), .A3(n34003), .A4(n34004), .ZN(
        n34000) );
  NAND4_X1 U34978 ( .A1(n34009), .A2(n34010), .A3(n34011), .A4(n34012), .ZN(
        n33999) );
  OAI22_X1 U34979 ( .A1(n16977), .A2(n39547), .B1(n35272), .B2(n39540), .ZN(
        n7238) );
  NOR2_X1 U34980 ( .A1(n35273), .A2(n35274), .ZN(n35272) );
  NAND4_X1 U34981 ( .A1(n35275), .A2(n35276), .A3(n35277), .A4(n35278), .ZN(
        n35274) );
  NAND4_X1 U34982 ( .A1(n35283), .A2(n35284), .A3(n35285), .A4(n35286), .ZN(
        n35273) );
  OAI22_X1 U34983 ( .A1(n17040), .A2(n39798), .B1(n34017), .B2(n39792), .ZN(
        n7301) );
  NOR2_X1 U34984 ( .A1(n34018), .A2(n34019), .ZN(n34017) );
  NAND4_X1 U34985 ( .A1(n34020), .A2(n34021), .A3(n34022), .A4(n34023), .ZN(
        n34019) );
  NAND4_X1 U34986 ( .A1(n34028), .A2(n34029), .A3(n34030), .A4(n34031), .ZN(
        n34018) );
  OAI22_X1 U34987 ( .A1(n16976), .A2(n39546), .B1(n35291), .B2(n39540), .ZN(
        n7237) );
  NOR2_X1 U34988 ( .A1(n35292), .A2(n35293), .ZN(n35291) );
  NAND4_X1 U34989 ( .A1(n35294), .A2(n35295), .A3(n35296), .A4(n35297), .ZN(
        n35293) );
  NAND4_X1 U34990 ( .A1(n35302), .A2(n35303), .A3(n35304), .A4(n35305), .ZN(
        n35292) );
  OAI22_X1 U34991 ( .A1(n17039), .A2(n39798), .B1(n34036), .B2(n39792), .ZN(
        n7300) );
  NOR2_X1 U34992 ( .A1(n34037), .A2(n34038), .ZN(n34036) );
  NAND4_X1 U34993 ( .A1(n34039), .A2(n34040), .A3(n34041), .A4(n34042), .ZN(
        n34038) );
  NAND4_X1 U34994 ( .A1(n34047), .A2(n34048), .A3(n34049), .A4(n34050), .ZN(
        n34037) );
  OAI22_X1 U34995 ( .A1(n16975), .A2(n39546), .B1(n35310), .B2(n39540), .ZN(
        n7236) );
  NOR2_X1 U34996 ( .A1(n35311), .A2(n35312), .ZN(n35310) );
  NAND4_X1 U34997 ( .A1(n35313), .A2(n35314), .A3(n35315), .A4(n35316), .ZN(
        n35312) );
  NAND4_X1 U34998 ( .A1(n35321), .A2(n35322), .A3(n35323), .A4(n35324), .ZN(
        n35311) );
  OAI22_X1 U34999 ( .A1(n17038), .A2(n39798), .B1(n34055), .B2(n39792), .ZN(
        n7299) );
  NOR2_X1 U35000 ( .A1(n34056), .A2(n34057), .ZN(n34055) );
  NAND4_X1 U35001 ( .A1(n34058), .A2(n34059), .A3(n34060), .A4(n34061), .ZN(
        n34057) );
  NAND4_X1 U35002 ( .A1(n34066), .A2(n34067), .A3(n34068), .A4(n34069), .ZN(
        n34056) );
  OAI22_X1 U35003 ( .A1(n16974), .A2(n39546), .B1(n35329), .B2(n39540), .ZN(
        n7235) );
  NOR2_X1 U35004 ( .A1(n35330), .A2(n35331), .ZN(n35329) );
  NAND4_X1 U35005 ( .A1(n35332), .A2(n35333), .A3(n35334), .A4(n35335), .ZN(
        n35331) );
  NAND4_X1 U35006 ( .A1(n35340), .A2(n35341), .A3(n35342), .A4(n35343), .ZN(
        n35330) );
  OAI22_X1 U35007 ( .A1(n17037), .A2(n39798), .B1(n34074), .B2(n39792), .ZN(
        n7298) );
  NOR2_X1 U35008 ( .A1(n34075), .A2(n34076), .ZN(n34074) );
  NAND4_X1 U35009 ( .A1(n34077), .A2(n34078), .A3(n34079), .A4(n34080), .ZN(
        n34076) );
  NAND4_X1 U35010 ( .A1(n34085), .A2(n34086), .A3(n34087), .A4(n34088), .ZN(
        n34075) );
  OAI22_X1 U35011 ( .A1(n16973), .A2(n39546), .B1(n35348), .B2(n39540), .ZN(
        n7234) );
  NOR2_X1 U35012 ( .A1(n35349), .A2(n35350), .ZN(n35348) );
  NAND4_X1 U35013 ( .A1(n35351), .A2(n35352), .A3(n35353), .A4(n35354), .ZN(
        n35350) );
  NAND4_X1 U35014 ( .A1(n35359), .A2(n35360), .A3(n35361), .A4(n35362), .ZN(
        n35349) );
  OAI22_X1 U35015 ( .A1(n17036), .A2(n39798), .B1(n34093), .B2(n39792), .ZN(
        n7297) );
  NOR2_X1 U35016 ( .A1(n34094), .A2(n34095), .ZN(n34093) );
  NAND4_X1 U35017 ( .A1(n34096), .A2(n34097), .A3(n34098), .A4(n34099), .ZN(
        n34095) );
  NAND4_X1 U35018 ( .A1(n34104), .A2(n34105), .A3(n34106), .A4(n34107), .ZN(
        n34094) );
  OAI22_X1 U35019 ( .A1(n16972), .A2(n39546), .B1(n35367), .B2(n39540), .ZN(
        n7233) );
  NOR2_X1 U35020 ( .A1(n35368), .A2(n35369), .ZN(n35367) );
  NAND4_X1 U35021 ( .A1(n35370), .A2(n35371), .A3(n35372), .A4(n35373), .ZN(
        n35369) );
  NAND4_X1 U35022 ( .A1(n35378), .A2(n35379), .A3(n35380), .A4(n35381), .ZN(
        n35368) );
  OAI22_X1 U35023 ( .A1(n17035), .A2(n39798), .B1(n34112), .B2(n39792), .ZN(
        n7296) );
  NOR2_X1 U35024 ( .A1(n34113), .A2(n34114), .ZN(n34112) );
  NAND4_X1 U35025 ( .A1(n34115), .A2(n34116), .A3(n34117), .A4(n34118), .ZN(
        n34114) );
  NAND4_X1 U35026 ( .A1(n34123), .A2(n34124), .A3(n34125), .A4(n34126), .ZN(
        n34113) );
  OAI22_X1 U35027 ( .A1(n16971), .A2(n39546), .B1(n35386), .B2(n39540), .ZN(
        n7232) );
  NOR2_X1 U35028 ( .A1(n35387), .A2(n35388), .ZN(n35386) );
  NAND4_X1 U35029 ( .A1(n35389), .A2(n35390), .A3(n35391), .A4(n35392), .ZN(
        n35388) );
  NAND4_X1 U35030 ( .A1(n35397), .A2(n35398), .A3(n35399), .A4(n35400), .ZN(
        n35387) );
  OAI22_X1 U35031 ( .A1(n17034), .A2(n39798), .B1(n34131), .B2(n39792), .ZN(
        n7295) );
  NOR2_X1 U35032 ( .A1(n34132), .A2(n34133), .ZN(n34131) );
  NAND4_X1 U35033 ( .A1(n34134), .A2(n34135), .A3(n34136), .A4(n34137), .ZN(
        n34133) );
  NAND4_X1 U35034 ( .A1(n34142), .A2(n34143), .A3(n34144), .A4(n34145), .ZN(
        n34132) );
  OAI22_X1 U35035 ( .A1(n16970), .A2(n39546), .B1(n35405), .B2(n39540), .ZN(
        n7231) );
  NOR2_X1 U35036 ( .A1(n35406), .A2(n35407), .ZN(n35405) );
  NAND4_X1 U35037 ( .A1(n35408), .A2(n35409), .A3(n35410), .A4(n35411), .ZN(
        n35407) );
  NAND4_X1 U35038 ( .A1(n35416), .A2(n35417), .A3(n35418), .A4(n35419), .ZN(
        n35406) );
  OAI22_X1 U35039 ( .A1(n17033), .A2(n39798), .B1(n34150), .B2(n39792), .ZN(
        n7294) );
  NOR2_X1 U35040 ( .A1(n34151), .A2(n34152), .ZN(n34150) );
  NAND4_X1 U35041 ( .A1(n34153), .A2(n34154), .A3(n34155), .A4(n34156), .ZN(
        n34152) );
  NAND4_X1 U35042 ( .A1(n34161), .A2(n34162), .A3(n34163), .A4(n34164), .ZN(
        n34151) );
  OAI22_X1 U35043 ( .A1(n16969), .A2(n39546), .B1(n35424), .B2(n39540), .ZN(
        n7230) );
  NOR2_X1 U35044 ( .A1(n35425), .A2(n35426), .ZN(n35424) );
  NAND4_X1 U35045 ( .A1(n35427), .A2(n35428), .A3(n35429), .A4(n35430), .ZN(
        n35426) );
  NAND4_X1 U35046 ( .A1(n35435), .A2(n35436), .A3(n35437), .A4(n35438), .ZN(
        n35425) );
  OAI22_X1 U35047 ( .A1(n17032), .A2(n39798), .B1(n34169), .B2(n39792), .ZN(
        n7293) );
  NOR2_X1 U35048 ( .A1(n34170), .A2(n34171), .ZN(n34169) );
  NAND4_X1 U35049 ( .A1(n34172), .A2(n34173), .A3(n34174), .A4(n34175), .ZN(
        n34171) );
  NAND4_X1 U35050 ( .A1(n34180), .A2(n34181), .A3(n34182), .A4(n34183), .ZN(
        n34170) );
  OAI22_X1 U35051 ( .A1(n16968), .A2(n39546), .B1(n35443), .B2(n39540), .ZN(
        n7229) );
  NOR2_X1 U35052 ( .A1(n35444), .A2(n35445), .ZN(n35443) );
  NAND4_X1 U35053 ( .A1(n35446), .A2(n35447), .A3(n35448), .A4(n35449), .ZN(
        n35445) );
  NAND4_X1 U35054 ( .A1(n35454), .A2(n35455), .A3(n35456), .A4(n35457), .ZN(
        n35444) );
  OAI22_X1 U35055 ( .A1(n17031), .A2(n39798), .B1(n34188), .B2(n39792), .ZN(
        n7292) );
  NOR2_X1 U35056 ( .A1(n34189), .A2(n34190), .ZN(n34188) );
  NAND4_X1 U35057 ( .A1(n34191), .A2(n34192), .A3(n34193), .A4(n34194), .ZN(
        n34190) );
  NAND4_X1 U35058 ( .A1(n34199), .A2(n34200), .A3(n34201), .A4(n34202), .ZN(
        n34189) );
  OAI22_X1 U35059 ( .A1(n16967), .A2(n39546), .B1(n35462), .B2(n39540), .ZN(
        n7228) );
  NOR2_X1 U35060 ( .A1(n35463), .A2(n35464), .ZN(n35462) );
  NAND4_X1 U35061 ( .A1(n35465), .A2(n35466), .A3(n35467), .A4(n35468), .ZN(
        n35464) );
  NAND4_X1 U35062 ( .A1(n35473), .A2(n35474), .A3(n35475), .A4(n35476), .ZN(
        n35463) );
  OAI22_X1 U35063 ( .A1(n17030), .A2(n39798), .B1(n34207), .B2(n39792), .ZN(
        n7291) );
  NOR2_X1 U35064 ( .A1(n34208), .A2(n34209), .ZN(n34207) );
  NAND4_X1 U35065 ( .A1(n34210), .A2(n34211), .A3(n34212), .A4(n34213), .ZN(
        n34209) );
  NAND4_X1 U35066 ( .A1(n34218), .A2(n34219), .A3(n34220), .A4(n34221), .ZN(
        n34208) );
  OAI22_X1 U35067 ( .A1(n16966), .A2(n39546), .B1(n35481), .B2(n39540), .ZN(
        n7227) );
  NOR2_X1 U35068 ( .A1(n35482), .A2(n35483), .ZN(n35481) );
  NAND4_X1 U35069 ( .A1(n35484), .A2(n35485), .A3(n35486), .A4(n35487), .ZN(
        n35483) );
  NAND4_X1 U35070 ( .A1(n35492), .A2(n35493), .A3(n35494), .A4(n35495), .ZN(
        n35482) );
  OAI22_X1 U35071 ( .A1(n17029), .A2(n39798), .B1(n34226), .B2(n39791), .ZN(
        n7290) );
  NOR2_X1 U35072 ( .A1(n34227), .A2(n34228), .ZN(n34226) );
  NAND4_X1 U35073 ( .A1(n34229), .A2(n34230), .A3(n34231), .A4(n34232), .ZN(
        n34228) );
  NAND4_X1 U35074 ( .A1(n34237), .A2(n34238), .A3(n34239), .A4(n34240), .ZN(
        n34227) );
  OAI22_X1 U35075 ( .A1(n16965), .A2(n39546), .B1(n35500), .B2(n39539), .ZN(
        n7226) );
  NOR2_X1 U35076 ( .A1(n35501), .A2(n35502), .ZN(n35500) );
  NAND4_X1 U35077 ( .A1(n35503), .A2(n35504), .A3(n35505), .A4(n35506), .ZN(
        n35502) );
  NAND4_X1 U35078 ( .A1(n35511), .A2(n35512), .A3(n35513), .A4(n35514), .ZN(
        n35501) );
  OAI22_X1 U35079 ( .A1(n17028), .A2(n39797), .B1(n34245), .B2(n39791), .ZN(
        n7289) );
  NOR2_X1 U35080 ( .A1(n34246), .A2(n34247), .ZN(n34245) );
  NAND4_X1 U35081 ( .A1(n34248), .A2(n34249), .A3(n34250), .A4(n34251), .ZN(
        n34247) );
  NAND4_X1 U35082 ( .A1(n34256), .A2(n34257), .A3(n34258), .A4(n34259), .ZN(
        n34246) );
  OAI22_X1 U35083 ( .A1(n16964), .A2(n39545), .B1(n35519), .B2(n39539), .ZN(
        n7225) );
  NOR2_X1 U35084 ( .A1(n35520), .A2(n35521), .ZN(n35519) );
  NAND4_X1 U35085 ( .A1(n35522), .A2(n35523), .A3(n35524), .A4(n35525), .ZN(
        n35521) );
  NAND4_X1 U35086 ( .A1(n35530), .A2(n35531), .A3(n35532), .A4(n35533), .ZN(
        n35520) );
  OAI22_X1 U35087 ( .A1(n17027), .A2(n39797), .B1(n34264), .B2(n39791), .ZN(
        n7288) );
  NOR2_X1 U35088 ( .A1(n34265), .A2(n34266), .ZN(n34264) );
  NAND4_X1 U35089 ( .A1(n34267), .A2(n34268), .A3(n34269), .A4(n34270), .ZN(
        n34266) );
  NAND4_X1 U35090 ( .A1(n34275), .A2(n34276), .A3(n34277), .A4(n34278), .ZN(
        n34265) );
  OAI22_X1 U35091 ( .A1(n16963), .A2(n39545), .B1(n35538), .B2(n39539), .ZN(
        n7224) );
  NOR2_X1 U35092 ( .A1(n35539), .A2(n35540), .ZN(n35538) );
  NAND4_X1 U35093 ( .A1(n35541), .A2(n35542), .A3(n35543), .A4(n35544), .ZN(
        n35540) );
  NAND4_X1 U35094 ( .A1(n35549), .A2(n35550), .A3(n35551), .A4(n35552), .ZN(
        n35539) );
  OAI22_X1 U35095 ( .A1(n17026), .A2(n39797), .B1(n34283), .B2(n39791), .ZN(
        n7287) );
  NOR2_X1 U35096 ( .A1(n34284), .A2(n34285), .ZN(n34283) );
  NAND4_X1 U35097 ( .A1(n34286), .A2(n34287), .A3(n34288), .A4(n34289), .ZN(
        n34285) );
  NAND4_X1 U35098 ( .A1(n34294), .A2(n34295), .A3(n34296), .A4(n34297), .ZN(
        n34284) );
  OAI22_X1 U35099 ( .A1(n16962), .A2(n39545), .B1(n35557), .B2(n39539), .ZN(
        n7223) );
  NOR2_X1 U35100 ( .A1(n35558), .A2(n35559), .ZN(n35557) );
  NAND4_X1 U35101 ( .A1(n35560), .A2(n35561), .A3(n35562), .A4(n35563), .ZN(
        n35559) );
  NAND4_X1 U35102 ( .A1(n35568), .A2(n35569), .A3(n35570), .A4(n35571), .ZN(
        n35558) );
  OAI22_X1 U35103 ( .A1(n17025), .A2(n39797), .B1(n34302), .B2(n39791), .ZN(
        n7286) );
  NOR2_X1 U35104 ( .A1(n34303), .A2(n34304), .ZN(n34302) );
  NAND4_X1 U35105 ( .A1(n34305), .A2(n34306), .A3(n34307), .A4(n34308), .ZN(
        n34304) );
  NAND4_X1 U35106 ( .A1(n34313), .A2(n34314), .A3(n34315), .A4(n34316), .ZN(
        n34303) );
  OAI22_X1 U35107 ( .A1(n16961), .A2(n39545), .B1(n35576), .B2(n39539), .ZN(
        n7222) );
  NOR2_X1 U35108 ( .A1(n35577), .A2(n35578), .ZN(n35576) );
  NAND4_X1 U35109 ( .A1(n35579), .A2(n35580), .A3(n35581), .A4(n35582), .ZN(
        n35578) );
  NAND4_X1 U35110 ( .A1(n35587), .A2(n35588), .A3(n35589), .A4(n35590), .ZN(
        n35577) );
  OAI22_X1 U35111 ( .A1(n17024), .A2(n39797), .B1(n34321), .B2(n39791), .ZN(
        n7285) );
  NOR2_X1 U35112 ( .A1(n34322), .A2(n34323), .ZN(n34321) );
  NAND4_X1 U35113 ( .A1(n34324), .A2(n34325), .A3(n34326), .A4(n34327), .ZN(
        n34323) );
  NAND4_X1 U35114 ( .A1(n34332), .A2(n34333), .A3(n34334), .A4(n34335), .ZN(
        n34322) );
  OAI22_X1 U35115 ( .A1(n16960), .A2(n39545), .B1(n35595), .B2(n39539), .ZN(
        n7221) );
  NOR2_X1 U35116 ( .A1(n35596), .A2(n35597), .ZN(n35595) );
  NAND4_X1 U35117 ( .A1(n35598), .A2(n35599), .A3(n35600), .A4(n35601), .ZN(
        n35597) );
  NAND4_X1 U35118 ( .A1(n35606), .A2(n35607), .A3(n35608), .A4(n35609), .ZN(
        n35596) );
  OAI22_X1 U35119 ( .A1(n17023), .A2(n39797), .B1(n34340), .B2(n39791), .ZN(
        n7284) );
  NOR2_X1 U35120 ( .A1(n34341), .A2(n34342), .ZN(n34340) );
  NAND4_X1 U35121 ( .A1(n34343), .A2(n34344), .A3(n34345), .A4(n34346), .ZN(
        n34342) );
  NAND4_X1 U35122 ( .A1(n34351), .A2(n34352), .A3(n34353), .A4(n34354), .ZN(
        n34341) );
  OAI22_X1 U35123 ( .A1(n16959), .A2(n39545), .B1(n35614), .B2(n39539), .ZN(
        n7220) );
  NOR2_X1 U35124 ( .A1(n35615), .A2(n35616), .ZN(n35614) );
  NAND4_X1 U35125 ( .A1(n35617), .A2(n35618), .A3(n35619), .A4(n35620), .ZN(
        n35616) );
  NAND4_X1 U35126 ( .A1(n35625), .A2(n35626), .A3(n35627), .A4(n35628), .ZN(
        n35615) );
  OAI22_X1 U35127 ( .A1(n17022), .A2(n39797), .B1(n34359), .B2(n39791), .ZN(
        n7283) );
  NOR2_X1 U35128 ( .A1(n34360), .A2(n34361), .ZN(n34359) );
  NAND4_X1 U35129 ( .A1(n34362), .A2(n34363), .A3(n34364), .A4(n34365), .ZN(
        n34361) );
  NAND4_X1 U35130 ( .A1(n34370), .A2(n34371), .A3(n34372), .A4(n34373), .ZN(
        n34360) );
  OAI22_X1 U35131 ( .A1(n16958), .A2(n39545), .B1(n35633), .B2(n39539), .ZN(
        n7219) );
  NOR2_X1 U35132 ( .A1(n35634), .A2(n35635), .ZN(n35633) );
  NAND4_X1 U35133 ( .A1(n35636), .A2(n35637), .A3(n35638), .A4(n35639), .ZN(
        n35635) );
  NAND4_X1 U35134 ( .A1(n35644), .A2(n35645), .A3(n35646), .A4(n35647), .ZN(
        n35634) );
  OAI22_X1 U35135 ( .A1(n17021), .A2(n39797), .B1(n34378), .B2(n39791), .ZN(
        n7282) );
  NOR2_X1 U35136 ( .A1(n34379), .A2(n34380), .ZN(n34378) );
  NAND4_X1 U35137 ( .A1(n34381), .A2(n34382), .A3(n34383), .A4(n34384), .ZN(
        n34380) );
  NAND4_X1 U35138 ( .A1(n34389), .A2(n34390), .A3(n34391), .A4(n34392), .ZN(
        n34379) );
  OAI22_X1 U35139 ( .A1(n16957), .A2(n39545), .B1(n35652), .B2(n39539), .ZN(
        n7218) );
  NOR2_X1 U35140 ( .A1(n35653), .A2(n35654), .ZN(n35652) );
  NAND4_X1 U35141 ( .A1(n35655), .A2(n35656), .A3(n35657), .A4(n35658), .ZN(
        n35654) );
  NAND4_X1 U35142 ( .A1(n35663), .A2(n35664), .A3(n35665), .A4(n35666), .ZN(
        n35653) );
  OAI22_X1 U35143 ( .A1(n17020), .A2(n39797), .B1(n34397), .B2(n39791), .ZN(
        n7281) );
  NOR2_X1 U35144 ( .A1(n34398), .A2(n34399), .ZN(n34397) );
  NAND4_X1 U35145 ( .A1(n34400), .A2(n34401), .A3(n34402), .A4(n34403), .ZN(
        n34399) );
  NAND4_X1 U35146 ( .A1(n34408), .A2(n34409), .A3(n34410), .A4(n34411), .ZN(
        n34398) );
  OAI22_X1 U35147 ( .A1(n16956), .A2(n39545), .B1(n35671), .B2(n39539), .ZN(
        n7217) );
  NOR2_X1 U35148 ( .A1(n35672), .A2(n35673), .ZN(n35671) );
  NAND4_X1 U35149 ( .A1(n35674), .A2(n35675), .A3(n35676), .A4(n35677), .ZN(
        n35673) );
  NAND4_X1 U35150 ( .A1(n35682), .A2(n35683), .A3(n35684), .A4(n35685), .ZN(
        n35672) );
  OAI22_X1 U35151 ( .A1(n17019), .A2(n39797), .B1(n34416), .B2(n39791), .ZN(
        n7280) );
  NOR2_X1 U35152 ( .A1(n34417), .A2(n34418), .ZN(n34416) );
  NAND4_X1 U35153 ( .A1(n34419), .A2(n34420), .A3(n34421), .A4(n34422), .ZN(
        n34418) );
  NAND4_X1 U35154 ( .A1(n34427), .A2(n34428), .A3(n34429), .A4(n34430), .ZN(
        n34417) );
  OAI22_X1 U35155 ( .A1(n16955), .A2(n39545), .B1(n35690), .B2(n39539), .ZN(
        n7216) );
  NOR2_X1 U35156 ( .A1(n35691), .A2(n35692), .ZN(n35690) );
  NAND4_X1 U35157 ( .A1(n35693), .A2(n35694), .A3(n35695), .A4(n35696), .ZN(
        n35692) );
  NAND4_X1 U35158 ( .A1(n35701), .A2(n35702), .A3(n35703), .A4(n35704), .ZN(
        n35691) );
  OAI22_X1 U35159 ( .A1(n17018), .A2(n39797), .B1(n34435), .B2(n39791), .ZN(
        n7279) );
  NOR2_X1 U35160 ( .A1(n34436), .A2(n34437), .ZN(n34435) );
  NAND4_X1 U35161 ( .A1(n34438), .A2(n34439), .A3(n34440), .A4(n34441), .ZN(
        n34437) );
  NAND4_X1 U35162 ( .A1(n34446), .A2(n34447), .A3(n34448), .A4(n34449), .ZN(
        n34436) );
  OAI22_X1 U35163 ( .A1(n16954), .A2(n39545), .B1(n35709), .B2(n39539), .ZN(
        n7215) );
  NOR2_X1 U35164 ( .A1(n35710), .A2(n35711), .ZN(n35709) );
  NAND4_X1 U35165 ( .A1(n35712), .A2(n35713), .A3(n35714), .A4(n35715), .ZN(
        n35711) );
  NAND4_X1 U35166 ( .A1(n35720), .A2(n35721), .A3(n35722), .A4(n35723), .ZN(
        n35710) );
  OAI22_X1 U35167 ( .A1(n17017), .A2(n39797), .B1(n34454), .B2(n39790), .ZN(
        n7278) );
  NOR2_X1 U35168 ( .A1(n34455), .A2(n34456), .ZN(n34454) );
  NAND4_X1 U35169 ( .A1(n34457), .A2(n34458), .A3(n34459), .A4(n34460), .ZN(
        n34456) );
  NAND4_X1 U35170 ( .A1(n34465), .A2(n34466), .A3(n34467), .A4(n34468), .ZN(
        n34455) );
  OAI22_X1 U35171 ( .A1(n16953), .A2(n39545), .B1(n35728), .B2(n39538), .ZN(
        n7214) );
  NOR2_X1 U35172 ( .A1(n35729), .A2(n35730), .ZN(n35728) );
  NAND4_X1 U35173 ( .A1(n35731), .A2(n35732), .A3(n35733), .A4(n35734), .ZN(
        n35730) );
  NAND4_X1 U35174 ( .A1(n35739), .A2(n35740), .A3(n35741), .A4(n35742), .ZN(
        n35729) );
  OAI22_X1 U35175 ( .A1(n17016), .A2(n39796), .B1(n34473), .B2(n39790), .ZN(
        n7277) );
  NOR2_X1 U35176 ( .A1(n34474), .A2(n34475), .ZN(n34473) );
  NAND4_X1 U35177 ( .A1(n34476), .A2(n34477), .A3(n34478), .A4(n34479), .ZN(
        n34475) );
  NAND4_X1 U35178 ( .A1(n34484), .A2(n34485), .A3(n34486), .A4(n34487), .ZN(
        n34474) );
  OAI22_X1 U35179 ( .A1(n16952), .A2(n39544), .B1(n35747), .B2(n39538), .ZN(
        n7213) );
  NOR2_X1 U35180 ( .A1(n35748), .A2(n35749), .ZN(n35747) );
  NAND4_X1 U35181 ( .A1(n35750), .A2(n35751), .A3(n35752), .A4(n35753), .ZN(
        n35749) );
  NAND4_X1 U35182 ( .A1(n35758), .A2(n35759), .A3(n35760), .A4(n35761), .ZN(
        n35748) );
  OAI22_X1 U35183 ( .A1(n17015), .A2(n39796), .B1(n34492), .B2(n39790), .ZN(
        n7276) );
  NOR2_X1 U35184 ( .A1(n34493), .A2(n34494), .ZN(n34492) );
  NAND4_X1 U35185 ( .A1(n34495), .A2(n34496), .A3(n34497), .A4(n34498), .ZN(
        n34494) );
  NAND4_X1 U35186 ( .A1(n34503), .A2(n34504), .A3(n34505), .A4(n34506), .ZN(
        n34493) );
  OAI22_X1 U35187 ( .A1(n16951), .A2(n39544), .B1(n35766), .B2(n39538), .ZN(
        n7212) );
  NOR2_X1 U35188 ( .A1(n35767), .A2(n35768), .ZN(n35766) );
  NAND4_X1 U35189 ( .A1(n35769), .A2(n35770), .A3(n35771), .A4(n35772), .ZN(
        n35768) );
  NAND4_X1 U35190 ( .A1(n35777), .A2(n35778), .A3(n35779), .A4(n35780), .ZN(
        n35767) );
  OAI22_X1 U35191 ( .A1(n17014), .A2(n39796), .B1(n34511), .B2(n39790), .ZN(
        n7275) );
  NOR2_X1 U35192 ( .A1(n34512), .A2(n34513), .ZN(n34511) );
  NAND4_X1 U35193 ( .A1(n34514), .A2(n34515), .A3(n34516), .A4(n34517), .ZN(
        n34513) );
  NAND4_X1 U35194 ( .A1(n34522), .A2(n34523), .A3(n34524), .A4(n34525), .ZN(
        n34512) );
  OAI22_X1 U35195 ( .A1(n16950), .A2(n39544), .B1(n35785), .B2(n39538), .ZN(
        n7211) );
  NOR2_X1 U35196 ( .A1(n35786), .A2(n35787), .ZN(n35785) );
  NAND4_X1 U35197 ( .A1(n35788), .A2(n35789), .A3(n35790), .A4(n35791), .ZN(
        n35787) );
  NAND4_X1 U35198 ( .A1(n35796), .A2(n35797), .A3(n35798), .A4(n35799), .ZN(
        n35786) );
  OAI22_X1 U35199 ( .A1(n17013), .A2(n39796), .B1(n34530), .B2(n39790), .ZN(
        n7274) );
  NOR2_X1 U35200 ( .A1(n34531), .A2(n34532), .ZN(n34530) );
  NAND4_X1 U35201 ( .A1(n34533), .A2(n34534), .A3(n34535), .A4(n34536), .ZN(
        n34532) );
  NAND4_X1 U35202 ( .A1(n34541), .A2(n34542), .A3(n34543), .A4(n34544), .ZN(
        n34531) );
  OAI22_X1 U35203 ( .A1(n16949), .A2(n39544), .B1(n35804), .B2(n39538), .ZN(
        n7210) );
  NOR2_X1 U35204 ( .A1(n35805), .A2(n35806), .ZN(n35804) );
  NAND4_X1 U35205 ( .A1(n35807), .A2(n35808), .A3(n35809), .A4(n35810), .ZN(
        n35806) );
  NAND4_X1 U35206 ( .A1(n35815), .A2(n35816), .A3(n35817), .A4(n35818), .ZN(
        n35805) );
  OAI22_X1 U35207 ( .A1(n17012), .A2(n39796), .B1(n34549), .B2(n39790), .ZN(
        n7273) );
  NOR2_X1 U35208 ( .A1(n34550), .A2(n34551), .ZN(n34549) );
  NAND4_X1 U35209 ( .A1(n34552), .A2(n34553), .A3(n34554), .A4(n34555), .ZN(
        n34551) );
  NAND4_X1 U35210 ( .A1(n34560), .A2(n34561), .A3(n34562), .A4(n34563), .ZN(
        n34550) );
  OAI22_X1 U35211 ( .A1(n16948), .A2(n39544), .B1(n35823), .B2(n39538), .ZN(
        n7209) );
  NOR2_X1 U35212 ( .A1(n35824), .A2(n35825), .ZN(n35823) );
  NAND4_X1 U35213 ( .A1(n35826), .A2(n35827), .A3(n35828), .A4(n35829), .ZN(
        n35825) );
  NAND4_X1 U35214 ( .A1(n35834), .A2(n35835), .A3(n35836), .A4(n35837), .ZN(
        n35824) );
  OAI22_X1 U35215 ( .A1(n17011), .A2(n39796), .B1(n34568), .B2(n39790), .ZN(
        n7272) );
  NOR2_X1 U35216 ( .A1(n34569), .A2(n34570), .ZN(n34568) );
  NAND4_X1 U35217 ( .A1(n34571), .A2(n34572), .A3(n34573), .A4(n34574), .ZN(
        n34570) );
  NAND4_X1 U35218 ( .A1(n34579), .A2(n34580), .A3(n34581), .A4(n34582), .ZN(
        n34569) );
  OAI22_X1 U35219 ( .A1(n16947), .A2(n39544), .B1(n35842), .B2(n39538), .ZN(
        n7208) );
  NOR2_X1 U35220 ( .A1(n35843), .A2(n35844), .ZN(n35842) );
  NAND4_X1 U35221 ( .A1(n35845), .A2(n35846), .A3(n35847), .A4(n35848), .ZN(
        n35844) );
  NAND4_X1 U35222 ( .A1(n35853), .A2(n35854), .A3(n35855), .A4(n35856), .ZN(
        n35843) );
  OAI22_X1 U35223 ( .A1(n17010), .A2(n39796), .B1(n34587), .B2(n39790), .ZN(
        n7271) );
  NOR2_X1 U35224 ( .A1(n34588), .A2(n34589), .ZN(n34587) );
  NAND4_X1 U35225 ( .A1(n34590), .A2(n34591), .A3(n34592), .A4(n34593), .ZN(
        n34589) );
  NAND4_X1 U35226 ( .A1(n34598), .A2(n34599), .A3(n34600), .A4(n34601), .ZN(
        n34588) );
  OAI22_X1 U35227 ( .A1(n16946), .A2(n39544), .B1(n35861), .B2(n39538), .ZN(
        n7207) );
  NOR2_X1 U35228 ( .A1(n35862), .A2(n35863), .ZN(n35861) );
  NAND4_X1 U35229 ( .A1(n35864), .A2(n35865), .A3(n35866), .A4(n35867), .ZN(
        n35863) );
  NAND4_X1 U35230 ( .A1(n35872), .A2(n35873), .A3(n35874), .A4(n35875), .ZN(
        n35862) );
  OAI22_X1 U35231 ( .A1(n17009), .A2(n39796), .B1(n34606), .B2(n39790), .ZN(
        n7270) );
  NOR2_X1 U35232 ( .A1(n34607), .A2(n34608), .ZN(n34606) );
  NAND4_X1 U35233 ( .A1(n34609), .A2(n34610), .A3(n34611), .A4(n34612), .ZN(
        n34608) );
  NAND4_X1 U35234 ( .A1(n34617), .A2(n34618), .A3(n34619), .A4(n34620), .ZN(
        n34607) );
  OAI22_X1 U35235 ( .A1(n16945), .A2(n39544), .B1(n35880), .B2(n39538), .ZN(
        n7206) );
  NOR2_X1 U35236 ( .A1(n35881), .A2(n35882), .ZN(n35880) );
  NAND4_X1 U35237 ( .A1(n35883), .A2(n35884), .A3(n35885), .A4(n35886), .ZN(
        n35882) );
  NAND4_X1 U35238 ( .A1(n35891), .A2(n35892), .A3(n35893), .A4(n35894), .ZN(
        n35881) );
  OAI22_X1 U35239 ( .A1(n17008), .A2(n39796), .B1(n34625), .B2(n39790), .ZN(
        n7269) );
  NOR2_X1 U35240 ( .A1(n34626), .A2(n34627), .ZN(n34625) );
  NAND4_X1 U35241 ( .A1(n34628), .A2(n34629), .A3(n34630), .A4(n34631), .ZN(
        n34627) );
  NAND4_X1 U35242 ( .A1(n34636), .A2(n34637), .A3(n34638), .A4(n34639), .ZN(
        n34626) );
  OAI22_X1 U35243 ( .A1(n16944), .A2(n39544), .B1(n35899), .B2(n39538), .ZN(
        n7205) );
  NOR2_X1 U35244 ( .A1(n35900), .A2(n35901), .ZN(n35899) );
  NAND4_X1 U35245 ( .A1(n35902), .A2(n35903), .A3(n35904), .A4(n35905), .ZN(
        n35901) );
  NAND4_X1 U35246 ( .A1(n35910), .A2(n35911), .A3(n35912), .A4(n35913), .ZN(
        n35900) );
  OAI22_X1 U35247 ( .A1(n17007), .A2(n39796), .B1(n34644), .B2(n39790), .ZN(
        n7268) );
  NOR2_X1 U35248 ( .A1(n34645), .A2(n34646), .ZN(n34644) );
  NAND4_X1 U35249 ( .A1(n34647), .A2(n34648), .A3(n34649), .A4(n34650), .ZN(
        n34646) );
  NAND4_X1 U35250 ( .A1(n34655), .A2(n34656), .A3(n34657), .A4(n34658), .ZN(
        n34645) );
  OAI22_X1 U35251 ( .A1(n16943), .A2(n39544), .B1(n35918), .B2(n39538), .ZN(
        n7204) );
  NOR2_X1 U35252 ( .A1(n35919), .A2(n35920), .ZN(n35918) );
  NAND4_X1 U35253 ( .A1(n35921), .A2(n35922), .A3(n35923), .A4(n35924), .ZN(
        n35920) );
  NAND4_X1 U35254 ( .A1(n35929), .A2(n35930), .A3(n35931), .A4(n35932), .ZN(
        n35919) );
  OAI22_X1 U35255 ( .A1(n17006), .A2(n39796), .B1(n34663), .B2(n39790), .ZN(
        n7267) );
  NOR2_X1 U35256 ( .A1(n34664), .A2(n34665), .ZN(n34663) );
  NAND4_X1 U35257 ( .A1(n34666), .A2(n34667), .A3(n34668), .A4(n34669), .ZN(
        n34665) );
  NAND4_X1 U35258 ( .A1(n34685), .A2(n34686), .A3(n34687), .A4(n34688), .ZN(
        n34664) );
  OAI22_X1 U35259 ( .A1(n16942), .A2(n39544), .B1(n35937), .B2(n39538), .ZN(
        n7203) );
  NOR2_X1 U35260 ( .A1(n35938), .A2(n35939), .ZN(n35937) );
  NAND4_X1 U35261 ( .A1(n35940), .A2(n35941), .A3(n35942), .A4(n35943), .ZN(
        n35939) );
  NAND4_X1 U35262 ( .A1(n35959), .A2(n35960), .A3(n35961), .A4(n35962), .ZN(
        n35938) );
  NOR2_X1 U35263 ( .A1(n2699), .A2(n2710), .ZN(n12791) );
  NOR2_X1 U35264 ( .A1(n2695), .A2(n32167), .ZN(\U3/U194/Z_4 ) );
  NOR2_X1 U35265 ( .A1(n2695), .A2(n32172), .ZN(\U3/U195/Z_4 ) );
  AND2_X1 U35266 ( .A1(n33301), .A2(WR), .ZN(n33330) );
  NOR2_X1 U35267 ( .A1(n2698), .A2(n32167), .ZN(\U3/U194/Z_1 ) );
  AND3_X1 U35268 ( .A1(ADD_RD1[0]), .A2(n32253), .A3(n33208), .ZN(\r504/n3 )
         );
  NOR2_X1 U35269 ( .A1(n2698), .A2(n32172), .ZN(\U3/U195/Z_1 ) );
  AND3_X1 U35270 ( .A1(ADD_RD2[0]), .A2(n32253), .A3(n33207), .ZN(\r510/n3 )
         );
  NOR2_X1 U35271 ( .A1(n2697), .A2(n32167), .ZN(\U3/U194/Z_2 ) );
  NOR2_X1 U35272 ( .A1(n2697), .A2(n32172), .ZN(\U3/U195/Z_2 ) );
  NOR2_X1 U35273 ( .A1(n2698), .A2(n32162), .ZN(\U3/U193/Z_1 ) );
  AND3_X1 U35274 ( .A1(ADD_WR[0]), .A2(n32253), .A3(n33209), .ZN(\r498/n1 ) );
  NAND2_X1 U35275 ( .A1(n2696), .A2(n33208), .ZN(\U3/U194/Z_3 ) );
  NAND2_X1 U35276 ( .A1(n2696), .A2(n33207), .ZN(\U3/U195/Z_3 ) );
  NOR2_X1 U35277 ( .A1(n2697), .A2(n32162), .ZN(\U3/U193/Z_2 ) );
  NAND2_X1 U35278 ( .A1(n2696), .A2(n33209), .ZN(\U3/U193/Z_3 ) );
  NOR3_X1 U35279 ( .A1(n32075), .A2(RESET), .A3(n33227), .ZN(n33223) );
  OAI222_X1 U35280 ( .A1(n32240), .A2(n33211), .B1(n33215), .B2(n33213), .C1(
        n2683), .C2(n33212), .ZN(n9902) );
  INV_X1 U35281 ( .A(n33215), .ZN(n32240) );
  OAI22_X1 U35282 ( .A1(n33250), .A2(\i[2] ), .B1(n2707), .B2(n33251), .ZN(
        n9891) );
  AOI211_X1 U35283 ( .C1(n2709), .C2(n33249), .A(n32077), .B(n32076), .ZN(
        n33251) );
  NAND4_X1 U35284 ( .A1(n2699), .A2(n2698), .A3(n35979), .A4(n2697), .ZN(
        n33218) );
  NOR2_X1 U35285 ( .A1(n2695), .A2(N661), .ZN(n35979) );
  XNOR2_X1 U35286 ( .A(n32244), .B(n2695), .ZN(n33215) );
  OAI21_X1 U35287 ( .B1(n23853), .B2(n32081), .A(n39297), .ZN(n33233) );
  NAND4_X1 U35288 ( .A1(n33238), .A2(n33239), .A3(n32238), .A4(n33240), .ZN(
        n33227) );
  NOR4_X1 U35289 ( .A1(n33241), .A2(n32083), .A3(n33242), .A4(n33243), .ZN(
        n33240) );
  INV_X1 U35290 ( .A(n33244), .ZN(n32238) );
  OAI211_X1 U35291 ( .C1(n35974), .C2(n35975), .A(ENABLE), .B(CALL), .ZN(
        n33232) );
  NOR4_X1 U35292 ( .A1(n35976), .A2(n33218), .A3(n32259), .A4(n32261), .ZN(
        n35975) );
  NOR4_X1 U35293 ( .A1(n35977), .A2(n35978), .A3(n33242), .A4(n33243), .ZN(
        n35974) );
  NAND4_X1 U35294 ( .A1(n2695), .A2(n2683), .A3(n33246), .A4(n2699), .ZN(
        n33216) );
  AND2_X1 U35295 ( .A1(n2696), .A2(n2697), .ZN(n33246) );
  XNOR2_X1 U35296 ( .A(n32322), .B(n2695), .ZN(n33238) );
  OAI211_X1 U35297 ( .C1(N659), .C2(n33216), .A(RETRN), .B(n33217), .ZN(n33213) );
  AND2_X1 U35298 ( .A1(n41370), .A2(n33212), .ZN(n33217) );
  OAI22_X1 U35299 ( .A1(n33220), .A2(n32323), .B1(n27870), .B2(n33221), .ZN(
        n9901) );
  AOI221_X1 U35300 ( .B1(n33223), .B2(n27872), .C1(n33222), .C2(n32322), .A(
        n32075), .ZN(n33220) );
  AOI22_X1 U35301 ( .A1(n33222), .A2(n27872), .B1(n33223), .B2(n32322), .ZN(
        n33221) );
  OAI22_X1 U35302 ( .A1(n2707), .A2(n33250), .B1(n2706), .B2(n37252), .ZN(
        n25394) );
  NOR2_X1 U35303 ( .A1(n33249), .A2(n32077), .ZN(n37252) );
  OR4_X1 U35304 ( .A1(n2706), .A2(n2707), .A3(n2709), .A4(n2710), .ZN(n33237)
         );
  OAI21_X1 U35305 ( .B1(n2695), .B2(n33212), .A(n33214), .ZN(n9903) );
  NAND2_X1 U35306 ( .A1(n33247), .A2(n33248), .ZN(n9892) );
  OAI21_X1 U35307 ( .B1(n32076), .B2(n32077), .A(\i[1] ), .ZN(n33247) );
  OAI21_X1 U35308 ( .B1(n23853), .B2(n33235), .A(n33236), .ZN(n9893) );
  OAI211_X1 U35309 ( .C1(n23853), .C2(n33237), .A(n33235), .B(n41368), .ZN(
        n33236) );
  OAI22_X1 U35310 ( .A1(n23853), .A2(n32081), .B1(n33231), .B2(n33230), .ZN(
        n33235) );
  OAI21_X1 U35311 ( .B1(n2700), .B2(n39296), .A(n35973), .ZN(n7202) );
  OAI221_X1 U35312 ( .B1(n32080), .B2(n39294), .C1(n2700), .C2(n33237), .A(
        n41364), .ZN(n35973) );
  INV_X1 U35313 ( .A(n33232), .ZN(n32080) );
  NAND2_X1 U35314 ( .A1(n2710), .A2(n33249), .ZN(n33234) );
  INV_X1 U35315 ( .A(n35972), .ZN(n39297) );
  OAI21_X1 U35316 ( .B1(n2700), .B2(n33231), .A(n41370), .ZN(n35972) );
  OAI21_X1 U35317 ( .B1(n2710), .B2(n33233), .A(n33234), .ZN(n9895) );
  AND4_X1 U35318 ( .A1(n33228), .A2(n33227), .A3(n33225), .A4(n41364), .ZN(
        n33222) );
  NAND4_X1 U35319 ( .A1(n27872), .A2(n27871), .A3(n33229), .A4(n27874), .ZN(
        n33228) );
  NOR2_X1 U35320 ( .A1(n38789), .A2(n38790), .ZN(n33229) );
  NOR2_X1 U35321 ( .A1(n2699), .A2(n33210), .ZN(n9907) );
  NOR2_X1 U35322 ( .A1(n2698), .A2(n33210), .ZN(n9906) );
  NOR2_X1 U35323 ( .A1(n2697), .A2(n33210), .ZN(n9905) );
  NOR2_X1 U35324 ( .A1(n2696), .A2(n33210), .ZN(n9904) );
  NOR2_X1 U35325 ( .A1(n27871), .A2(n33224), .ZN(n9900) );
  NOR2_X1 U35326 ( .A1(n27874), .A2(n33224), .ZN(n9898) );
  NOR2_X1 U35327 ( .A1(n32082), .A2(RESET), .ZN(n33230) );
  INV_X1 U35328 ( .A(n33227), .ZN(n32082) );
  OAI21_X1 U35329 ( .B1(n33231), .B2(n32148), .A(n41370), .ZN(n33424) );
  INV_X1 U35330 ( .A(RD1), .ZN(n32148) );
  OAI21_X1 U35331 ( .B1(n33231), .B2(n32149), .A(n41370), .ZN(n34698) );
  INV_X1 U35332 ( .A(RD2), .ZN(n32149) );
  NOR2_X1 U35333 ( .A1(ENABLE), .A2(RESET), .ZN(n33231) );
  NAND2_X1 U35334 ( .A1(n41370), .A2(n33219), .ZN(n33212) );
  OAI21_X1 U35335 ( .B1(CALL), .B2(RETRN), .A(ENABLE), .ZN(n33219) );
  NAND2_X1 U35336 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n33208) );
  NAND2_X1 U35337 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n33207) );
  NAND2_X1 U35338 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(n33209) );
  INV_X1 U35339 ( .A(RESET), .ZN(n32079) );
  INV_X1 U35340 ( .A(ENABLE), .ZN(n32081) );
  INV_X1 U35341 ( .A(RETRN), .ZN(n32083) );
  AND2_X1 U35342 ( .A1(WR), .A2(n41370), .ZN(n33300) );
  AND2_X1 U35343 ( .A1(WR), .A2(ENABLE), .ZN(n33299) );
  INV_X1 U35344 ( .A(BUSin[23]), .ZN(n32124) );
  INV_X1 U35345 ( .A(DATAIN[23]), .ZN(n32214) );
  INV_X1 U35346 ( .A(BUSin[24]), .ZN(n32123) );
  INV_X1 U35347 ( .A(DATAIN[24]), .ZN(n32213) );
  INV_X1 U35348 ( .A(BUSin[25]), .ZN(n32122) );
  INV_X1 U35349 ( .A(DATAIN[25]), .ZN(n32212) );
  INV_X1 U35350 ( .A(BUSin[26]), .ZN(n32121) );
  INV_X1 U35351 ( .A(DATAIN[26]), .ZN(n32211) );
  INV_X1 U35352 ( .A(BUSin[27]), .ZN(n32120) );
  INV_X1 U35353 ( .A(DATAIN[27]), .ZN(n32210) );
  INV_X1 U35354 ( .A(BUSin[28]), .ZN(n32119) );
  INV_X1 U35355 ( .A(DATAIN[28]), .ZN(n32209) );
  INV_X1 U35356 ( .A(BUSin[29]), .ZN(n32118) );
  INV_X1 U35357 ( .A(DATAIN[29]), .ZN(n32208) );
  INV_X1 U35358 ( .A(BUSin[30]), .ZN(n32117) );
  INV_X1 U35359 ( .A(DATAIN[30]), .ZN(n32207) );
  INV_X1 U35360 ( .A(BUSin[31]), .ZN(n32116) );
  INV_X1 U35361 ( .A(DATAIN[31]), .ZN(n32206) );
  INV_X1 U35362 ( .A(BUSin[32]), .ZN(n32115) );
  INV_X1 U35363 ( .A(DATAIN[32]), .ZN(n32205) );
  INV_X1 U35364 ( .A(BUSin[33]), .ZN(n32114) );
  INV_X1 U35365 ( .A(DATAIN[33]), .ZN(n32204) );
  INV_X1 U35366 ( .A(BUSin[34]), .ZN(n32113) );
  INV_X1 U35367 ( .A(DATAIN[34]), .ZN(n32203) );
  INV_X1 U35368 ( .A(BUSin[35]), .ZN(n32112) );
  INV_X1 U35369 ( .A(DATAIN[35]), .ZN(n32202) );
  INV_X1 U35370 ( .A(BUSin[36]), .ZN(n32111) );
  INV_X1 U35371 ( .A(DATAIN[36]), .ZN(n32201) );
  INV_X1 U35372 ( .A(BUSin[37]), .ZN(n32110) );
  INV_X1 U35373 ( .A(DATAIN[37]), .ZN(n32200) );
  INV_X1 U35374 ( .A(BUSin[38]), .ZN(n32109) );
  INV_X1 U35375 ( .A(DATAIN[38]), .ZN(n32199) );
  INV_X1 U35376 ( .A(BUSin[39]), .ZN(n32108) );
  INV_X1 U35377 ( .A(DATAIN[39]), .ZN(n32198) );
  INV_X1 U35378 ( .A(BUSin[40]), .ZN(n32107) );
  INV_X1 U35379 ( .A(DATAIN[40]), .ZN(n32197) );
  INV_X1 U35380 ( .A(BUSin[41]), .ZN(n32106) );
  INV_X1 U35381 ( .A(DATAIN[41]), .ZN(n32196) );
  INV_X1 U35382 ( .A(BUSin[42]), .ZN(n32105) );
  INV_X1 U35383 ( .A(DATAIN[42]), .ZN(n32195) );
  INV_X1 U35384 ( .A(BUSin[43]), .ZN(n32104) );
  INV_X1 U35385 ( .A(DATAIN[43]), .ZN(n32194) );
  INV_X1 U35386 ( .A(BUSin[44]), .ZN(n32103) );
  INV_X1 U35387 ( .A(DATAIN[44]), .ZN(n32193) );
  INV_X1 U35388 ( .A(BUSin[45]), .ZN(n32102) );
  INV_X1 U35389 ( .A(DATAIN[45]), .ZN(n32192) );
  INV_X1 U35390 ( .A(BUSin[46]), .ZN(n32101) );
  INV_X1 U35391 ( .A(DATAIN[46]), .ZN(n32191) );
  INV_X1 U35392 ( .A(BUSin[47]), .ZN(n32100) );
  INV_X1 U35393 ( .A(DATAIN[47]), .ZN(n32190) );
  INV_X1 U35394 ( .A(BUSin[48]), .ZN(n32099) );
  INV_X1 U35395 ( .A(DATAIN[48]), .ZN(n32189) );
  INV_X1 U35396 ( .A(BUSin[49]), .ZN(n32098) );
  INV_X1 U35397 ( .A(DATAIN[49]), .ZN(n32188) );
  INV_X1 U35398 ( .A(BUSin[50]), .ZN(n32097) );
  INV_X1 U35399 ( .A(DATAIN[50]), .ZN(n32187) );
  INV_X1 U35400 ( .A(BUSin[51]), .ZN(n32096) );
  INV_X1 U35401 ( .A(DATAIN[51]), .ZN(n32186) );
  INV_X1 U35402 ( .A(BUSin[52]), .ZN(n32095) );
  INV_X1 U35403 ( .A(DATAIN[52]), .ZN(n32185) );
  INV_X1 U35404 ( .A(BUSin[53]), .ZN(n32094) );
  INV_X1 U35405 ( .A(DATAIN[53]), .ZN(n32184) );
  INV_X1 U35406 ( .A(BUSin[54]), .ZN(n32093) );
  INV_X1 U35407 ( .A(DATAIN[54]), .ZN(n32183) );
  INV_X1 U35408 ( .A(BUSin[55]), .ZN(n32092) );
  INV_X1 U35409 ( .A(DATAIN[55]), .ZN(n32182) );
  INV_X1 U35410 ( .A(BUSin[56]), .ZN(n32091) );
  INV_X1 U35411 ( .A(DATAIN[56]), .ZN(n32181) );
  INV_X1 U35412 ( .A(BUSin[57]), .ZN(n32090) );
  INV_X1 U35413 ( .A(DATAIN[57]), .ZN(n32180) );
  INV_X1 U35414 ( .A(BUSin[58]), .ZN(n32089) );
  INV_X1 U35415 ( .A(DATAIN[58]), .ZN(n32179) );
  INV_X1 U35416 ( .A(BUSin[59]), .ZN(n32088) );
  INV_X1 U35417 ( .A(DATAIN[59]), .ZN(n32178) );
  INV_X1 U35418 ( .A(BUSin[60]), .ZN(n32087) );
  INV_X1 U35419 ( .A(DATAIN[60]), .ZN(n32177) );
  INV_X1 U35420 ( .A(BUSin[61]), .ZN(n32086) );
  INV_X1 U35421 ( .A(DATAIN[61]), .ZN(n32176) );
  INV_X1 U35422 ( .A(BUSin[62]), .ZN(n32085) );
  INV_X1 U35423 ( .A(DATAIN[62]), .ZN(n32175) );
  INV_X1 U35424 ( .A(BUSin[63]), .ZN(n32084) );
  INV_X1 U35425 ( .A(DATAIN[63]), .ZN(n32174) );
  INV_X1 U35426 ( .A(BUSin[0]), .ZN(n32147) );
  INV_X1 U35427 ( .A(DATAIN[0]), .ZN(n32237) );
  INV_X1 U35428 ( .A(BUSin[1]), .ZN(n32146) );
  INV_X1 U35429 ( .A(DATAIN[1]), .ZN(n32236) );
  INV_X1 U35430 ( .A(BUSin[2]), .ZN(n32145) );
  INV_X1 U35431 ( .A(DATAIN[2]), .ZN(n32235) );
  INV_X1 U35432 ( .A(BUSin[3]), .ZN(n32144) );
  INV_X1 U35433 ( .A(DATAIN[3]), .ZN(n32234) );
  INV_X1 U35434 ( .A(BUSin[4]), .ZN(n32143) );
  INV_X1 U35435 ( .A(DATAIN[4]), .ZN(n32233) );
  INV_X1 U35436 ( .A(BUSin[5]), .ZN(n32142) );
  INV_X1 U35437 ( .A(DATAIN[5]), .ZN(n32232) );
  INV_X1 U35438 ( .A(BUSin[6]), .ZN(n32141) );
  INV_X1 U35439 ( .A(DATAIN[6]), .ZN(n32231) );
  INV_X1 U35440 ( .A(BUSin[7]), .ZN(n32140) );
  INV_X1 U35441 ( .A(DATAIN[7]), .ZN(n32230) );
  INV_X1 U35442 ( .A(BUSin[8]), .ZN(n32139) );
  INV_X1 U35443 ( .A(DATAIN[8]), .ZN(n32229) );
  INV_X1 U35444 ( .A(BUSin[9]), .ZN(n32138) );
  INV_X1 U35445 ( .A(DATAIN[9]), .ZN(n32228) );
  INV_X1 U35446 ( .A(BUSin[10]), .ZN(n32137) );
  INV_X1 U35447 ( .A(DATAIN[10]), .ZN(n32227) );
  INV_X1 U35448 ( .A(BUSin[11]), .ZN(n32136) );
  INV_X1 U35449 ( .A(DATAIN[11]), .ZN(n32226) );
  INV_X1 U35450 ( .A(BUSin[12]), .ZN(n32135) );
  INV_X1 U35451 ( .A(DATAIN[12]), .ZN(n32225) );
  INV_X1 U35452 ( .A(BUSin[13]), .ZN(n32134) );
  INV_X1 U35453 ( .A(DATAIN[13]), .ZN(n32224) );
  INV_X1 U35454 ( .A(BUSin[14]), .ZN(n32133) );
  INV_X1 U35455 ( .A(DATAIN[14]), .ZN(n32223) );
  INV_X1 U35456 ( .A(BUSin[15]), .ZN(n32132) );
  INV_X1 U35457 ( .A(DATAIN[15]), .ZN(n32222) );
  INV_X1 U35458 ( .A(BUSin[16]), .ZN(n32131) );
  INV_X1 U35459 ( .A(DATAIN[16]), .ZN(n32221) );
  INV_X1 U35460 ( .A(BUSin[17]), .ZN(n32130) );
  INV_X1 U35461 ( .A(DATAIN[17]), .ZN(n32220) );
  INV_X1 U35462 ( .A(BUSin[18]), .ZN(n32129) );
  INV_X1 U35463 ( .A(DATAIN[18]), .ZN(n32219) );
  INV_X1 U35464 ( .A(BUSin[19]), .ZN(n32128) );
  INV_X1 U35465 ( .A(DATAIN[19]), .ZN(n32218) );
  INV_X1 U35466 ( .A(BUSin[20]), .ZN(n32127) );
  INV_X1 U35467 ( .A(DATAIN[20]), .ZN(n32217) );
  INV_X1 U35468 ( .A(BUSin[21]), .ZN(n32126) );
  INV_X1 U35469 ( .A(DATAIN[21]), .ZN(n32216) );
  INV_X1 U35470 ( .A(BUSin[22]), .ZN(n32125) );
  INV_X1 U35471 ( .A(DATAIN[22]), .ZN(n32215) );
  CLKBUF_X1 U35472 ( .A(n36039), .Z(n39053) );
  CLKBUF_X1 U35473 ( .A(n36038), .Z(n39059) );
  CLKBUF_X1 U35474 ( .A(n36037), .Z(n39065) );
  CLKBUF_X1 U35475 ( .A(n36035), .Z(n39071) );
  CLKBUF_X1 U35476 ( .A(n36034), .Z(n39077) );
  CLKBUF_X1 U35477 ( .A(n36033), .Z(n39083) );
  CLKBUF_X1 U35478 ( .A(n36032), .Z(n39089) );
  CLKBUF_X1 U35479 ( .A(n36031), .Z(n39095) );
  CLKBUF_X1 U35480 ( .A(n36029), .Z(n39101) );
  CLKBUF_X1 U35481 ( .A(n36028), .Z(n39107) );
  CLKBUF_X1 U35482 ( .A(n36027), .Z(n39113) );
  CLKBUF_X1 U35483 ( .A(n36026), .Z(n39119) );
  CLKBUF_X1 U35484 ( .A(n36025), .Z(n39125) );
  CLKBUF_X1 U35485 ( .A(n36023), .Z(n39131) );
  CLKBUF_X1 U35486 ( .A(n36022), .Z(n39137) );
  CLKBUF_X1 U35487 ( .A(n36021), .Z(n39143) );
  CLKBUF_X1 U35488 ( .A(n36020), .Z(n39149) );
  CLKBUF_X1 U35489 ( .A(n36019), .Z(n39155) );
  CLKBUF_X1 U35490 ( .A(n36017), .Z(n39161) );
  CLKBUF_X1 U35491 ( .A(n36016), .Z(n39167) );
  CLKBUF_X1 U35492 ( .A(n36011), .Z(n39173) );
  CLKBUF_X1 U35493 ( .A(n36010), .Z(n39179) );
  CLKBUF_X1 U35494 ( .A(n36009), .Z(n39185) );
  CLKBUF_X1 U35495 ( .A(n36007), .Z(n39191) );
  CLKBUF_X1 U35496 ( .A(n36006), .Z(n39197) );
  CLKBUF_X1 U35497 ( .A(n36005), .Z(n39203) );
  CLKBUF_X1 U35498 ( .A(n36004), .Z(n39209) );
  CLKBUF_X1 U35499 ( .A(n36003), .Z(n39215) );
  CLKBUF_X1 U35500 ( .A(n36001), .Z(n39221) );
  CLKBUF_X1 U35501 ( .A(n36000), .Z(n39227) );
  CLKBUF_X1 U35502 ( .A(n35999), .Z(n39233) );
  CLKBUF_X1 U35503 ( .A(n35998), .Z(n39239) );
  CLKBUF_X1 U35504 ( .A(n35997), .Z(n39245) );
  CLKBUF_X1 U35505 ( .A(n35995), .Z(n39251) );
  CLKBUF_X1 U35506 ( .A(n35994), .Z(n39257) );
  CLKBUF_X1 U35507 ( .A(n35993), .Z(n39263) );
  CLKBUF_X1 U35508 ( .A(n35992), .Z(n39269) );
  CLKBUF_X1 U35509 ( .A(n35991), .Z(n39275) );
  CLKBUF_X1 U35510 ( .A(n35989), .Z(n39281) );
  CLKBUF_X1 U35511 ( .A(n35988), .Z(n39287) );
  CLKBUF_X1 U35512 ( .A(n35981), .Z(n39293) );
  CLKBUF_X1 U35513 ( .A(n34758), .Z(n39303) );
  CLKBUF_X1 U35514 ( .A(n34757), .Z(n39309) );
  CLKBUF_X1 U35515 ( .A(n34756), .Z(n39315) );
  CLKBUF_X1 U35516 ( .A(n34754), .Z(n39321) );
  CLKBUF_X1 U35517 ( .A(n34753), .Z(n39327) );
  CLKBUF_X1 U35518 ( .A(n34752), .Z(n39333) );
  CLKBUF_X1 U35519 ( .A(n34751), .Z(n39339) );
  CLKBUF_X1 U35520 ( .A(n34750), .Z(n39345) );
  CLKBUF_X1 U35521 ( .A(n34748), .Z(n39351) );
  CLKBUF_X1 U35522 ( .A(n34747), .Z(n39357) );
  CLKBUF_X1 U35523 ( .A(n34746), .Z(n39363) );
  CLKBUF_X1 U35524 ( .A(n34745), .Z(n39369) );
  CLKBUF_X1 U35525 ( .A(n34744), .Z(n39375) );
  CLKBUF_X1 U35526 ( .A(n34742), .Z(n39381) );
  CLKBUF_X1 U35527 ( .A(n34741), .Z(n39387) );
  CLKBUF_X1 U35528 ( .A(n34740), .Z(n39393) );
  CLKBUF_X1 U35529 ( .A(n34739), .Z(n39399) );
  CLKBUF_X1 U35530 ( .A(n34738), .Z(n39405) );
  CLKBUF_X1 U35531 ( .A(n34736), .Z(n39411) );
  CLKBUF_X1 U35532 ( .A(n34735), .Z(n39417) );
  CLKBUF_X1 U35533 ( .A(n34730), .Z(n39423) );
  CLKBUF_X1 U35534 ( .A(n34729), .Z(n39429) );
  CLKBUF_X1 U35535 ( .A(n34728), .Z(n39435) );
  CLKBUF_X1 U35536 ( .A(n34726), .Z(n39441) );
  CLKBUF_X1 U35537 ( .A(n34725), .Z(n39447) );
  CLKBUF_X1 U35538 ( .A(n34724), .Z(n39453) );
  CLKBUF_X1 U35539 ( .A(n34723), .Z(n39459) );
  CLKBUF_X1 U35540 ( .A(n34722), .Z(n39465) );
  CLKBUF_X1 U35541 ( .A(n34720), .Z(n39471) );
  CLKBUF_X1 U35542 ( .A(n34719), .Z(n39477) );
  CLKBUF_X1 U35543 ( .A(n34718), .Z(n39483) );
  CLKBUF_X1 U35544 ( .A(n34717), .Z(n39489) );
  CLKBUF_X1 U35545 ( .A(n34716), .Z(n39495) );
  CLKBUF_X1 U35546 ( .A(n34714), .Z(n39501) );
  CLKBUF_X1 U35547 ( .A(n34713), .Z(n39507) );
  CLKBUF_X1 U35548 ( .A(n34712), .Z(n39513) );
  CLKBUF_X1 U35549 ( .A(n34711), .Z(n39519) );
  CLKBUF_X1 U35550 ( .A(n34710), .Z(n39525) );
  CLKBUF_X1 U35551 ( .A(n34708), .Z(n39531) );
  CLKBUF_X1 U35552 ( .A(n34707), .Z(n39537) );
  CLKBUF_X1 U35553 ( .A(n34700), .Z(n39543) );
  CLKBUF_X1 U35554 ( .A(n34698), .Z(n39549) );
  CLKBUF_X1 U35555 ( .A(n33484), .Z(n39555) );
  CLKBUF_X1 U35556 ( .A(n33483), .Z(n39561) );
  CLKBUF_X1 U35557 ( .A(n33482), .Z(n39567) );
  CLKBUF_X1 U35558 ( .A(n33480), .Z(n39573) );
  CLKBUF_X1 U35559 ( .A(n33479), .Z(n39579) );
  CLKBUF_X1 U35560 ( .A(n33478), .Z(n39585) );
  CLKBUF_X1 U35561 ( .A(n33477), .Z(n39591) );
  CLKBUF_X1 U35562 ( .A(n33476), .Z(n39597) );
  CLKBUF_X1 U35563 ( .A(n33474), .Z(n39603) );
  CLKBUF_X1 U35564 ( .A(n33473), .Z(n39609) );
  CLKBUF_X1 U35565 ( .A(n33472), .Z(n39615) );
  CLKBUF_X1 U35566 ( .A(n33471), .Z(n39621) );
  CLKBUF_X1 U35567 ( .A(n33470), .Z(n39627) );
  CLKBUF_X1 U35568 ( .A(n33468), .Z(n39633) );
  CLKBUF_X1 U35569 ( .A(n33467), .Z(n39639) );
  CLKBUF_X1 U35570 ( .A(n33466), .Z(n39645) );
  CLKBUF_X1 U35571 ( .A(n33465), .Z(n39651) );
  CLKBUF_X1 U35572 ( .A(n33464), .Z(n39657) );
  CLKBUF_X1 U35573 ( .A(n33462), .Z(n39663) );
  CLKBUF_X1 U35574 ( .A(n33461), .Z(n39669) );
  CLKBUF_X1 U35575 ( .A(n33456), .Z(n39675) );
  CLKBUF_X1 U35576 ( .A(n33455), .Z(n39681) );
  CLKBUF_X1 U35577 ( .A(n33454), .Z(n39687) );
  CLKBUF_X1 U35578 ( .A(n33452), .Z(n39693) );
  CLKBUF_X1 U35579 ( .A(n33451), .Z(n39699) );
  CLKBUF_X1 U35580 ( .A(n33450), .Z(n39705) );
  CLKBUF_X1 U35581 ( .A(n33449), .Z(n39711) );
  CLKBUF_X1 U35582 ( .A(n33448), .Z(n39717) );
  CLKBUF_X1 U35583 ( .A(n33446), .Z(n39723) );
  CLKBUF_X1 U35584 ( .A(n33445), .Z(n39729) );
  CLKBUF_X1 U35585 ( .A(n33444), .Z(n39735) );
  CLKBUF_X1 U35586 ( .A(n33443), .Z(n39741) );
  CLKBUF_X1 U35587 ( .A(n33442), .Z(n39747) );
  CLKBUF_X1 U35588 ( .A(n33440), .Z(n39753) );
  CLKBUF_X1 U35589 ( .A(n33439), .Z(n39759) );
  CLKBUF_X1 U35590 ( .A(n33438), .Z(n39765) );
  CLKBUF_X1 U35591 ( .A(n33437), .Z(n39771) );
  CLKBUF_X1 U35592 ( .A(n33436), .Z(n39777) );
  CLKBUF_X1 U35593 ( .A(n33434), .Z(n39783) );
  CLKBUF_X1 U35594 ( .A(n33433), .Z(n39789) );
  CLKBUF_X1 U35595 ( .A(n33426), .Z(n39795) );
  CLKBUF_X1 U35596 ( .A(n33424), .Z(n39801) );
  CLKBUF_X1 U35597 ( .A(n39807), .Z(n39813) );
  CLKBUF_X1 U35598 ( .A(n39814), .Z(n39820) );
  CLKBUF_X1 U35599 ( .A(n33417), .Z(n39826) );
  CLKBUF_X1 U35600 ( .A(n39827), .Z(n39833) );
  CLKBUF_X1 U35601 ( .A(n39834), .Z(n39840) );
  CLKBUF_X1 U35602 ( .A(n33414), .Z(n39846) );
  CLKBUF_X1 U35603 ( .A(n39847), .Z(n39853) );
  CLKBUF_X1 U35604 ( .A(n39854), .Z(n39860) );
  CLKBUF_X1 U35605 ( .A(n33411), .Z(n39866) );
  CLKBUF_X1 U35606 ( .A(n39867), .Z(n39873) );
  CLKBUF_X1 U35607 ( .A(n39874), .Z(n39880) );
  CLKBUF_X1 U35608 ( .A(n33408), .Z(n39886) );
  CLKBUF_X1 U35609 ( .A(n39887), .Z(n39893) );
  CLKBUF_X1 U35610 ( .A(n39894), .Z(n39900) );
  CLKBUF_X1 U35611 ( .A(n39906), .Z(n39912) );
  CLKBUF_X1 U35612 ( .A(n39913), .Z(n39919) );
  CLKBUF_X1 U35613 ( .A(n39925), .Z(n39931) );
  CLKBUF_X1 U35614 ( .A(n39932), .Z(n39938) );
  CLKBUF_X1 U35615 ( .A(n33393), .Z(n39944) );
  CLKBUF_X1 U35616 ( .A(n39945), .Z(n39951) );
  CLKBUF_X1 U35617 ( .A(n39952), .Z(n39958) );
  CLKBUF_X1 U35618 ( .A(n33390), .Z(n39964) );
  CLKBUF_X1 U35619 ( .A(n39965), .Z(n39971) );
  CLKBUF_X1 U35620 ( .A(n39972), .Z(n39978) );
  CLKBUF_X1 U35621 ( .A(n33387), .Z(n39984) );
  CLKBUF_X1 U35622 ( .A(n39985), .Z(n39991) );
  CLKBUF_X1 U35623 ( .A(n39992), .Z(n39998) );
  CLKBUF_X1 U35624 ( .A(n40004), .Z(n40010) );
  CLKBUF_X1 U35625 ( .A(n40011), .Z(n40017) );
  CLKBUF_X1 U35626 ( .A(n40023), .Z(n40029) );
  CLKBUF_X1 U35627 ( .A(n40030), .Z(n40036) );
  CLKBUF_X1 U35628 ( .A(n33378), .Z(n40042) );
  CLKBUF_X1 U35629 ( .A(n40043), .Z(n40049) );
  CLKBUF_X1 U35630 ( .A(n40050), .Z(n40056) );
  CLKBUF_X1 U35631 ( .A(n33375), .Z(n40062) );
  CLKBUF_X1 U35632 ( .A(n40063), .Z(n40069) );
  CLKBUF_X1 U35633 ( .A(n40070), .Z(n40076) );
  CLKBUF_X1 U35634 ( .A(n33372), .Z(n40082) );
  CLKBUF_X1 U35635 ( .A(n40083), .Z(n40089) );
  CLKBUF_X1 U35636 ( .A(n40090), .Z(n40096) );
  CLKBUF_X1 U35637 ( .A(n40102), .Z(n40108) );
  CLKBUF_X1 U35638 ( .A(n40109), .Z(n40115) );
  CLKBUF_X1 U35639 ( .A(n33361), .Z(n40121) );
  CLKBUF_X1 U35640 ( .A(n40122), .Z(n40128) );
  CLKBUF_X1 U35641 ( .A(n40129), .Z(n40135) );
  CLKBUF_X1 U35642 ( .A(n33358), .Z(n40141) );
  CLKBUF_X1 U35643 ( .A(n40142), .Z(n40148) );
  CLKBUF_X1 U35644 ( .A(n40149), .Z(n40155) );
  CLKBUF_X1 U35645 ( .A(n33355), .Z(n40161) );
  CLKBUF_X1 U35646 ( .A(n40162), .Z(n40168) );
  CLKBUF_X1 U35647 ( .A(n40169), .Z(n40175) );
  CLKBUF_X1 U35648 ( .A(n33352), .Z(n40181) );
  CLKBUF_X1 U35649 ( .A(n40182), .Z(n40188) );
  CLKBUF_X1 U35650 ( .A(n40189), .Z(n40195) );
  CLKBUF_X1 U35651 ( .A(n33349), .Z(n40201) );
  CLKBUF_X1 U35652 ( .A(n40202), .Z(n40208) );
  CLKBUF_X1 U35653 ( .A(n40209), .Z(n40215) );
  CLKBUF_X1 U35654 ( .A(n33346), .Z(n40221) );
  CLKBUF_X1 U35655 ( .A(n40222), .Z(n40228) );
  CLKBUF_X1 U35656 ( .A(n40229), .Z(n40235) );
  CLKBUF_X1 U35657 ( .A(n33343), .Z(n40241) );
  CLKBUF_X1 U35658 ( .A(n40242), .Z(n40248) );
  CLKBUF_X1 U35659 ( .A(n40249), .Z(n40255) );
  CLKBUF_X1 U35660 ( .A(n33336), .Z(n40261) );
  CLKBUF_X1 U35661 ( .A(n40262), .Z(n40268) );
  CLKBUF_X1 U35662 ( .A(n40269), .Z(n40275) );
  CLKBUF_X1 U35663 ( .A(n33329), .Z(n40281) );
  CLKBUF_X1 U35664 ( .A(n40282), .Z(n40288) );
  CLKBUF_X1 U35665 ( .A(n40289), .Z(n40295) );
  CLKBUF_X1 U35666 ( .A(n33326), .Z(n40301) );
  CLKBUF_X1 U35667 ( .A(n40302), .Z(n40308) );
  CLKBUF_X1 U35668 ( .A(n40309), .Z(n40315) );
  CLKBUF_X1 U35669 ( .A(n33323), .Z(n40321) );
  CLKBUF_X1 U35670 ( .A(n40322), .Z(n40328) );
  CLKBUF_X1 U35671 ( .A(n40329), .Z(n40335) );
  CLKBUF_X1 U35672 ( .A(n33320), .Z(n40341) );
  CLKBUF_X1 U35673 ( .A(n40342), .Z(n40348) );
  CLKBUF_X1 U35674 ( .A(n40349), .Z(n40355) );
  CLKBUF_X1 U35675 ( .A(n33317), .Z(n40361) );
  CLKBUF_X1 U35676 ( .A(n40362), .Z(n40368) );
  CLKBUF_X1 U35677 ( .A(n40369), .Z(n40375) );
  CLKBUF_X1 U35678 ( .A(n33314), .Z(n40381) );
  CLKBUF_X1 U35679 ( .A(n40382), .Z(n40388) );
  CLKBUF_X1 U35680 ( .A(n40389), .Z(n40395) );
  CLKBUF_X1 U35681 ( .A(n33311), .Z(n40401) );
  CLKBUF_X1 U35682 ( .A(n40402), .Z(n40408) );
  CLKBUF_X1 U35683 ( .A(n40409), .Z(n40415) );
  CLKBUF_X1 U35684 ( .A(n33304), .Z(n40421) );
  CLKBUF_X1 U35685 ( .A(n40422), .Z(n40428) );
  CLKBUF_X1 U35686 ( .A(n40429), .Z(n40435) );
  CLKBUF_X1 U35687 ( .A(n33293), .Z(n40441) );
  CLKBUF_X1 U35688 ( .A(n40442), .Z(n40448) );
  CLKBUF_X1 U35689 ( .A(n40449), .Z(n40455) );
  CLKBUF_X1 U35690 ( .A(n33288), .Z(n40461) );
  CLKBUF_X1 U35691 ( .A(n40462), .Z(n40468) );
  CLKBUF_X1 U35692 ( .A(n40469), .Z(n40475) );
  CLKBUF_X1 U35693 ( .A(n33283), .Z(n40481) );
  CLKBUF_X1 U35694 ( .A(n40482), .Z(n40488) );
  CLKBUF_X1 U35695 ( .A(n40489), .Z(n40495) );
  CLKBUF_X1 U35696 ( .A(n33278), .Z(n40501) );
  CLKBUF_X1 U35697 ( .A(n40502), .Z(n40508) );
  CLKBUF_X1 U35698 ( .A(n40509), .Z(n40515) );
  CLKBUF_X1 U35699 ( .A(n33273), .Z(n40521) );
  CLKBUF_X1 U35700 ( .A(n40522), .Z(n40528) );
  CLKBUF_X1 U35701 ( .A(n40529), .Z(n40535) );
  CLKBUF_X1 U35702 ( .A(n33268), .Z(n40541) );
  CLKBUF_X1 U35703 ( .A(n40542), .Z(n40548) );
  CLKBUF_X1 U35704 ( .A(n40549), .Z(n40555) );
  CLKBUF_X1 U35705 ( .A(n33263), .Z(n40561) );
  CLKBUF_X1 U35706 ( .A(n40562), .Z(n40568) );
  CLKBUF_X1 U35707 ( .A(n40569), .Z(n40575) );
  CLKBUF_X1 U35708 ( .A(n33254), .Z(n40581) );
  CLKBUF_X1 U35709 ( .A(n40582), .Z(n40588) );
  CLKBUF_X1 U35710 ( .A(n40589), .Z(n40595) );
endmodule

