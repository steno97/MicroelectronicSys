
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type matrix_mux is array (INTEGER range <>) of std_logic_vector (63 downto 0);
type matrix_out_shifter is array (1 downto 0) of std_logic_vector (63 downto 0)
   ;

end CONV_PACK_BOOTHMUL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_15 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_15;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_15 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, net15667, net15665, net15663, net15661, net15659, net15657, 
      net16563, net16581, net16579, net16577, net16575, net16597, net16593, 
      net16591, net16589, net16587, net16609, net16607, net16605, net16603, 
      net16601, net16599, net18142, net18141, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284 : 
      std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => net16563, Z => n136);
   U2 : INV_X1 port map( A => n149, ZN => net16563);
   U3 : BUF_X2 port map( A => n142, Z => net18142);
   U4 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(32));
   U5 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(48));
   U6 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(50));
   U7 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(38));
   U8 : INV_X1 port map( A => INPUT(253), ZN => n150);
   U9 : AOI21_X1 port map( B1 => n158, B2 => INPUT(125), A => n151, ZN => n146)
                           ;
   U10 : NOR2_X1 port map( A1 => n150, A2 => n143, ZN => n151);
   U11 : NOR2_X1 port map( A1 => n156, A2 => n155, ZN => n153);
   U12 : INV_X1 port map( A => net15657, ZN => n154);
   U13 : AND2_X1 port map( A1 => n156, A2 => n155, ZN => n137);
   U14 : AND2_X1 port map( A1 => n153, A2 => n154, ZN => n138);
   U15 : INV_X1 port map( A => n18, ZN => n152);
   U16 : INV_X1 port map( A => n158, ZN => n139);
   U17 : INV_X1 port map( A => n139, ZN => n140);
   U18 : INV_X1 port map( A => n139, ZN => n141);
   U19 : AND2_X2 port map( A1 => n144, A2 => n147, ZN => n142);
   U20 : AOI21_X1 port map( B1 => n142, B2 => INPUT(189), A => n152, ZN => n145
                           );
   U21 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(58));
   U22 : INV_X1 port map( A => net16575, ZN => n143);
   U23 : BUF_X4 port map( A => n137, Z => net16581);
   U24 : BUF_X1 port map( A => SEL(1), Z => n144);
   U25 : NAND2_X1 port map( A1 => n145, A2 => n146, ZN => Y(61));
   U26 : NAND2_X1 port map( A1 => SEL(2), A2 => n148, ZN => n149);
   U27 : INV_X1 port map( A => n149, ZN => n158);
   U28 : INV_X1 port map( A => SEL(2), ZN => n147);
   U29 : INV_X1 port map( A => n147, ZN => n155);
   U30 : CLKBUF_X1 port map( A => net16597, Z => n157);
   U31 : INV_X1 port map( A => SEL(1), ZN => n148);
   U32 : INV_X1 port map( A => n148, ZN => n156);
   U33 : BUF_X2 port map( A => n142, Z => net18141);
   U34 : AOI222_X1 port map( A1 => INPUT(80), A2 => n141, B1 => INPUT(208), B2 
                           => net16579, C1 => INPUT(144), C2 => n157, ZN => 
                           n173);
   U35 : AOI222_X1 port map( A1 => INPUT(79), A2 => n141, B1 => INPUT(207), B2 
                           => net16581, C1 => INPUT(143), C2 => net18141, ZN =>
                           n171);
   U36 : AOI222_X1 port map( A1 => INPUT(115), A2 => net16563, B1 => INPUT(243)
                           , B2 => net16581, C1 => INPUT(179), C2 => net18141, 
                           ZN => n251);
   U37 : AOI222_X1 port map( A1 => INPUT(116), A2 => n140, B1 => INPUT(244), B2
                           => net16581, C1 => INPUT(180), C2 => net18142, ZN =>
                           n253);
   U38 : AOI222_X1 port map( A1 => INPUT(111), A2 => net16563, B1 => INPUT(239)
                           , B2 => net16581, C1 => INPUT(175), C2 => net16587, 
                           ZN => n241);
   U39 : AOI222_X1 port map( A1 => INPUT(110), A2 => n141, B1 => INPUT(238), B2
                           => net16581, C1 => INPUT(174), C2 => net18142, ZN =>
                           n239);
   U40 : AOI222_X1 port map( A1 => INPUT(109), A2 => n136, B1 => INPUT(237), B2
                           => net16581, C1 => INPUT(173), C2 => net18142, ZN =>
                           n237);
   U41 : AOI222_X1 port map( A1 => INPUT(108), A2 => n141, B1 => INPUT(236), B2
                           => net16581, C1 => INPUT(172), C2 => net18141, ZN =>
                           n235);
   U42 : AOI222_X1 port map( A1 => INPUT(107), A2 => n136, B1 => INPUT(235), B2
                           => net16581, C1 => INPUT(171), C2 => net18142, ZN =>
                           n233);
   U43 : AOI222_X1 port map( A1 => INPUT(106), A2 => n141, B1 => INPUT(234), B2
                           => net16581, C1 => INPUT(170), C2 => net18142, ZN =>
                           n231);
   U44 : AOI222_X1 port map( A1 => INPUT(94), A2 => n141, B1 => INPUT(222), B2 
                           => net16581, C1 => INPUT(158), C2 => net18141, ZN =>
                           n205);
   U45 : AOI222_X1 port map( A1 => INPUT(95), A2 => n136, B1 => INPUT(223), B2 
                           => net16579, C1 => INPUT(159), C2 => net18142, ZN =>
                           n207);
   U46 : AOI222_X1 port map( A1 => INPUT(96), A2 => n141, B1 => INPUT(224), B2 
                           => net16581, C1 => INPUT(160), C2 => net18141, ZN =>
                           n209);
   U47 : AOI222_X1 port map( A1 => INPUT(97), A2 => n136, B1 => INPUT(225), B2 
                           => net16579, C1 => INPUT(161), C2 => net18141, ZN =>
                           n211);
   U48 : AOI222_X1 port map( A1 => INPUT(98), A2 => n141, B1 => INPUT(226), B2 
                           => net16581, C1 => INPUT(162), C2 => net18141, ZN =>
                           n213);
   U49 : AOI222_X1 port map( A1 => INPUT(99), A2 => n136, B1 => INPUT(227), B2 
                           => net16579, C1 => INPUT(163), C2 => net18141, ZN =>
                           n215);
   U50 : AOI222_X1 port map( A1 => INPUT(100), A2 => n141, B1 => INPUT(228), B2
                           => net16581, C1 => INPUT(164), C2 => net16587, ZN =>
                           n217);
   U51 : AOI222_X1 port map( A1 => INPUT(101), A2 => n136, B1 => INPUT(229), B2
                           => net16579, C1 => INPUT(165), C2 => net16591, ZN =>
                           n219);
   U52 : AOI222_X1 port map( A1 => INPUT(105), A2 => n136, B1 => INPUT(233), B2
                           => net16581, C1 => INPUT(169), C2 => net18141, ZN =>
                           n229);
   U53 : AOI222_X1 port map( A1 => INPUT(104), A2 => n141, B1 => INPUT(232), B2
                           => net16581, C1 => INPUT(168), C2 => n157, ZN => 
                           n227);
   U54 : AOI222_X1 port map( A1 => INPUT(103), A2 => n136, B1 => INPUT(231), B2
                           => net16581, C1 => INPUT(167), C2 => net16597, ZN =>
                           n223);
   U55 : AOI222_X1 port map( A1 => INPUT(102), A2 => n141, B1 => INPUT(230), B2
                           => net16579, C1 => INPUT(166), C2 => net16589, ZN =>
                           n221);
   U56 : CLKBUF_X1 port map( A => n142, Z => net16593);
   U57 : CLKBUF_X1 port map( A => n142, Z => net16591);
   U58 : CLKBUF_X1 port map( A => n137, Z => net16579);
   U59 : AOI222_X1 port map( A1 => INPUT(91), A2 => n136, B1 => INPUT(219), B2 
                           => net16581, C1 => INPUT(155), C2 => net16591, ZN =>
                           n197);
   U60 : AOI222_X1 port map( A1 => INPUT(90), A2 => n141, B1 => INPUT(218), B2 
                           => net16579, C1 => INPUT(154), C2 => net16587, ZN =>
                           n195);
   U61 : AOI222_X1 port map( A1 => INPUT(89), A2 => n136, B1 => INPUT(217), B2 
                           => net16581, C1 => INPUT(153), C2 => n157, ZN => 
                           n193);
   U62 : AOI222_X1 port map( A1 => INPUT(87), A2 => n136, B1 => INPUT(215), B2 
                           => net16581, C1 => INPUT(151), C2 => net18141, ZN =>
                           n189);
   U63 : AOI222_X1 port map( A1 => INPUT(86), A2 => n141, B1 => INPUT(214), B2 
                           => net16579, C1 => INPUT(150), C2 => net18142, ZN =>
                           n187);
   U64 : AOI222_X1 port map( A1 => INPUT(85), A2 => n136, B1 => INPUT(213), B2 
                           => net16581, C1 => INPUT(149), C2 => net18141, ZN =>
                           n185);
   U65 : AOI222_X1 port map( A1 => INPUT(88), A2 => n141, B1 => INPUT(216), B2 
                           => net16579, C1 => INPUT(152), C2 => net18142, ZN =>
                           n191);
   U66 : AOI222_X1 port map( A1 => INPUT(92), A2 => n141, B1 => INPUT(220), B2 
                           => net16579, C1 => INPUT(156), C2 => net16589, ZN =>
                           n199);
   U67 : AOI222_X1 port map( A1 => INPUT(84), A2 => n141, B1 => INPUT(212), B2 
                           => net16579, C1 => INPUT(148), C2 => net16597, ZN =>
                           n183);
   U68 : AOI222_X1 port map( A1 => INPUT(93), A2 => n136, B1 => INPUT(221), B2 
                           => net16579, C1 => INPUT(157), C2 => net16597, ZN =>
                           n201);
   U69 : CLKBUF_X1 port map( A => n142, Z => net16589);
   U70 : CLKBUF_X1 port map( A => n137, Z => net16577);
   U71 : AOI222_X1 port map( A1 => INPUT(74), A2 => n141, B1 => INPUT(202), B2 
                           => net16579, C1 => INPUT(138), C2 => net16597, ZN =>
                           n161);
   U72 : AOI222_X1 port map( A1 => INPUT(83), A2 => n136, B1 => INPUT(211), B2 
                           => net16581, C1 => INPUT(147), C2 => net16589, ZN =>
                           n179);
   U73 : AOI222_X1 port map( A1 => INPUT(73), A2 => n136, B1 => INPUT(201), B2 
                           => net16581, C1 => INPUT(137), C2 => net16589, ZN =>
                           n283);
   U74 : AOI222_X1 port map( A1 => INPUT(76), A2 => n141, B1 => INPUT(204), B2 
                           => net16581, C1 => INPUT(140), C2 => net18142, ZN =>
                           n165);
   U75 : AOI222_X1 port map( A1 => INPUT(75), A2 => n136, B1 => INPUT(203), B2 
                           => net16579, C1 => INPUT(139), C2 => net18141, ZN =>
                           n163);
   U76 : AOI222_X1 port map( A1 => INPUT(78), A2 => n141, B1 => INPUT(206), B2 
                           => net16579, C1 => INPUT(142), C2 => net18142, ZN =>
                           n169);
   U77 : AOI222_X1 port map( A1 => INPUT(77), A2 => n136, B1 => INPUT(205), B2 
                           => net16581, C1 => INPUT(141), C2 => net18141, ZN =>
                           n167);
   U78 : AOI222_X1 port map( A1 => INPUT(82), A2 => n136, B1 => INPUT(210), B2 
                           => net16581, C1 => INPUT(146), C2 => net16591, ZN =>
                           n177);
   U79 : AOI222_X1 port map( A1 => INPUT(81), A2 => n136, B1 => INPUT(209), B2 
                           => net16579, C1 => INPUT(145), C2 => net16587, ZN =>
                           n175);
   U80 : CLKBUF_X1 port map( A => n137, Z => net16575);
   U81 : CLKBUF_X1 port map( A => n142, Z => net16587);
   U82 : AOI222_X1 port map( A1 => INPUT(70), A2 => n141, B1 => INPUT(198), B2 
                           => net16581, C1 => INPUT(134), C2 => net18142, ZN =>
                           n277);
   U83 : AOI222_X1 port map( A1 => INPUT(68), A2 => n141, B1 => INPUT(196), B2 
                           => net16579, C1 => INPUT(132), C2 => net16597, ZN =>
                           n247);
   U84 : AOI222_X1 port map( A1 => INPUT(67), A2 => n136, B1 => INPUT(195), B2 
                           => net16581, C1 => INPUT(131), C2 => net16589, ZN =>
                           n225);
   U85 : AOI222_X1 port map( A1 => INPUT(72), A2 => n141, B1 => INPUT(200), B2 
                           => net16579, C1 => INPUT(136), C2 => net16591, ZN =>
                           n281);
   U86 : AOI222_X1 port map( A1 => INPUT(71), A2 => n136, B1 => INPUT(199), B2 
                           => net16581, C1 => INPUT(135), C2 => net16587, ZN =>
                           n279);
   U87 : AOI222_X1 port map( A1 => INPUT(66), A2 => n141, B1 => INPUT(194), B2 
                           => net16581, C1 => INPUT(130), C2 => net16591, ZN =>
                           n203);
   U88 : AOI222_X1 port map( A1 => INPUT(65), A2 => n136, B1 => INPUT(193), B2 
                           => net16579, C1 => INPUT(129), C2 => net16587, ZN =>
                           n181);
   U89 : AOI222_X1 port map( A1 => INPUT(64), A2 => n136, B1 => INPUT(192), B2 
                           => net16581, C1 => INPUT(128), C2 => net18142, ZN =>
                           n159);
   U90 : BUF_X1 port map( A => n138, Z => net16605);
   U91 : BUF_X1 port map( A => n138, Z => net16603);
   U92 : BUF_X1 port map( A => n138, Z => net16601);
   U93 : BUF_X1 port map( A => n138, Z => net16599);
   U94 : CLKBUF_X1 port map( A => n138, Z => net16607);
   U95 : AOI222_X1 port map( A1 => INPUT(114), A2 => n140, B1 => INPUT(242), B2
                           => net16581, C1 => INPUT(178), C2 => net16589, ZN =>
                           n249);
   U96 : BUF_X2 port map( A => SEL(0), Z => net15665);
   U97 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(7));
   U98 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(6));
   U99 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(4));
   U100 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(5));
   U101 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(29));
   U102 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(28));
   U103 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(27));
   U104 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(26));
   U105 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(25));
   U106 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(24));
   U107 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(23));
   U108 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(22));
   U109 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(21));
   U110 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(30));
   U111 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(20));
   U112 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(16));
   U113 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(15));
   U114 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(14));
   U115 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(13));
   U116 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => Y(12));
   U117 : NAND2_X1 port map( A1 => n164, A2 => n163, ZN => Y(11));
   U118 : NAND2_X1 port map( A1 => n162, A2 => n161, ZN => Y(10));
   U119 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(9));
   U120 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(8));
   U121 : AOI222_X1 port map( A1 => INPUT(113), A2 => net16563, B1 => 
                           INPUT(241), B2 => net16581, C1 => INPUT(177), C2 => 
                           n157, ZN => n245);
   U122 : AOI222_X1 port map( A1 => INPUT(112), A2 => n140, B1 => INPUT(240), 
                           B2 => net16581, C1 => INPUT(176), C2 => net16591, ZN
                           => n243);
   U123 : CLKBUF_X1 port map( A => SEL(0), Z => net15663);
   U124 : CLKBUF_X1 port map( A => SEL(0), Z => net15661);
   U125 : CLKBUF_X1 port map( A => SEL(0), Z => net15659);
   U126 : CLKBUF_X1 port map( A => SEL(0), Z => net15657);
   U127 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(3));
   U128 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(2));
   U129 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(1));
   U130 : NAND2_X1 port map( A1 => n160, A2 => n159, ZN => Y(0));
   U131 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(19));
   U132 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(18));
   U133 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(17));
   U134 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(31));
   U135 : AOI22_X1 port map( A1 => INPUT(31), A2 => net16603, B1 => INPUT(287),
                           B2 => net15661, ZN => n208);
   U136 : AOI22_X1 port map( A1 => INPUT(32), A2 => net16603, B1 => INPUT(288),
                           B2 => net15661, ZN => n210);
   U137 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(33));
   U138 : AOI22_X1 port map( A1 => INPUT(33), A2 => net16603, B1 => INPUT(289),
                           B2 => net15661, ZN => n212);
   U139 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(34));
   U140 : AOI22_X1 port map( A1 => INPUT(34), A2 => net16603, B1 => INPUT(290),
                           B2 => net15661, ZN => n214);
   U141 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(35));
   U142 : AOI22_X1 port map( A1 => INPUT(35), A2 => net16603, B1 => INPUT(291),
                           B2 => net15661, ZN => n216);
   U143 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(36));
   U144 : AOI22_X1 port map( A1 => INPUT(36), A2 => net16603, B1 => INPUT(292),
                           B2 => net15661, ZN => n218);
   U145 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(37));
   U146 : AOI22_X1 port map( A1 => INPUT(37), A2 => net16603, B1 => INPUT(293),
                           B2 => net15661, ZN => n220);
   U147 : AOI22_X1 port map( A1 => INPUT(38), A2 => net16603, B1 => INPUT(294),
                           B2 => net15661, ZN => n222);
   U148 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(39));
   U149 : AOI22_X1 port map( A1 => INPUT(39), A2 => net16603, B1 => INPUT(295),
                           B2 => net15661, ZN => n224);
   U150 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(42));
   U151 : AOI22_X1 port map( A1 => INPUT(42), A2 => net16605, B1 => INPUT(298),
                           B2 => net15663, ZN => n232);
   U152 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(41));
   U153 : AOI22_X1 port map( A1 => INPUT(41), A2 => net16603, B1 => INPUT(297),
                           B2 => net15663, ZN => n230);
   U154 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(40));
   U155 : AOI22_X1 port map( A1 => INPUT(40), A2 => net16603, B1 => INPUT(296),
                           B2 => net15661, ZN => n228);
   U156 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(56));
   U157 : AOI22_X1 port map( A1 => INPUT(56), A2 => net16607, B1 => INPUT(312),
                           B2 => net15665, ZN => n262);
   U158 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(55));
   U159 : AOI22_X1 port map( A1 => INPUT(55), A2 => net16607, B1 => INPUT(311),
                           B2 => net15665, ZN => n260);
   U160 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(54));
   U161 : AOI22_X1 port map( A1 => INPUT(54), A2 => net16607, B1 => INPUT(310),
                           B2 => net15665, ZN => n258);
   U162 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(53));
   U163 : AOI22_X1 port map( A1 => INPUT(53), A2 => net16607, B1 => INPUT(309),
                           B2 => net15665, ZN => n256);
   U164 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(52));
   U165 : AOI22_X1 port map( A1 => INPUT(52), A2 => net16605, B1 => INPUT(308),
                           B2 => net15665, ZN => n254);
   U166 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(51));
   U167 : AOI22_X1 port map( A1 => INPUT(51), A2 => net16605, B1 => INPUT(307),
                           B2 => net15663, ZN => n252);
   U168 : AOI22_X1 port map( A1 => INPUT(50), A2 => net16605, B1 => INPUT(306),
                           B2 => net15663, ZN => n250);
   U169 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(49));
   U170 : AOI22_X1 port map( A1 => INPUT(49), A2 => net16605, B1 => INPUT(305),
                           B2 => net15663, ZN => n246);
   U171 : AOI22_X1 port map( A1 => INPUT(48), A2 => net16605, B1 => INPUT(304),
                           B2 => net15663, ZN => n244);
   U172 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(47));
   U173 : AOI22_X1 port map( A1 => INPUT(47), A2 => net16605, B1 => INPUT(303),
                           B2 => net15663, ZN => n242);
   U174 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(46));
   U175 : AOI22_X1 port map( A1 => INPUT(46), A2 => net16605, B1 => INPUT(302),
                           B2 => net15663, ZN => n240);
   U176 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(45));
   U177 : AOI22_X1 port map( A1 => INPUT(45), A2 => net16605, B1 => INPUT(301),
                           B2 => net15663, ZN => n238);
   U178 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(44));
   U179 : AOI22_X1 port map( A1 => INPUT(44), A2 => net16605, B1 => INPUT(300),
                           B2 => net15663, ZN => n236);
   U180 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(43));
   U181 : AOI22_X1 port map( A1 => INPUT(43), A2 => net16605, B1 => INPUT(299),
                           B2 => net15663, ZN => n234);
   U182 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(57));
   U183 : AOI22_X1 port map( A1 => INPUT(57), A2 => net16607, B1 => INPUT(313),
                           B2 => net15665, ZN => n264);
   U184 : AOI22_X1 port map( A1 => INPUT(59), A2 => net16607, B1 => INPUT(315),
                           B2 => net15665, ZN => n268);
   U185 : AOI22_X1 port map( A1 => INPUT(29), A2 => net16601, B1 => INPUT(285),
                           B2 => net15659, ZN => n202);
   U186 : AOI22_X1 port map( A1 => INPUT(30), A2 => net16601, B1 => INPUT(286),
                           B2 => net15661, ZN => n206);
   U187 : AOI22_X1 port map( A1 => INPUT(26), A2 => net16601, B1 => INPUT(282),
                           B2 => net15659, ZN => n196);
   U188 : AOI22_X1 port map( A1 => INPUT(25), A2 => net16601, B1 => INPUT(281),
                           B2 => net15659, ZN => n194);
   U189 : AOI22_X1 port map( A1 => INPUT(24), A2 => net16601, B1 => INPUT(280),
                           B2 => net15659, ZN => n192);
   U190 : AOI22_X1 port map( A1 => INPUT(22), A2 => net16601, B1 => INPUT(278),
                           B2 => net15659, ZN => n188);
   U191 : AOI22_X1 port map( A1 => INPUT(21), A2 => net16601, B1 => INPUT(277),
                           B2 => net15659, ZN => n186);
   U192 : AOI22_X1 port map( A1 => INPUT(20), A2 => net16601, B1 => INPUT(276),
                           B2 => net15659, ZN => n184);
   U193 : AOI22_X1 port map( A1 => INPUT(23), A2 => net16601, B1 => INPUT(279),
                           B2 => net15659, ZN => n190);
   U194 : AOI22_X1 port map( A1 => INPUT(27), A2 => net16601, B1 => INPUT(283),
                           B2 => net15659, ZN => n198);
   U195 : AOI22_X1 port map( A1 => INPUT(28), A2 => net16601, B1 => INPUT(284),
                           B2 => net15659, ZN => n200);
   U196 : AOI22_X1 port map( A1 => INPUT(9), A2 => net16609, B1 => net15667, B2
                           => INPUT(265), ZN => n284);
   U197 : AOI22_X1 port map( A1 => INPUT(18), A2 => net16599, B1 => INPUT(274),
                           B2 => net15657, ZN => n178);
   U198 : AOI22_X1 port map( A1 => INPUT(19), A2 => net16599, B1 => INPUT(275),
                           B2 => net15657, ZN => n180);
   U199 : AOI22_X1 port map( A1 => INPUT(11), A2 => net16599, B1 => INPUT(267),
                           B2 => net15657, ZN => n164);
   U200 : AOI22_X1 port map( A1 => INPUT(10), A2 => net16599, B1 => INPUT(266),
                           B2 => net15657, ZN => n162);
   U201 : AOI22_X1 port map( A1 => INPUT(13), A2 => net16599, B1 => INPUT(269),
                           B2 => net15657, ZN => n168);
   U202 : AOI22_X1 port map( A1 => INPUT(12), A2 => net16599, B1 => INPUT(268),
                           B2 => net15657, ZN => n166);
   U203 : AOI22_X1 port map( A1 => INPUT(15), A2 => net16599, B1 => INPUT(271),
                           B2 => net15657, ZN => n172);
   U204 : AOI22_X1 port map( A1 => INPUT(16), A2 => net16599, B1 => INPUT(272),
                           B2 => net15657, ZN => n174);
   U205 : AOI22_X1 port map( A1 => INPUT(14), A2 => net16599, B1 => INPUT(270),
                           B2 => net15657, ZN => n170);
   U206 : AOI22_X1 port map( A1 => INPUT(17), A2 => net16599, B1 => INPUT(273),
                           B2 => net15657, ZN => n176);
   U207 : AOI22_X1 port map( A1 => INPUT(5), A2 => net16607, B1 => INPUT(261), 
                           B2 => net15665, ZN => n270);
   U208 : AOI22_X1 port map( A1 => INPUT(3), A2 => net16603, B1 => INPUT(259), 
                           B2 => net15661, ZN => n226);
   U209 : AOI22_X1 port map( A1 => INPUT(2), A2 => net16601, B1 => INPUT(258), 
                           B2 => net15659, ZN => n204);
   U210 : AOI22_X1 port map( A1 => INPUT(8), A2 => net16609, B1 => INPUT(264), 
                           B2 => net15667, ZN => n282);
   U211 : AOI22_X1 port map( A1 => INPUT(7), A2 => net16609, B1 => INPUT(263), 
                           B2 => net15667, ZN => n280);
   U212 : AOI22_X1 port map( A1 => INPUT(6), A2 => net16609, B1 => INPUT(262), 
                           B2 => net15667, ZN => n278);
   U213 : AOI22_X1 port map( A1 => INPUT(4), A2 => net16605, B1 => INPUT(260), 
                           B2 => net15663, ZN => n248);
   U214 : AOI22_X1 port map( A1 => INPUT(1), A2 => net16599, B1 => INPUT(257), 
                           B2 => net15659, ZN => n182);
   U215 : AOI22_X1 port map( A1 => INPUT(0), A2 => net16599, B1 => INPUT(256), 
                           B2 => net15657, ZN => n160);
   U216 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(63));
   U217 : AOI22_X1 port map( A1 => INPUT(63), A2 => net16607, B1 => INPUT(319),
                           B2 => net15667, ZN => n276);
   U218 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(62));
   U219 : AOI22_X1 port map( A1 => INPUT(62), A2 => net16607, B1 => INPUT(318),
                           B2 => net15665, ZN => n274);
   U220 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(60));
   U221 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(59));
   U222 : AOI22_X1 port map( A1 => INPUT(61), A2 => net16607, B1 => INPUT(317),
                           B2 => net15665, ZN => n18);
   U223 : AOI222_X1 port map( A1 => INPUT(126), A2 => n141, B1 => INPUT(254), 
                           B2 => net16579, C1 => INPUT(190), C2 => n157, ZN => 
                           n273);
   U224 : AOI222_X1 port map( A1 => INPUT(127), A2 => n141, B1 => INPUT(255), 
                           B2 => net16579, C1 => INPUT(191), C2 => n157, ZN => 
                           n275);
   U225 : AOI222_X1 port map( A1 => INPUT(69), A2 => n136, B1 => INPUT(197), B2
                           => net16579, C1 => INPUT(133), C2 => net18141, ZN =>
                           n269);
   U226 : AOI222_X1 port map( A1 => INPUT(117), A2 => net16563, B1 => 
                           INPUT(245), B2 => net16581, C1 => INPUT(181), C2 => 
                           net18141, ZN => n255);
   U227 : AOI222_X1 port map( A1 => INPUT(118), A2 => n140, B1 => INPUT(246), 
                           B2 => net16581, C1 => INPUT(182), C2 => net16597, ZN
                           => n257);
   U228 : AOI222_X1 port map( A1 => INPUT(119), A2 => net16563, B1 => 
                           INPUT(247), B2 => net16579, C1 => INPUT(183), C2 => 
                           net18141, ZN => n259);
   U229 : AOI222_X1 port map( A1 => INPUT(120), A2 => n140, B1 => INPUT(248), 
                           B2 => net16575, C1 => INPUT(184), C2 => net16587, ZN
                           => n261);
   U230 : AOI222_X1 port map( A1 => INPUT(121), A2 => net16563, B1 => 
                           INPUT(249), B2 => net16577, C1 => INPUT(185), C2 => 
                           net16591, ZN => n263);
   U231 : AOI222_X1 port map( A1 => INPUT(122), A2 => n140, B1 => INPUT(250), 
                           B2 => n137, C1 => INPUT(186), C2 => net16589, ZN => 
                           n265);
   U232 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n137, C1 => INPUT(188), C2 => net16593, ZN => 
                           n271);
   U233 : AOI22_X1 port map( A1 => INPUT(60), A2 => net16607, B1 => INPUT(316),
                           B2 => net15665, ZN => n272);
   U234 : AOI22_X1 port map( A1 => INPUT(58), A2 => net16607, B1 => INPUT(314),
                           B2 => net15665, ZN => n266);
   U235 : AOI222_X1 port map( A1 => INPUT(123), A2 => net16563, B1 => 
                           INPUT(251), B2 => net16577, C1 => INPUT(187), C2 => 
                           net18142, ZN => n267);
   U236 : CLKBUF_X1 port map( A => n138, Z => net16609);
   U237 : CLKBUF_X1 port map( A => n142, Z => net16597);
   U238 : CLKBUF_X1 port map( A => SEL(0), Z => net15667);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_14 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_14;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_14 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U2 : NAND2_X2 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U3 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U4 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U5 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U6 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U7 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U8 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U9 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U10 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U11 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U12 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U13 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U14 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U15 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U16 : BUF_X1 port map( A => n295, Z => n152);
   U17 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U18 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U19 : BUF_X2 port map( A => n296, Z => n158);
   U20 : BUF_X2 port map( A => n294, Z => n146);
   U21 : CLKBUF_X1 port map( A => n296, Z => n157);
   U22 : CLKBUF_X1 port map( A => n296, Z => n156);
   U23 : CLKBUF_X1 port map( A => n294, Z => n145);
   U24 : CLKBUF_X1 port map( A => n294, Z => n144);
   U25 : CLKBUF_X1 port map( A => n296, Z => n155);
   U26 : CLKBUF_X1 port map( A => n294, Z => n143);
   U27 : CLKBUF_X1 port map( A => n296, Z => n154);
   U28 : CLKBUF_X1 port map( A => n294, Z => n142);
   U29 : CLKBUF_X1 port map( A => SEL(0), Z => n163);
   U30 : CLKBUF_X1 port map( A => SEL(0), Z => n162);
   U31 : CLKBUF_X1 port map( A => SEL(0), Z => n161);
   U32 : CLKBUF_X1 port map( A => SEL(0), Z => n160);
   U33 : CLKBUF_X1 port map( A => n295, Z => n151);
   U34 : CLKBUF_X1 port map( A => n295, Z => n150);
   U35 : CLKBUF_X1 port map( A => n295, Z => n149);
   U36 : CLKBUF_X1 port map( A => n295, Z => n148);
   U37 : BUF_X1 port map( A => n293, Z => n139);
   U38 : BUF_X1 port map( A => n293, Z => n138);
   U39 : BUF_X1 port map( A => n293, Z => n137);
   U40 : BUF_X1 port map( A => n293, Z => n136);
   U41 : BUF_X1 port map( A => n293, Z => n140);
   U42 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U43 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U44 : INV_X1 port map( A => SEL(2), ZN => n166);
   U45 : BUF_X1 port map( A => SEL(0), Z => n164);
   U46 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U47 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U48 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U49 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U50 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U51 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U52 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U53 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U54 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U55 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U56 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U57 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U58 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U59 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U60 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U61 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U62 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U63 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U64 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U65 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U66 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U67 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U68 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U69 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U70 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U71 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U72 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U73 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U74 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U75 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U76 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U77 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U78 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U79 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U80 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U81 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U82 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U83 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U84 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U85 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U86 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U87 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U88 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U89 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U90 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U91 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U92 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U93 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2 
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U94 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U95 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U96 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U97 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U98 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U99 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2 
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U100 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U101 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U102 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U103 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U104 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 
                           => n165, ZN => n288);
   U105 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U106 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U107 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U108 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U109 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U110 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U111 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U112 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 
                           => n164, ZN => n278);
   U113 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U114 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U115 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U116 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U117 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 
                           => n163, ZN => n256);
   U118 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U119 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U120 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U121 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U122 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U123 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U124 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U125 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U126 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U127 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U128 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U129 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U130 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U131 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U132 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U133 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U134 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U135 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U136 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U137 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U138 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U139 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U140 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U141 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U142 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U143 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U144 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U145 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U146 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U147 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U148 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U149 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U150 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U151 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U152 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U153 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U154 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U155 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U156 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U157 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U158 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U159 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U160 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U161 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U162 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U163 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U164 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U165 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U166 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U167 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U168 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U169 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U170 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U171 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U172 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U173 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U174 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U175 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U176 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U177 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U178 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U179 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U180 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U181 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U182 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U183 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U184 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U185 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U186 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U187 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U188 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U189 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U190 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U191 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U192 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U193 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 
                           => n162, ZN => n234);
   U194 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U195 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U196 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 
                           => n161, ZN => n212);
   U197 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U198 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U199 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 
                           => n161, ZN => n190);
   U200 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U201 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U202 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U203 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U204 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U205 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U206 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U207 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U208 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U209 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U210 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U211 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U212 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U213 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U214 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U215 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U216 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U217 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U218 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U219 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U220 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U221 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U222 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_13 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_13;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_13 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U2 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U3 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U4 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U5 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U6 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U7 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U8 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U9 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U10 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U11 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U12 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U13 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U14 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U15 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U16 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U17 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U18 : BUF_X1 port map( A => n295, Z => n152);
   U19 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U20 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U21 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U22 : BUF_X2 port map( A => n296, Z => n158);
   U23 : CLKBUF_X1 port map( A => n296, Z => n157);
   U24 : CLKBUF_X1 port map( A => n296, Z => n156);
   U25 : CLKBUF_X1 port map( A => n295, Z => n151);
   U26 : BUF_X2 port map( A => n294, Z => n146);
   U27 : CLKBUF_X1 port map( A => n294, Z => n145);
   U28 : CLKBUF_X1 port map( A => n294, Z => n144);
   U29 : CLKBUF_X1 port map( A => n296, Z => n155);
   U30 : CLKBUF_X1 port map( A => n294, Z => n143);
   U31 : CLKBUF_X1 port map( A => n296, Z => n154);
   U32 : CLKBUF_X1 port map( A => n294, Z => n142);
   U33 : CLKBUF_X1 port map( A => SEL(0), Z => n163);
   U34 : CLKBUF_X1 port map( A => SEL(0), Z => n162);
   U35 : CLKBUF_X1 port map( A => SEL(0), Z => n161);
   U36 : CLKBUF_X1 port map( A => SEL(0), Z => n160);
   U37 : CLKBUF_X1 port map( A => n295, Z => n150);
   U38 : CLKBUF_X1 port map( A => n295, Z => n149);
   U39 : CLKBUF_X1 port map( A => n295, Z => n148);
   U40 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U41 : BUF_X1 port map( A => n293, Z => n139);
   U42 : BUF_X1 port map( A => n293, Z => n138);
   U43 : BUF_X1 port map( A => n293, Z => n137);
   U44 : BUF_X1 port map( A => n293, Z => n136);
   U45 : BUF_X1 port map( A => n293, Z => n140);
   U46 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U47 : BUF_X1 port map( A => SEL(0), Z => n164);
   U48 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U49 : INV_X1 port map( A => SEL(2), ZN => n166);
   U50 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U51 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U52 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U53 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U54 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U55 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U56 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U57 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U58 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U59 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U60 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U61 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U62 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U63 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U64 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U65 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U66 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U67 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U68 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U69 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U70 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U71 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U72 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U73 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U74 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U75 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U76 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U77 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U78 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U79 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U80 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U81 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U82 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U83 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U84 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U85 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U86 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U87 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U88 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U89 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U90 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U91 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U92 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U93 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U94 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U95 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U96 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U97 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U98 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U99 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U100 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U101 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U102 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U103 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 
                           => n165, ZN => n292);
   U104 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U105 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U106 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U107 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U108 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U109 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 
                           => n165, ZN => n290);
   U110 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U111 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U112 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U113 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U114 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U115 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U116 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U117 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U118 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U119 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U120 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U121 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U122 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U123 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U124 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U125 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U126 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U127 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U128 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U129 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U130 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U131 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U132 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U133 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U134 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U135 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U136 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U137 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U138 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U139 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U140 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U141 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U142 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U143 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U144 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U145 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U146 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U147 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U148 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U149 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U150 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U151 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U152 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U153 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U154 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U155 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U156 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U157 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U158 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U159 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U160 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U161 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U162 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U163 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U164 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U165 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U166 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U167 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U168 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U169 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U170 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U171 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U172 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U173 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U174 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U175 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U176 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U177 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U178 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U179 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U180 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U181 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U182 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U183 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U184 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U185 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U186 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U187 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U188 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U189 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U190 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U191 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U192 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U193 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U194 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U195 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U196 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U197 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U198 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U199 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U200 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U201 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U202 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U203 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U204 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U205 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U206 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U207 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U208 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U209 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U210 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U211 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U212 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U213 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U214 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U215 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U216 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U217 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U218 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U219 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U220 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U221 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U222 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_12 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_12;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_12 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U2 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U3 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U4 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U5 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U6 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U7 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U8 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U9 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U10 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U11 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U12 : BUF_X2 port map( A => n296, Z => n158);
   U13 : CLKBUF_X1 port map( A => n296, Z => n157);
   U14 : CLKBUF_X1 port map( A => n296, Z => n156);
   U15 : BUF_X2 port map( A => n294, Z => n146);
   U16 : CLKBUF_X1 port map( A => n294, Z => n145);
   U17 : CLKBUF_X1 port map( A => n294, Z => n144);
   U18 : CLKBUF_X1 port map( A => n296, Z => n155);
   U19 : CLKBUF_X1 port map( A => n294, Z => n143);
   U20 : CLKBUF_X1 port map( A => n296, Z => n154);
   U21 : CLKBUF_X1 port map( A => n294, Z => n142);
   U22 : CLKBUF_X1 port map( A => SEL(0), Z => n163);
   U23 : CLKBUF_X1 port map( A => SEL(0), Z => n162);
   U24 : CLKBUF_X1 port map( A => SEL(0), Z => n161);
   U25 : CLKBUF_X1 port map( A => SEL(0), Z => n160);
   U26 : BUF_X1 port map( A => n295, Z => n151);
   U27 : BUF_X2 port map( A => n295, Z => n152);
   U28 : CLKBUF_X1 port map( A => n295, Z => n150);
   U29 : CLKBUF_X1 port map( A => n295, Z => n149);
   U30 : CLKBUF_X1 port map( A => n295, Z => n148);
   U31 : BUF_X1 port map( A => n293, Z => n138);
   U32 : BUF_X1 port map( A => n293, Z => n137);
   U33 : BUF_X1 port map( A => n293, Z => n136);
   U34 : BUF_X1 port map( A => n293, Z => n140);
   U35 : BUF_X1 port map( A => n293, Z => n139);
   U36 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U37 : BUF_X1 port map( A => SEL(0), Z => n164);
   U38 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U39 : INV_X1 port map( A => SEL(2), ZN => n166);
   U40 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U41 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U42 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U43 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U44 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U45 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U46 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U47 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U48 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U49 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U50 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U51 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U52 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U53 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U54 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U55 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U56 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U57 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U58 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U59 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U60 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U61 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U62 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U63 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U64 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U65 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U66 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U67 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U68 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U69 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U70 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U71 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U72 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U73 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U74 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U75 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U76 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U77 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U78 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U79 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U80 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U81 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U82 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U83 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U84 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U85 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U86 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U87 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U88 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U89 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U90 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U91 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U92 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U93 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U94 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U95 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U96 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U97 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U98 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U99 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2 
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U100 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 
                           => n163, ZN => n256);
   U101 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U102 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U103 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U104 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U105 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U106 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U107 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U108 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U109 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U110 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U111 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U112 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U113 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U114 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 
                           => n162, ZN => n234);
   U115 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U116 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U117 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U118 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U119 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U120 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U121 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U122 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U123 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U124 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U125 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U126 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U127 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U128 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U129 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U130 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U131 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U132 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U133 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U134 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U135 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U136 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U137 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U138 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U139 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U140 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U141 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U142 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U143 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U144 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U145 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U146 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U147 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U148 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U149 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U150 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U151 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U152 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U153 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U154 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U155 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U156 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U157 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U158 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U159 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U160 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U161 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U162 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U163 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U164 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U165 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U166 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U167 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U168 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U169 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U170 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U171 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U172 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U173 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U174 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U175 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U176 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U177 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U178 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U179 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U180 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U181 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U182 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U183 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U184 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 
                           => n161, ZN => n212);
   U185 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U186 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U187 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 
                           => n161, ZN => n190);
   U188 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U189 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U190 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U191 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U192 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U193 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U194 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U195 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U196 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U197 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U198 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U199 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U200 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U201 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U202 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U203 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U204 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U205 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U206 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U207 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U208 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U209 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U210 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U211 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U212 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U213 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U214 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U215 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U216 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U217 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U218 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U219 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U220 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U221 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U222 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_11 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_11;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_11 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U2 : BUF_X1 port map( A => n294, Z => n146);
   U3 : BUF_X1 port map( A => n296, Z => n158);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U5 : CLKBUF_X1 port map( A => n296, Z => n156);
   U6 : CLKBUF_X1 port map( A => n295, Z => n150);
   U7 : CLKBUF_X1 port map( A => n296, Z => n155);
   U8 : CLKBUF_X1 port map( A => n295, Z => n149);
   U9 : CLKBUF_X1 port map( A => n296, Z => n154);
   U10 : CLKBUF_X1 port map( A => n295, Z => n148);
   U11 : CLKBUF_X1 port map( A => n295, Z => n152);
   U12 : CLKBUF_X1 port map( A => n294, Z => n144);
   U13 : CLKBUF_X1 port map( A => n294, Z => n143);
   U14 : CLKBUF_X1 port map( A => n294, Z => n142);
   U15 : BUF_X1 port map( A => n295, Z => n151);
   U16 : BUF_X1 port map( A => n294, Z => n145);
   U17 : BUF_X1 port map( A => n296, Z => n157);
   U18 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U19 : BUF_X1 port map( A => n293, Z => n140);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : BUF_X1 port map( A => n293, Z => n139);
   U24 : BUF_X1 port map( A => SEL(0), Z => n164);
   U25 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U26 : BUF_X1 port map( A => SEL(0), Z => n163);
   U27 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U28 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U29 : INV_X1 port map( A => SEL(2), ZN => n166);
   U30 : BUF_X1 port map( A => SEL(0), Z => n162);
   U31 : BUF_X1 port map( A => SEL(0), Z => n161);
   U32 : BUF_X1 port map( A => SEL(0), Z => n160);
   U33 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U34 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U35 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U36 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U37 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U38 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U39 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U40 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U41 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U42 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U43 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U44 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U45 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U46 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U47 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U48 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U49 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U50 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U51 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U52 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U53 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U54 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U55 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U56 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U57 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U58 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U59 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U60 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U61 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U62 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U63 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U64 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U65 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U66 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U67 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U68 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U69 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U70 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U71 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U72 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U73 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U74 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U75 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U76 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U77 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U78 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U79 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U80 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U81 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U82 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U83 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U84 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U85 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U86 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U87 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U88 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U89 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U90 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U91 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U92 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U93 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U94 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U95 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U96 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U97 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U98 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U99 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U100 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U101 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U102 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U103 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U104 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U105 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U106 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U107 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U108 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U109 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U110 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U111 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U112 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U113 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U114 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U115 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U116 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U117 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U118 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U119 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U120 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U121 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U122 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U123 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U124 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U125 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U126 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U127 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U128 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U129 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U130 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U131 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U132 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U133 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U134 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U135 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U136 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U137 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U138 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U139 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U140 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U141 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U142 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U143 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U144 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U145 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U146 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U147 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U148 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U149 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U150 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U151 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U152 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U153 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U154 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U155 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U156 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U157 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U158 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U159 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U160 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U161 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U162 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U163 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U164 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U165 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U166 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U167 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U168 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U169 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U170 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U171 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U172 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U173 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U174 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U175 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U176 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U177 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U178 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U179 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U180 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U181 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U182 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U183 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U184 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U185 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U186 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U187 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U188 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U189 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U190 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U191 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U192 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U193 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U194 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U195 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U196 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U197 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U198 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U199 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U200 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U201 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U202 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U203 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U204 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U205 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U206 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U207 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U208 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U209 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U210 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U211 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U212 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U213 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U214 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U215 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U216 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U217 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U218 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U219 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U220 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U221 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U222 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_10 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_10;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_10 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U2 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U3 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U5 : BUF_X1 port map( A => n294, Z => n144);
   U6 : BUF_X1 port map( A => n295, Z => n151);
   U7 : BUF_X1 port map( A => n294, Z => n145);
   U8 : BUF_X1 port map( A => n296, Z => n157);
   U9 : BUF_X1 port map( A => n294, Z => n143);
   U10 : BUF_X1 port map( A => n296, Z => n156);
   U11 : BUF_X1 port map( A => n295, Z => n150);
   U12 : BUF_X1 port map( A => n296, Z => n155);
   U13 : BUF_X1 port map( A => n295, Z => n149);
   U14 : BUF_X1 port map( A => n294, Z => n142);
   U15 : BUF_X1 port map( A => n295, Z => n148);
   U16 : BUF_X1 port map( A => n296, Z => n154);
   U17 : BUF_X1 port map( A => n295, Z => n152);
   U18 : BUF_X1 port map( A => n294, Z => n146);
   U19 : BUF_X1 port map( A => n296, Z => n158);
   U20 : BUF_X1 port map( A => n293, Z => n140);
   U21 : BUF_X1 port map( A => n293, Z => n138);
   U22 : BUF_X1 port map( A => n293, Z => n137);
   U23 : BUF_X1 port map( A => n293, Z => n136);
   U24 : BUF_X1 port map( A => n293, Z => n139);
   U25 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U26 : BUF_X1 port map( A => SEL(0), Z => n163);
   U27 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U28 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U29 : INV_X1 port map( A => SEL(2), ZN => n166);
   U30 : BUF_X1 port map( A => SEL(0), Z => n162);
   U31 : BUF_X1 port map( A => SEL(0), Z => n161);
   U32 : BUF_X1 port map( A => SEL(0), Z => n160);
   U33 : BUF_X1 port map( A => SEL(0), Z => n164);
   U34 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U35 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U36 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U37 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U38 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U39 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U40 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U41 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U42 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U43 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U44 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U45 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U46 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U47 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U48 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U49 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U50 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U51 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U52 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U53 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U54 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U55 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U56 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U57 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U58 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U59 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U60 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U61 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U62 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U63 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U64 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U65 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U66 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U67 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U68 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U69 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U70 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U71 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U72 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U73 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U74 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U75 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U76 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U77 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U78 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U79 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U80 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U81 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U82 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U83 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U84 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U85 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U86 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U87 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U88 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U89 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U90 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U91 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U92 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U93 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U94 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U95 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U96 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2 
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U97 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U98 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U99 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2 
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U100 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U101 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U102 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U103 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U104 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U105 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U106 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U107 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U108 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U109 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U110 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U111 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U112 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U113 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U114 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U115 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U116 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U117 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U118 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U119 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 
                           => n162, ZN => n234);
   U120 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U121 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U122 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U123 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U124 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U125 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U126 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U127 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U128 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U129 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U130 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U131 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U132 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U133 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U134 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U135 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U136 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U137 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U138 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U139 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U140 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U141 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U142 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U143 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U144 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U145 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U146 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U147 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U148 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U149 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U150 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U151 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U152 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U153 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U154 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U155 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U156 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U157 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U158 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U159 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U160 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U161 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U162 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U163 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U164 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U165 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U166 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U167 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U168 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U169 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U170 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U171 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U172 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 
                           => n161, ZN => n212);
   U173 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U174 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U175 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 
                           => n161, ZN => n190);
   U176 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U177 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U178 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U179 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U180 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U181 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U182 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U183 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U184 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U185 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U186 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U187 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U188 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U189 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U190 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U191 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U192 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U193 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U194 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U195 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U196 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U197 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U198 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U199 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U200 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U201 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U202 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U203 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U204 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U205 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U206 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U207 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U208 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U209 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U210 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U211 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U212 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U213 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U214 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U215 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U216 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U217 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U218 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U219 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U220 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U221 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U222 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_9 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_9;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_9 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U2 : BUF_X1 port map( A => n295, Z => n151);
   U3 : BUF_X1 port map( A => n294, Z => n145);
   U4 : BUF_X1 port map( A => n296, Z => n157);
   U5 : BUF_X1 port map( A => n294, Z => n144);
   U6 : BUF_X1 port map( A => n296, Z => n156);
   U7 : BUF_X1 port map( A => n295, Z => n150);
   U8 : BUF_X1 port map( A => n294, Z => n143);
   U9 : BUF_X1 port map( A => n296, Z => n155);
   U10 : BUF_X1 port map( A => n295, Z => n149);
   U11 : BUF_X1 port map( A => n295, Z => n148);
   U12 : BUF_X1 port map( A => n294, Z => n142);
   U13 : BUF_X1 port map( A => n296, Z => n154);
   U14 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U15 : BUF_X1 port map( A => n295, Z => n152);
   U16 : BUF_X1 port map( A => n294, Z => n146);
   U17 : BUF_X1 port map( A => n296, Z => n158);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : BUF_X1 port map( A => SEL(0), Z => n163);
   U25 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U26 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U27 : INV_X1 port map( A => SEL(2), ZN => n166);
   U28 : BUF_X1 port map( A => SEL(0), Z => n162);
   U29 : BUF_X1 port map( A => SEL(0), Z => n161);
   U30 : BUF_X1 port map( A => SEL(0), Z => n160);
   U31 : BUF_X1 port map( A => SEL(0), Z => n164);
   U32 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U33 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U34 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U35 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U36 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U37 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U38 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U39 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U40 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U41 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U42 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U43 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U44 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U45 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U46 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U47 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U48 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U49 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U50 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U51 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U52 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U53 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U54 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U55 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U56 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U57 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U58 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U59 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U60 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U61 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U62 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U63 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U64 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U65 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U66 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U67 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U68 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U69 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U70 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U71 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U72 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U73 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U74 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U75 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U76 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U77 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U78 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U79 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U80 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U81 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U82 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U83 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U84 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U85 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U86 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U87 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U88 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U89 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U90 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U91 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U92 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U93 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U94 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U95 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U96 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U97 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U98 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U99 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U100 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U101 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U102 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U103 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U104 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U105 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U106 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U107 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U108 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U109 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U110 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U111 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U112 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U113 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U114 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U115 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U116 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U117 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U118 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U119 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U120 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U121 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U122 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U123 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U124 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U125 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U126 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U127 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U128 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U129 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U130 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U131 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U132 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U133 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U134 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U135 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U136 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U137 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U138 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U139 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U140 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U141 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U142 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U143 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U144 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U145 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U146 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U147 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U148 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U149 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U150 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U151 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U152 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U153 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U154 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U155 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U156 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U157 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U158 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U159 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U160 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U161 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U162 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U163 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U164 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U165 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U166 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U167 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U168 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U169 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U170 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U171 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U172 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U173 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U174 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U175 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U176 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U177 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U178 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U179 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U180 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U181 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U182 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U183 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U184 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U185 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U186 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U187 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U188 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U189 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U190 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U191 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U192 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U193 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U194 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U195 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U196 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U197 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U198 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U199 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U200 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U201 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U202 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U203 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U204 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U205 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U206 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U207 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U208 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U209 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U210 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U211 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U212 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U213 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U214 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U215 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U216 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U217 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U218 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U219 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U220 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U221 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U222 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_8 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_8;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_8 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U2 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U3 : BUF_X1 port map( A => n295, Z => n151);
   U4 : BUF_X1 port map( A => n294, Z => n145);
   U5 : BUF_X1 port map( A => n296, Z => n157);
   U6 : BUF_X1 port map( A => n294, Z => n144);
   U7 : BUF_X1 port map( A => n296, Z => n156);
   U8 : BUF_X1 port map( A => n295, Z => n150);
   U9 : BUF_X1 port map( A => n294, Z => n143);
   U10 : BUF_X1 port map( A => n296, Z => n155);
   U11 : BUF_X1 port map( A => n295, Z => n149);
   U12 : BUF_X1 port map( A => n295, Z => n148);
   U13 : BUF_X1 port map( A => n294, Z => n142);
   U14 : BUF_X1 port map( A => n296, Z => n154);
   U15 : BUF_X1 port map( A => n295, Z => n152);
   U16 : BUF_X1 port map( A => n294, Z => n146);
   U17 : BUF_X1 port map( A => n296, Z => n158);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : BUF_X1 port map( A => SEL(0), Z => n163);
   U25 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U26 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U27 : INV_X1 port map( A => SEL(2), ZN => n166);
   U28 : BUF_X1 port map( A => SEL(0), Z => n162);
   U29 : BUF_X1 port map( A => SEL(0), Z => n161);
   U30 : BUF_X1 port map( A => SEL(0), Z => n160);
   U31 : BUF_X1 port map( A => SEL(0), Z => n164);
   U32 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U34 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U35 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U36 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U37 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U38 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U39 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U40 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U41 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U42 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U43 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U44 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U45 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U46 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U47 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U48 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U49 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U50 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U51 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U52 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U53 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U54 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U55 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U56 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U57 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U58 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U59 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U60 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U61 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U62 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U63 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U64 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U65 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U66 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U67 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U68 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U69 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U70 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U71 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U72 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U73 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U74 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U75 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U76 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U77 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U78 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U79 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U80 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U81 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U82 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U83 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U84 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U85 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U86 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U87 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U88 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U89 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U90 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U91 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U92 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U93 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U94 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U95 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U96 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U97 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2 
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U98 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U99 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U100 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U101 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U102 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U103 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U104 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U105 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U106 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U107 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U108 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U109 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U110 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U111 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U112 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U113 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U114 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U115 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U116 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U117 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U118 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U119 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U120 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U121 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U122 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U123 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U124 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U125 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U126 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U127 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U128 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U129 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U130 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U131 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U132 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U133 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U134 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U135 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U136 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U137 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U138 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U139 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U140 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U141 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U142 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U143 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U144 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U145 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U146 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U147 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U148 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U149 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U150 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U151 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U152 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U153 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U154 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U155 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U156 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U157 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U158 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U159 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U160 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U161 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U162 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 
                           => n161, ZN => n212);
   U163 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U164 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U165 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 
                           => n161, ZN => n190);
   U166 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U167 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U168 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U169 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U170 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U171 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U172 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U173 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U174 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U175 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U176 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U177 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U178 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U179 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U180 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U181 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U182 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U183 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U184 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U185 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U186 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U187 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U188 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U189 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U190 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U191 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U192 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U193 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U194 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U195 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U196 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U197 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U198 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U199 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U200 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U201 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U202 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U203 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U204 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U205 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U206 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U207 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U208 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U209 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U210 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U211 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U212 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U213 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U214 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U215 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U216 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U217 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U218 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U219 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U220 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U221 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U222 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_7 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_7;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_7 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U2 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U3 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U4 : BUF_X1 port map( A => n294, Z => n145);
   U5 : BUF_X1 port map( A => n295, Z => n151);
   U6 : BUF_X1 port map( A => n294, Z => n144);
   U7 : BUF_X1 port map( A => n296, Z => n157);
   U8 : BUF_X1 port map( A => n296, Z => n156);
   U9 : BUF_X1 port map( A => n295, Z => n150);
   U10 : BUF_X1 port map( A => n294, Z => n143);
   U11 : BUF_X1 port map( A => n296, Z => n155);
   U12 : BUF_X1 port map( A => n295, Z => n149);
   U13 : BUF_X1 port map( A => n295, Z => n148);
   U14 : BUF_X1 port map( A => n294, Z => n142);
   U15 : BUF_X1 port map( A => n296, Z => n154);
   U16 : BUF_X1 port map( A => n295, Z => n152);
   U17 : BUF_X1 port map( A => n294, Z => n146);
   U18 : BUF_X1 port map( A => n296, Z => n158);
   U19 : BUF_X1 port map( A => n293, Z => n140);
   U20 : BUF_X1 port map( A => n293, Z => n139);
   U21 : BUF_X1 port map( A => n293, Z => n138);
   U22 : BUF_X1 port map( A => n293, Z => n137);
   U23 : BUF_X1 port map( A => n293, Z => n136);
   U24 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U25 : INV_X1 port map( A => SEL(2), ZN => n166);
   U26 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U27 : BUF_X1 port map( A => SEL(0), Z => n163);
   U28 : BUF_X1 port map( A => SEL(0), Z => n162);
   U29 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U30 : BUF_X1 port map( A => SEL(0), Z => n161);
   U31 : BUF_X1 port map( A => SEL(0), Z => n160);
   U32 : BUF_X1 port map( A => SEL(0), Z => n164);
   U33 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U34 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U35 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U36 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U37 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U38 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U39 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U40 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U41 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U42 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U43 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U44 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U45 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U46 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U47 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U48 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U49 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U50 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U51 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U52 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U53 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U54 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U55 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U56 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U57 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U58 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U59 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U60 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U61 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U62 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U63 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U64 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U65 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U66 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U67 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U68 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U69 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U70 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U71 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U72 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U73 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U74 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U75 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U76 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U77 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U78 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U79 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U80 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U81 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U82 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U83 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U84 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U85 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U86 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U87 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U88 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U89 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U90 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U91 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U92 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U93 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U94 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U95 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U96 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U97 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U98 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U99 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U100 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U101 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U102 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U103 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U104 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U105 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U106 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U107 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U108 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U109 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U110 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U111 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U112 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U113 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U114 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U115 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U116 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U117 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U118 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U119 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U120 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U121 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U122 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U123 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U124 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U125 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U126 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U127 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U128 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U129 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U130 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U131 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U132 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U133 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U134 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U135 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U136 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U137 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U138 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U139 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U140 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U141 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U142 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U143 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U144 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U145 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U146 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U147 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U148 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U149 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U150 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U151 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U152 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U153 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U154 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U155 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U156 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U157 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U158 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U159 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U160 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U161 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U162 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U163 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U164 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U165 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U166 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U167 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U168 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U169 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U170 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U171 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U172 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U173 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U174 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U175 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U176 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U177 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U178 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U179 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U180 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U181 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U182 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U183 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U184 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U185 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U186 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U187 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U188 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U189 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U190 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U191 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U192 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U193 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U194 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U195 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U196 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U197 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U198 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U199 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U200 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U201 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U202 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U203 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U204 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U205 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U206 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U207 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U208 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U209 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U210 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U211 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U212 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U213 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U214 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U215 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U216 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U217 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U218 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U219 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U220 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U221 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U222 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_6 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_6;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_6 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U2 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U3 : BUF_X1 port map( A => n295, Z => n151);
   U4 : BUF_X1 port map( A => n294, Z => n145);
   U5 : BUF_X1 port map( A => n294, Z => n144);
   U6 : BUF_X1 port map( A => n296, Z => n157);
   U7 : BUF_X1 port map( A => n296, Z => n156);
   U8 : BUF_X1 port map( A => n295, Z => n150);
   U9 : BUF_X1 port map( A => n294, Z => n143);
   U10 : BUF_X1 port map( A => n296, Z => n155);
   U11 : BUF_X1 port map( A => n295, Z => n149);
   U12 : BUF_X1 port map( A => n295, Z => n148);
   U13 : BUF_X1 port map( A => n294, Z => n142);
   U14 : BUF_X1 port map( A => n296, Z => n154);
   U15 : BUF_X1 port map( A => n295, Z => n152);
   U16 : BUF_X1 port map( A => n294, Z => n146);
   U17 : BUF_X1 port map( A => n296, Z => n158);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : BUF_X1 port map( A => SEL(0), Z => n163);
   U25 : BUF_X1 port map( A => SEL(0), Z => n162);
   U26 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U27 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U28 : INV_X1 port map( A => SEL(2), ZN => n166);
   U29 : BUF_X1 port map( A => SEL(0), Z => n161);
   U30 : BUF_X1 port map( A => SEL(0), Z => n160);
   U31 : BUF_X1 port map( A => SEL(0), Z => n164);
   U32 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U33 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U34 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U35 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U36 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U37 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U38 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U39 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U40 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U41 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U42 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U43 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U44 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U45 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U46 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U47 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U48 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U49 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U50 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U51 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U52 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U53 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U54 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U55 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U56 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U57 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U58 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U59 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U60 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U61 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U62 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U63 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U64 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U65 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U66 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U67 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U68 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U69 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U70 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U71 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U72 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U73 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U74 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U75 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U76 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U77 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U78 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U79 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U80 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U81 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U82 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U83 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U84 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U85 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U86 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U87 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U88 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U89 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U90 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U91 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U92 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U93 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U94 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U95 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U96 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U97 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U98 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U99 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U100 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U101 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U102 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U103 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U104 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U105 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U106 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U107 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U108 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U109 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U110 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U111 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U112 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U113 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U114 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U115 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U116 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U117 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U118 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U119 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U120 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U121 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U122 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U123 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U124 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U125 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U126 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U127 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U128 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U129 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U130 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U131 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U132 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U133 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U134 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U135 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U136 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U137 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U138 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U139 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U140 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U141 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U142 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U143 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U144 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U145 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U146 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U147 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U148 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U149 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U150 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U151 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U152 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U153 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 
                           => n161, ZN => n190);
   U154 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U155 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U156 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U157 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U158 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U159 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U160 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U161 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U162 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U163 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U164 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U165 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U166 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U167 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U168 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U169 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U170 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U171 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U172 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U173 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U174 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U175 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U176 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U177 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U178 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U179 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U180 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U181 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U182 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U183 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U184 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U185 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U186 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U187 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U188 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U189 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U190 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U191 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U192 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U193 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U194 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U195 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U196 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U197 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U198 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U199 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U200 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U201 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U202 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U203 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U204 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U205 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U206 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U207 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U208 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U209 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U210 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U211 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U212 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U213 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U214 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U215 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U216 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U217 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U218 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U219 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U220 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U221 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U222 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_5 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_5;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U2 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U3 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U4 : BUF_X1 port map( A => n294, Z => n144);
   U5 : BUF_X1 port map( A => n296, Z => n156);
   U6 : BUF_X1 port map( A => n295, Z => n150);
   U7 : BUF_X1 port map( A => n294, Z => n143);
   U8 : BUF_X1 port map( A => n296, Z => n155);
   U9 : BUF_X1 port map( A => n295, Z => n149);
   U10 : BUF_X1 port map( A => n295, Z => n148);
   U11 : BUF_X1 port map( A => n294, Z => n142);
   U12 : BUF_X1 port map( A => n296, Z => n154);
   U13 : BUF_X1 port map( A => n295, Z => n152);
   U14 : BUF_X1 port map( A => n294, Z => n146);
   U15 : BUF_X1 port map( A => n296, Z => n158);
   U16 : BUF_X1 port map( A => n295, Z => n151);
   U17 : BUF_X1 port map( A => n294, Z => n145);
   U18 : BUF_X1 port map( A => n296, Z => n157);
   U19 : BUF_X1 port map( A => n293, Z => n140);
   U20 : BUF_X1 port map( A => n293, Z => n139);
   U21 : BUF_X1 port map( A => n293, Z => n138);
   U22 : BUF_X1 port map( A => n293, Z => n137);
   U23 : BUF_X1 port map( A => n293, Z => n136);
   U24 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U25 : BUF_X1 port map( A => SEL(0), Z => n162);
   U26 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U27 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U28 : INV_X1 port map( A => SEL(2), ZN => n166);
   U29 : BUF_X1 port map( A => SEL(0), Z => n161);
   U30 : BUF_X1 port map( A => SEL(0), Z => n160);
   U31 : BUF_X1 port map( A => SEL(0), Z => n164);
   U32 : BUF_X1 port map( A => SEL(0), Z => n163);
   U33 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U34 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U35 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U36 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U37 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U38 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U39 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U40 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U41 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U42 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U43 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U44 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U45 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U46 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U47 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U48 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U49 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U50 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U51 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U52 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U53 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U54 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U55 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U56 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U57 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U58 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U59 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U60 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U61 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U62 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U63 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U64 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U65 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U66 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U67 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U68 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U69 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U70 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U71 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U72 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U73 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U74 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U75 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U76 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U77 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U78 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U79 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U80 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U81 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U82 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U83 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U84 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U85 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U86 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U87 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U88 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U89 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U90 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U91 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U92 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U93 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U94 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U95 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U96 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U97 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U98 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U99 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U100 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U101 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U102 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U103 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U104 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U105 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U106 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U107 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U108 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U109 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U110 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U111 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U112 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U113 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U114 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U115 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U116 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U117 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U118 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U119 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U120 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U121 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U122 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U123 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U124 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U125 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U126 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U127 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U128 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U129 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U130 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U131 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U132 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U133 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U134 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U135 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U136 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U137 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U138 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U139 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U140 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U141 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U142 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U143 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U144 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U145 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U146 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U147 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U148 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U149 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U150 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U151 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U152 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U153 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U154 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U155 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U156 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U157 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U158 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U159 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U160 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U161 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U162 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U163 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U164 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U165 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U166 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U167 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U168 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U169 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U170 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U171 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U172 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U173 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U174 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U175 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U176 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U177 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U178 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U179 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U180 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U181 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U182 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U183 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U184 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U185 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U186 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U187 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U188 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U189 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U190 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U191 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U192 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U193 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U194 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U195 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U196 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U197 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U198 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U199 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U200 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U201 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U202 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U203 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U204 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U205 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U206 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U207 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U208 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U209 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U210 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U211 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U212 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U213 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U214 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U215 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U216 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U217 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U218 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U219 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U220 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U221 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U222 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_4 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_4;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U2 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U3 : BUF_X1 port map( A => n294, Z => n144);
   U4 : BUF_X1 port map( A => n296, Z => n156);
   U5 : BUF_X1 port map( A => n294, Z => n143);
   U6 : BUF_X1 port map( A => n296, Z => n155);
   U7 : BUF_X1 port map( A => n295, Z => n150);
   U8 : BUF_X1 port map( A => n295, Z => n149);
   U9 : BUF_X1 port map( A => n295, Z => n148);
   U10 : BUF_X1 port map( A => n294, Z => n142);
   U11 : BUF_X1 port map( A => n296, Z => n154);
   U12 : BUF_X1 port map( A => n295, Z => n152);
   U13 : BUF_X1 port map( A => n295, Z => n151);
   U14 : BUF_X1 port map( A => n294, Z => n146);
   U15 : BUF_X1 port map( A => n294, Z => n145);
   U16 : BUF_X1 port map( A => n296, Z => n158);
   U17 : BUF_X1 port map( A => n296, Z => n157);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U25 : INV_X1 port map( A => SEL(2), ZN => n166);
   U26 : BUF_X1 port map( A => SEL(0), Z => n162);
   U27 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U28 : BUF_X1 port map( A => SEL(0), Z => n160);
   U29 : BUF_X1 port map( A => SEL(0), Z => n161);
   U30 : BUF_X1 port map( A => SEL(0), Z => n164);
   U31 : BUF_X1 port map( A => SEL(0), Z => n163);
   U32 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U33 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U34 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U35 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U36 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U37 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U38 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U39 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U40 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U41 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U42 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U43 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U44 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U45 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U46 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U47 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U48 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U49 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U50 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U51 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U52 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U53 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U54 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U55 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U56 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U57 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U58 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U59 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U60 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U61 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U62 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U63 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U64 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U65 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U66 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U67 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U68 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U69 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U70 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U71 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U72 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U73 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U74 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U75 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U76 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U77 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U78 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U79 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U80 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U81 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U82 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U83 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U84 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U85 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U86 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U87 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U88 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U89 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U90 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U91 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U92 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U93 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U94 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U95 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U96 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U97 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U98 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U99 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U100 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U101 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U102 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U103 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U104 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U105 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U106 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U107 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U108 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U109 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U110 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U111 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U112 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U113 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U114 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U115 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U116 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U117 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U118 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U119 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U120 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U121 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U122 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U123 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U124 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U125 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U126 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U127 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U128 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U129 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U130 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U131 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U132 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U133 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U134 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U135 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U136 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U137 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U138 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U139 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U140 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U141 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U142 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U143 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U144 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U145 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U146 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U147 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U148 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U149 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U150 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U151 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U152 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U153 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U154 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U155 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U156 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U157 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U158 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U159 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U160 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U161 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U162 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U163 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U164 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U165 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U166 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U167 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U168 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U169 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U170 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U171 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U172 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U173 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U174 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U175 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U176 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U177 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U178 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U179 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U180 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U181 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U182 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U183 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U184 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U185 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U186 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U187 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U188 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U189 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U190 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U191 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U192 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U193 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U194 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U195 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U196 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U197 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U198 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U199 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U200 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U201 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U202 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U203 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U204 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U205 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U206 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U207 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U208 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U209 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U210 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U211 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U212 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U213 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U214 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U215 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U216 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U217 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U218 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U219 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U220 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U221 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U222 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_3 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_3;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U2 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U3 : BUF_X1 port map( A => n294, Z => n144);
   U4 : BUF_X1 port map( A => n294, Z => n143);
   U5 : BUF_X1 port map( A => n296, Z => n156);
   U6 : BUF_X1 port map( A => n296, Z => n155);
   U7 : BUF_X1 port map( A => n295, Z => n150);
   U8 : BUF_X1 port map( A => n295, Z => n149);
   U9 : BUF_X1 port map( A => n295, Z => n148);
   U10 : BUF_X1 port map( A => n294, Z => n142);
   U11 : BUF_X1 port map( A => n296, Z => n154);
   U12 : BUF_X1 port map( A => n295, Z => n152);
   U13 : BUF_X1 port map( A => n295, Z => n151);
   U14 : BUF_X1 port map( A => n294, Z => n146);
   U15 : BUF_X1 port map( A => n294, Z => n145);
   U16 : BUF_X1 port map( A => n296, Z => n158);
   U17 : BUF_X1 port map( A => n296, Z => n157);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : BUF_X1 port map( A => SEL(0), Z => n162);
   U25 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U26 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U27 : INV_X1 port map( A => SEL(2), ZN => n166);
   U28 : BUF_X1 port map( A => SEL(0), Z => n161);
   U29 : BUF_X1 port map( A => SEL(0), Z => n160);
   U30 : BUF_X1 port map( A => SEL(0), Z => n164);
   U31 : BUF_X1 port map( A => SEL(0), Z => n163);
   U32 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U33 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U34 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U35 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U36 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 =>
                           n160, ZN => n168);
   U37 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U38 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U39 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U40 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U41 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U42 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U43 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U44 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U45 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U46 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U47 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U48 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U49 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U50 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U51 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U52 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U53 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U54 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U55 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U56 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U57 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U58 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U59 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U60 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U61 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U62 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U63 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U64 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U65 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U66 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U67 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U68 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U69 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U70 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U71 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U72 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U73 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U74 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U75 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U76 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U77 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U78 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U79 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U80 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U81 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U82 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U83 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U84 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U85 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U86 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U87 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U88 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U89 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U90 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U91 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U92 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U93 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U94 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U95 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U96 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U97 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U98 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U99 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U100 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U101 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U102 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U103 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U104 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U105 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U106 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U107 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U108 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U109 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U110 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U111 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U112 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U113 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U114 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U115 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U116 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U117 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U118 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U119 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U120 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U121 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U122 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U123 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U124 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U125 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U126 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U127 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U128 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U129 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U130 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U131 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U132 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U133 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U134 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U135 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U136 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U137 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U138 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U139 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U140 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U141 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U142 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U143 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U144 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U145 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U146 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U147 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U148 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U149 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U150 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U151 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U152 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U153 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U154 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U155 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U156 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U157 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U158 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U159 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U160 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U161 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U162 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U163 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U164 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U165 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U166 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U167 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U168 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U169 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U170 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U171 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U172 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U173 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U174 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U175 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U176 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U177 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U178 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U179 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U180 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U181 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U182 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U183 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U184 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U185 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U186 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U187 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U188 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U189 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U190 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U191 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U192 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U193 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U194 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U195 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U196 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U197 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U198 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U199 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U200 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U201 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U202 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U203 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U204 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U205 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U206 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U207 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U208 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U209 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U210 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U211 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U212 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U213 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U214 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U215 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U216 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U217 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U218 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U219 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U220 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U221 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U222 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_2 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_2;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_2 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U2 : BUF_X1 port map( A => n294, Z => n144);
   U3 : BUF_X1 port map( A => n296, Z => n156);
   U4 : BUF_X1 port map( A => n295, Z => n150);
   U5 : BUF_X1 port map( A => n294, Z => n143);
   U6 : BUF_X1 port map( A => n296, Z => n155);
   U7 : BUF_X1 port map( A => n295, Z => n149);
   U8 : BUF_X1 port map( A => n295, Z => n148);
   U9 : BUF_X1 port map( A => n294, Z => n142);
   U10 : BUF_X1 port map( A => n296, Z => n154);
   U11 : BUF_X1 port map( A => n295, Z => n152);
   U12 : BUF_X1 port map( A => n295, Z => n151);
   U13 : BUF_X1 port map( A => n294, Z => n146);
   U14 : BUF_X1 port map( A => n294, Z => n145);
   U15 : BUF_X1 port map( A => n296, Z => n158);
   U16 : BUF_X1 port map( A => n296, Z => n157);
   U17 : BUF_X1 port map( A => n293, Z => n140);
   U18 : BUF_X1 port map( A => n293, Z => n139);
   U19 : BUF_X1 port map( A => n293, Z => n138);
   U20 : BUF_X1 port map( A => n293, Z => n137);
   U21 : BUF_X1 port map( A => n293, Z => n136);
   U22 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U23 : BUF_X1 port map( A => SEL(0), Z => n162);
   U24 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U25 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U26 : INV_X1 port map( A => SEL(2), ZN => n166);
   U27 : BUF_X1 port map( A => SEL(0), Z => n161);
   U28 : BUF_X1 port map( A => SEL(0), Z => n160);
   U29 : BUF_X1 port map( A => SEL(0), Z => n164);
   U30 : BUF_X1 port map( A => SEL(0), Z => n163);
   U31 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U32 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U33 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U34 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U35 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U36 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U37 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U38 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U39 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U40 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U41 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U42 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U43 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U44 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U45 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U46 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U47 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U48 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U49 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U50 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U51 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U52 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U53 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U54 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U55 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U56 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U57 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U58 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U59 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U60 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U61 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U62 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U63 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U64 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U65 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U66 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U67 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U68 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U69 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U70 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U71 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U72 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U73 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U74 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U75 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U76 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U77 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U78 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U79 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U80 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U81 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U82 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U83 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U84 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U85 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U86 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U87 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2 
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U88 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U89 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U90 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2 
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U91 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U92 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U93 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2 
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U94 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U95 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U96 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2 
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U97 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U98 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U99 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2 
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U100 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U101 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U102 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U103 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U104 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U105 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U106 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U107 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U108 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U109 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U110 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U111 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U112 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U113 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U114 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U115 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U116 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U117 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U118 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U119 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U120 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U121 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U122 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U123 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U124 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U125 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U126 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U127 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U128 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U129 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U130 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U131 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U132 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U133 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U134 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U135 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U136 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U137 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U138 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U139 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U140 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U141 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U142 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U143 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U144 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U145 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U146 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U147 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U148 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U149 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U150 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U151 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U152 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U153 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U154 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U155 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U156 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U157 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U158 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U159 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U160 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U161 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U162 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U163 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U164 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U165 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U166 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U167 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U168 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U169 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U170 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U171 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U172 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U173 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U174 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U175 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U176 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U177 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U178 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U179 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U180 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U181 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U182 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U183 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U184 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U185 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U186 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U187 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U188 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U189 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U190 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U191 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U192 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U193 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U194 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U195 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U196 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U197 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U198 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U199 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U200 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U201 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U202 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U203 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U204 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U205 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U206 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U207 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U208 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U209 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U210 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U211 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U212 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U213 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U214 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U215 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U216 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U217 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U218 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U219 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U220 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U221 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U222 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_1 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_1;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n160, ZN => n293);
   U2 : AOI222_X1 port map( A1 => INPUT(64), A2 => n154, B1 => INPUT(192), B2 
                           => n148, C1 => INPUT(128), C2 => n142, ZN => n167);
   U3 : BUF_X1 port map( A => n294, Z => n144);
   U4 : BUF_X1 port map( A => n296, Z => n156);
   U5 : BUF_X1 port map( A => n294, Z => n143);
   U6 : BUF_X1 port map( A => n296, Z => n155);
   U7 : BUF_X1 port map( A => n295, Z => n150);
   U8 : BUF_X1 port map( A => n295, Z => n149);
   U9 : BUF_X1 port map( A => n295, Z => n148);
   U10 : BUF_X1 port map( A => n294, Z => n142);
   U11 : BUF_X1 port map( A => n296, Z => n154);
   U12 : BUF_X1 port map( A => n295, Z => n152);
   U13 : BUF_X1 port map( A => n295, Z => n151);
   U14 : BUF_X1 port map( A => n294, Z => n146);
   U15 : BUF_X1 port map( A => n294, Z => n145);
   U16 : BUF_X1 port map( A => n296, Z => n158);
   U17 : BUF_X1 port map( A => n296, Z => n157);
   U18 : BUF_X1 port map( A => n293, Z => n140);
   U19 : BUF_X1 port map( A => n293, Z => n139);
   U20 : BUF_X1 port map( A => n293, Z => n138);
   U21 : BUF_X1 port map( A => n293, Z => n137);
   U22 : BUF_X1 port map( A => n293, Z => n136);
   U23 : NOR2_X1 port map( A1 => n166, A2 => SEL(1), ZN => n296);
   U24 : AND2_X1 port map( A1 => SEL(1), A2 => n166, ZN => n294);
   U25 : INV_X1 port map( A => SEL(2), ZN => n166);
   U26 : BUF_X1 port map( A => SEL(0), Z => n162);
   U27 : BUF_X1 port map( A => SEL(0), Z => n161);
   U28 : AND2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => n295);
   U29 : BUF_X1 port map( A => SEL(0), Z => n160);
   U30 : BUF_X1 port map( A => SEL(0), Z => n164);
   U31 : BUF_X1 port map( A => SEL(0), Z => n163);
   U32 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(1));
   U33 : AOI222_X1 port map( A1 => INPUT(65), A2 => n154, B1 => INPUT(193), B2 
                           => n148, C1 => INPUT(129), C2 => n142, ZN => n189);
   U34 : AOI22_X1 port map( A1 => INPUT(1), A2 => n136, B1 => INPUT(257), B2 =>
                           n161, ZN => n190);
   U35 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(2));
   U36 : AOI22_X1 port map( A1 => INPUT(2), A2 => n137, B1 => INPUT(258), B2 =>
                           n161, ZN => n212);
   U37 : AOI222_X1 port map( A1 => INPUT(66), A2 => n155, B1 => INPUT(194), B2 
                           => n149, C1 => INPUT(130), C2 => n143, ZN => n211);
   U38 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(3));
   U39 : AOI22_X1 port map( A1 => INPUT(3), A2 => n138, B1 => INPUT(259), B2 =>
                           n162, ZN => n234);
   U40 : AOI222_X1 port map( A1 => INPUT(67), A2 => n156, B1 => INPUT(195), B2 
                           => n150, C1 => INPUT(131), C2 => n144, ZN => n233);
   U41 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(4));
   U42 : AOI22_X1 port map( A1 => INPUT(4), A2 => n139, B1 => INPUT(260), B2 =>
                           n163, ZN => n256);
   U43 : AOI222_X1 port map( A1 => INPUT(68), A2 => n157, B1 => INPUT(196), B2 
                           => n151, C1 => INPUT(132), C2 => n145, ZN => n255);
   U44 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(5));
   U45 : AOI22_X1 port map( A1 => INPUT(5), A2 => n140, B1 => INPUT(261), B2 =>
                           n164, ZN => n278);
   U46 : AOI222_X1 port map( A1 => INPUT(69), A2 => n158, B1 => INPUT(197), B2 
                           => n152, C1 => INPUT(133), C2 => n146, ZN => n277);
   U47 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(6));
   U48 : AOI22_X1 port map( A1 => INPUT(6), A2 => n141, B1 => INPUT(262), B2 =>
                           n165, ZN => n288);
   U49 : AOI222_X1 port map( A1 => INPUT(70), A2 => n159, B1 => INPUT(198), B2 
                           => n153, C1 => INPUT(134), C2 => n147, ZN => n287);
   U50 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(7));
   U51 : AOI22_X1 port map( A1 => INPUT(7), A2 => n141, B1 => INPUT(263), B2 =>
                           n165, ZN => n290);
   U52 : AOI222_X1 port map( A1 => INPUT(71), A2 => n159, B1 => INPUT(199), B2 
                           => n153, C1 => INPUT(135), C2 => n147, ZN => n289);
   U53 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(8));
   U54 : AOI22_X1 port map( A1 => INPUT(8), A2 => n141, B1 => INPUT(264), B2 =>
                           n165, ZN => n292);
   U55 : AOI222_X1 port map( A1 => INPUT(72), A2 => n159, B1 => INPUT(200), B2 
                           => n153, C1 => INPUT(136), C2 => n147, ZN => n291);
   U56 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(9));
   U57 : AOI22_X1 port map( A1 => INPUT(9), A2 => n141, B1 => n165, B2 => 
                           INPUT(265), ZN => n298);
   U58 : AOI222_X1 port map( A1 => INPUT(73), A2 => n159, B1 => INPUT(201), B2 
                           => n153, C1 => INPUT(137), C2 => n147, ZN => n297);
   U59 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => Y(10));
   U60 : AOI22_X1 port map( A1 => INPUT(10), A2 => n136, B1 => INPUT(266), B2 
                           => n160, ZN => n170);
   U61 : AOI222_X1 port map( A1 => INPUT(74), A2 => n154, B1 => INPUT(202), B2 
                           => n148, C1 => INPUT(138), C2 => n142, ZN => n169);
   U62 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(11));
   U63 : AOI22_X1 port map( A1 => INPUT(11), A2 => n136, B1 => INPUT(267), B2 
                           => n160, ZN => n172);
   U64 : AOI222_X1 port map( A1 => INPUT(75), A2 => n154, B1 => INPUT(203), B2 
                           => n148, C1 => INPUT(139), C2 => n142, ZN => n171);
   U65 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(12));
   U66 : AOI22_X1 port map( A1 => INPUT(12), A2 => n136, B1 => INPUT(268), B2 
                           => n160, ZN => n174);
   U67 : AOI222_X1 port map( A1 => INPUT(76), A2 => n154, B1 => INPUT(204), B2 
                           => n148, C1 => INPUT(140), C2 => n142, ZN => n173);
   U68 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(18));
   U69 : AOI22_X1 port map( A1 => INPUT(18), A2 => n136, B1 => INPUT(274), B2 
                           => n160, ZN => n186);
   U70 : AOI222_X1 port map( A1 => INPUT(82), A2 => n154, B1 => INPUT(210), B2 
                           => n148, C1 => INPUT(146), C2 => n142, ZN => n185);
   U71 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(17));
   U72 : AOI22_X1 port map( A1 => INPUT(17), A2 => n136, B1 => INPUT(273), B2 
                           => n160, ZN => n184);
   U73 : AOI222_X1 port map( A1 => INPUT(81), A2 => n154, B1 => INPUT(209), B2 
                           => n148, C1 => INPUT(145), C2 => n142, ZN => n183);
   U74 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(16));
   U75 : AOI22_X1 port map( A1 => INPUT(16), A2 => n136, B1 => INPUT(272), B2 
                           => n160, ZN => n182);
   U76 : AOI222_X1 port map( A1 => INPUT(80), A2 => n154, B1 => INPUT(208), B2 
                           => n148, C1 => INPUT(144), C2 => n142, ZN => n181);
   U77 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(13));
   U78 : AOI22_X1 port map( A1 => INPUT(13), A2 => n136, B1 => INPUT(269), B2 
                           => n160, ZN => n176);
   U79 : AOI222_X1 port map( A1 => INPUT(77), A2 => n154, B1 => INPUT(205), B2 
                           => n148, C1 => INPUT(141), C2 => n142, ZN => n175);
   U80 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(14));
   U81 : AOI22_X1 port map( A1 => INPUT(14), A2 => n136, B1 => INPUT(270), B2 
                           => n160, ZN => n178);
   U82 : AOI222_X1 port map( A1 => INPUT(78), A2 => n154, B1 => INPUT(206), B2 
                           => n148, C1 => INPUT(142), C2 => n142, ZN => n177);
   U83 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(15));
   U84 : AOI22_X1 port map( A1 => INPUT(15), A2 => n136, B1 => INPUT(271), B2 
                           => n160, ZN => n180);
   U85 : AOI222_X1 port map( A1 => INPUT(79), A2 => n154, B1 => INPUT(207), B2 
                           => n148, C1 => INPUT(143), C2 => n142, ZN => n179);
   U86 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(32));
   U87 : AOI222_X1 port map( A1 => INPUT(96), A2 => n156, B1 => INPUT(224), B2 
                           => n150, C1 => INPUT(160), C2 => n144, ZN => n217);
   U88 : AOI22_X1 port map( A1 => INPUT(32), A2 => n138, B1 => INPUT(288), B2 
                           => n162, ZN => n218);
   U89 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(31));
   U90 : AOI22_X1 port map( A1 => INPUT(31), A2 => n138, B1 => INPUT(287), B2 
                           => n162, ZN => n216);
   U91 : AOI222_X1 port map( A1 => INPUT(95), A2 => n156, B1 => INPUT(223), B2 
                           => n150, C1 => INPUT(159), C2 => n144, ZN => n215);
   U92 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(30));
   U93 : AOI22_X1 port map( A1 => INPUT(30), A2 => n137, B1 => INPUT(286), B2 
                           => n162, ZN => n214);
   U94 : AOI222_X1 port map( A1 => INPUT(94), A2 => n155, B1 => INPUT(222), B2 
                           => n149, C1 => INPUT(158), C2 => n143, ZN => n213);
   U95 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(29));
   U96 : AOI22_X1 port map( A1 => INPUT(29), A2 => n137, B1 => INPUT(285), B2 
                           => n161, ZN => n210);
   U97 : AOI222_X1 port map( A1 => INPUT(93), A2 => n155, B1 => INPUT(221), B2 
                           => n149, C1 => INPUT(157), C2 => n143, ZN => n209);
   U98 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(28));
   U99 : AOI22_X1 port map( A1 => INPUT(28), A2 => n137, B1 => INPUT(284), B2 
                           => n161, ZN => n208);
   U100 : AOI222_X1 port map( A1 => INPUT(92), A2 => n155, B1 => INPUT(220), B2
                           => n149, C1 => INPUT(156), C2 => n143, ZN => n207);
   U101 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(27));
   U102 : AOI22_X1 port map( A1 => INPUT(27), A2 => n137, B1 => INPUT(283), B2 
                           => n161, ZN => n206);
   U103 : AOI222_X1 port map( A1 => INPUT(91), A2 => n155, B1 => INPUT(219), B2
                           => n149, C1 => INPUT(155), C2 => n143, ZN => n205);
   U104 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(26));
   U105 : AOI22_X1 port map( A1 => INPUT(26), A2 => n137, B1 => INPUT(282), B2 
                           => n161, ZN => n204);
   U106 : AOI222_X1 port map( A1 => INPUT(90), A2 => n155, B1 => INPUT(218), B2
                           => n149, C1 => INPUT(154), C2 => n143, ZN => n203);
   U107 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(25));
   U108 : AOI22_X1 port map( A1 => INPUT(25), A2 => n137, B1 => INPUT(281), B2 
                           => n161, ZN => n202);
   U109 : AOI222_X1 port map( A1 => INPUT(89), A2 => n155, B1 => INPUT(217), B2
                           => n149, C1 => INPUT(153), C2 => n143, ZN => n201);
   U110 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(24));
   U111 : AOI22_X1 port map( A1 => INPUT(24), A2 => n137, B1 => INPUT(280), B2 
                           => n161, ZN => n200);
   U112 : AOI222_X1 port map( A1 => INPUT(88), A2 => n155, B1 => INPUT(216), B2
                           => n149, C1 => INPUT(152), C2 => n143, ZN => n199);
   U113 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(23));
   U114 : AOI22_X1 port map( A1 => INPUT(23), A2 => n137, B1 => INPUT(279), B2 
                           => n161, ZN => n198);
   U115 : AOI222_X1 port map( A1 => INPUT(87), A2 => n155, B1 => INPUT(215), B2
                           => n149, C1 => INPUT(151), C2 => n143, ZN => n197);
   U116 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(22));
   U117 : AOI22_X1 port map( A1 => INPUT(22), A2 => n137, B1 => INPUT(278), B2 
                           => n161, ZN => n196);
   U118 : AOI222_X1 port map( A1 => INPUT(86), A2 => n155, B1 => INPUT(214), B2
                           => n149, C1 => INPUT(150), C2 => n143, ZN => n195);
   U119 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(21));
   U120 : AOI22_X1 port map( A1 => INPUT(21), A2 => n137, B1 => INPUT(277), B2 
                           => n161, ZN => n194);
   U121 : AOI222_X1 port map( A1 => INPUT(85), A2 => n155, B1 => INPUT(213), B2
                           => n149, C1 => INPUT(149), C2 => n143, ZN => n193);
   U122 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(20));
   U123 : AOI22_X1 port map( A1 => INPUT(20), A2 => n137, B1 => INPUT(276), B2 
                           => n161, ZN => n192);
   U124 : AOI222_X1 port map( A1 => INPUT(84), A2 => n155, B1 => INPUT(212), B2
                           => n149, C1 => INPUT(148), C2 => n143, ZN => n191);
   U125 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(19));
   U126 : AOI22_X1 port map( A1 => INPUT(19), A2 => n136, B1 => INPUT(275), B2 
                           => n160, ZN => n188);
   U127 : AOI222_X1 port map( A1 => INPUT(83), A2 => n154, B1 => INPUT(211), B2
                           => n148, C1 => INPUT(147), C2 => n142, ZN => n187);
   U128 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(33));
   U129 : AOI22_X1 port map( A1 => INPUT(33), A2 => n138, B1 => INPUT(289), B2 
                           => n162, ZN => n220);
   U130 : AOI222_X1 port map( A1 => INPUT(97), A2 => n156, B1 => INPUT(225), B2
                           => n150, C1 => INPUT(161), C2 => n144, ZN => n219);
   U131 : NAND2_X1 port map( A1 => n168, A2 => n167, ZN => Y(0));
   U132 : AOI22_X1 port map( A1 => INPUT(0), A2 => n136, B1 => INPUT(256), B2 
                           => n160, ZN => n168);
   U133 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(37));
   U134 : AOI22_X1 port map( A1 => INPUT(37), A2 => n138, B1 => INPUT(293), B2 
                           => n162, ZN => n228);
   U135 : AOI222_X1 port map( A1 => INPUT(101), A2 => n156, B1 => INPUT(229), 
                           B2 => n150, C1 => INPUT(165), C2 => n144, ZN => n227
                           );
   U136 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(36));
   U137 : AOI22_X1 port map( A1 => INPUT(36), A2 => n138, B1 => INPUT(292), B2 
                           => n162, ZN => n226);
   U138 : AOI222_X1 port map( A1 => INPUT(100), A2 => n156, B1 => INPUT(228), 
                           B2 => n150, C1 => INPUT(164), C2 => n144, ZN => n225
                           );
   U139 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(35));
   U140 : AOI22_X1 port map( A1 => INPUT(35), A2 => n138, B1 => INPUT(291), B2 
                           => n162, ZN => n224);
   U141 : AOI222_X1 port map( A1 => INPUT(99), A2 => n156, B1 => INPUT(227), B2
                           => n150, C1 => INPUT(163), C2 => n144, ZN => n223);
   U142 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(34));
   U143 : AOI22_X1 port map( A1 => INPUT(34), A2 => n138, B1 => INPUT(290), B2 
                           => n162, ZN => n222);
   U144 : AOI222_X1 port map( A1 => INPUT(98), A2 => n156, B1 => INPUT(226), B2
                           => n150, C1 => INPUT(162), C2 => n144, ZN => n221);
   U145 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(48));
   U146 : AOI22_X1 port map( A1 => INPUT(48), A2 => n139, B1 => INPUT(304), B2 
                           => n163, ZN => n252);
   U147 : AOI222_X1 port map( A1 => INPUT(112), A2 => n157, B1 => INPUT(240), 
                           B2 => n151, C1 => INPUT(176), C2 => n145, ZN => n251
                           );
   U148 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(47));
   U149 : AOI22_X1 port map( A1 => INPUT(47), A2 => n139, B1 => INPUT(303), B2 
                           => n163, ZN => n250);
   U150 : AOI222_X1 port map( A1 => INPUT(111), A2 => n157, B1 => INPUT(239), 
                           B2 => n151, C1 => INPUT(175), C2 => n145, ZN => n249
                           );
   U151 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(46));
   U152 : AOI22_X1 port map( A1 => INPUT(46), A2 => n139, B1 => INPUT(302), B2 
                           => n163, ZN => n248);
   U153 : AOI222_X1 port map( A1 => INPUT(110), A2 => n157, B1 => INPUT(238), 
                           B2 => n151, C1 => INPUT(174), C2 => n145, ZN => n247
                           );
   U154 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(45));
   U155 : AOI22_X1 port map( A1 => INPUT(45), A2 => n139, B1 => INPUT(301), B2 
                           => n163, ZN => n246);
   U156 : AOI222_X1 port map( A1 => INPUT(109), A2 => n157, B1 => INPUT(237), 
                           B2 => n151, C1 => INPUT(173), C2 => n145, ZN => n245
                           );
   U157 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(44));
   U158 : AOI22_X1 port map( A1 => INPUT(44), A2 => n139, B1 => INPUT(300), B2 
                           => n163, ZN => n244);
   U159 : AOI222_X1 port map( A1 => INPUT(108), A2 => n157, B1 => INPUT(236), 
                           B2 => n151, C1 => INPUT(172), C2 => n145, ZN => n243
                           );
   U160 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(43));
   U161 : AOI22_X1 port map( A1 => INPUT(43), A2 => n139, B1 => INPUT(299), B2 
                           => n163, ZN => n242);
   U162 : AOI222_X1 port map( A1 => INPUT(107), A2 => n157, B1 => INPUT(235), 
                           B2 => n151, C1 => INPUT(171), C2 => n145, ZN => n241
                           );
   U163 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(42));
   U164 : AOI22_X1 port map( A1 => INPUT(42), A2 => n139, B1 => INPUT(298), B2 
                           => n163, ZN => n240);
   U165 : AOI222_X1 port map( A1 => INPUT(106), A2 => n157, B1 => INPUT(234), 
                           B2 => n151, C1 => INPUT(170), C2 => n145, ZN => n239
                           );
   U166 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(41));
   U167 : AOI22_X1 port map( A1 => INPUT(41), A2 => n138, B1 => INPUT(297), B2 
                           => n163, ZN => n238);
   U168 : AOI222_X1 port map( A1 => INPUT(105), A2 => n156, B1 => INPUT(233), 
                           B2 => n150, C1 => INPUT(169), C2 => n144, ZN => n237
                           );
   U169 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(40));
   U170 : AOI22_X1 port map( A1 => INPUT(40), A2 => n138, B1 => INPUT(296), B2 
                           => n162, ZN => n236);
   U171 : AOI222_X1 port map( A1 => INPUT(104), A2 => n156, B1 => INPUT(232), 
                           B2 => n150, C1 => INPUT(168), C2 => n144, ZN => n235
                           );
   U172 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(39));
   U173 : AOI22_X1 port map( A1 => INPUT(39), A2 => n138, B1 => INPUT(295), B2 
                           => n162, ZN => n232);
   U174 : AOI222_X1 port map( A1 => INPUT(103), A2 => n156, B1 => INPUT(231), 
                           B2 => n150, C1 => INPUT(167), C2 => n144, ZN => n231
                           );
   U175 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(38));
   U176 : AOI22_X1 port map( A1 => INPUT(38), A2 => n138, B1 => INPUT(294), B2 
                           => n162, ZN => n230);
   U177 : AOI222_X1 port map( A1 => INPUT(102), A2 => n156, B1 => INPUT(230), 
                           B2 => n150, C1 => INPUT(166), C2 => n144, ZN => n229
                           );
   U178 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(59));
   U179 : AOI22_X1 port map( A1 => INPUT(59), A2 => n140, B1 => INPUT(315), B2 
                           => n164, ZN => n276);
   U180 : AOI222_X1 port map( A1 => INPUT(123), A2 => n158, B1 => INPUT(251), 
                           B2 => n152, C1 => INPUT(187), C2 => n146, ZN => n275
                           );
   U181 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(58));
   U182 : AOI22_X1 port map( A1 => INPUT(58), A2 => n140, B1 => INPUT(314), B2 
                           => n164, ZN => n274);
   U183 : AOI222_X1 port map( A1 => INPUT(122), A2 => n158, B1 => INPUT(250), 
                           B2 => n152, C1 => INPUT(186), C2 => n146, ZN => n273
                           );
   U184 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(57));
   U185 : AOI22_X1 port map( A1 => INPUT(57), A2 => n140, B1 => INPUT(313), B2 
                           => n164, ZN => n272);
   U186 : AOI222_X1 port map( A1 => INPUT(121), A2 => n158, B1 => INPUT(249), 
                           B2 => n152, C1 => INPUT(185), C2 => n146, ZN => n271
                           );
   U187 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(56));
   U188 : AOI22_X1 port map( A1 => INPUT(56), A2 => n140, B1 => INPUT(312), B2 
                           => n164, ZN => n270);
   U189 : AOI222_X1 port map( A1 => INPUT(120), A2 => n158, B1 => INPUT(248), 
                           B2 => n152, C1 => INPUT(184), C2 => n146, ZN => n269
                           );
   U190 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(55));
   U191 : AOI22_X1 port map( A1 => INPUT(55), A2 => n140, B1 => INPUT(311), B2 
                           => n164, ZN => n268);
   U192 : AOI222_X1 port map( A1 => INPUT(119), A2 => n158, B1 => INPUT(247), 
                           B2 => n152, C1 => INPUT(183), C2 => n146, ZN => n267
                           );
   U193 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(54));
   U194 : AOI22_X1 port map( A1 => INPUT(54), A2 => n140, B1 => INPUT(310), B2 
                           => n164, ZN => n266);
   U195 : AOI222_X1 port map( A1 => INPUT(118), A2 => n158, B1 => INPUT(246), 
                           B2 => n152, C1 => INPUT(182), C2 => n146, ZN => n265
                           );
   U196 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(53));
   U197 : AOI22_X1 port map( A1 => INPUT(53), A2 => n140, B1 => INPUT(309), B2 
                           => n164, ZN => n264);
   U198 : AOI222_X1 port map( A1 => INPUT(117), A2 => n158, B1 => INPUT(245), 
                           B2 => n152, C1 => INPUT(181), C2 => n146, ZN => n263
                           );
   U199 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(52));
   U200 : AOI22_X1 port map( A1 => INPUT(52), A2 => n139, B1 => INPUT(308), B2 
                           => n164, ZN => n262);
   U201 : AOI222_X1 port map( A1 => INPUT(116), A2 => n157, B1 => INPUT(244), 
                           B2 => n151, C1 => INPUT(180), C2 => n145, ZN => n261
                           );
   U202 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(51));
   U203 : AOI22_X1 port map( A1 => INPUT(51), A2 => n139, B1 => INPUT(307), B2 
                           => n163, ZN => n260);
   U204 : AOI222_X1 port map( A1 => INPUT(115), A2 => n157, B1 => INPUT(243), 
                           B2 => n151, C1 => INPUT(179), C2 => n145, ZN => n259
                           );
   U205 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(50));
   U206 : AOI22_X1 port map( A1 => INPUT(50), A2 => n139, B1 => INPUT(306), B2 
                           => n163, ZN => n258);
   U207 : AOI222_X1 port map( A1 => INPUT(114), A2 => n157, B1 => INPUT(242), 
                           B2 => n151, C1 => INPUT(178), C2 => n145, ZN => n257
                           );
   U208 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(49));
   U209 : AOI22_X1 port map( A1 => INPUT(49), A2 => n139, B1 => INPUT(305), B2 
                           => n163, ZN => n254);
   U210 : AOI222_X1 port map( A1 => INPUT(113), A2 => n157, B1 => INPUT(241), 
                           B2 => n151, C1 => INPUT(177), C2 => n145, ZN => n253
                           );
   U211 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(63));
   U212 : AOI22_X1 port map( A1 => INPUT(63), A2 => n140, B1 => INPUT(319), B2 
                           => n165, ZN => n286);
   U213 : AOI222_X1 port map( A1 => INPUT(127), A2 => n158, B1 => INPUT(255), 
                           B2 => n152, C1 => INPUT(191), C2 => n146, ZN => n285
                           );
   U214 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(62));
   U215 : AOI22_X1 port map( A1 => INPUT(62), A2 => n140, B1 => INPUT(318), B2 
                           => n164, ZN => n284);
   U216 : AOI222_X1 port map( A1 => INPUT(126), A2 => n158, B1 => INPUT(254), 
                           B2 => n152, C1 => INPUT(190), C2 => n146, ZN => n283
                           );
   U217 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(61));
   U218 : AOI22_X1 port map( A1 => INPUT(61), A2 => n140, B1 => INPUT(317), B2 
                           => n164, ZN => n282);
   U219 : AOI222_X1 port map( A1 => INPUT(125), A2 => n158, B1 => INPUT(253), 
                           B2 => n152, C1 => INPUT(189), C2 => n146, ZN => n281
                           );
   U220 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(60));
   U221 : AOI22_X1 port map( A1 => INPUT(60), A2 => n140, B1 => INPUT(316), B2 
                           => n164, ZN => n280);
   U222 : AOI222_X1 port map( A1 => INPUT(124), A2 => n158, B1 => INPUT(252), 
                           B2 => n152, C1 => INPUT(188), C2 => n146, ZN => n279
                           );
   U223 : CLKBUF_X1 port map( A => n293, Z => n141);
   U224 : CLKBUF_X1 port map( A => n294, Z => n147);
   U225 : CLKBUF_X1 port map( A => n295, Z => n153);
   U226 : CLKBUF_X1 port map( A => n296, Z => n159);
   U227 : CLKBUF_X1 port map( A => SEL(0), Z => n165);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_14 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_14;

architecture SYN_Behavior of Shifter_NBIT64_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_31 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_31;

architecture SYN_Behavior of Shifter_NBIT64_31 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_30 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_30;

architecture SYN_Behavior of Shifter_NBIT64_30 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_29 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_29;

architecture SYN_Behavior of Shifter_NBIT64_29 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_28 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_28;

architecture SYN_Behavior of Shifter_NBIT64_28 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_27 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_27;

architecture SYN_Behavior of Shifter_NBIT64_27 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_26 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_26;

architecture SYN_Behavior of Shifter_NBIT64_26 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_25 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_25;

architecture SYN_Behavior of Shifter_NBIT64_25 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_16_port, RESULT_1_17_port, RESULT_1_18_port, 
      RESULT_1_19_port, RESULT_1_20_port, RESULT_1_21_port, RESULT_1_22_port, 
      RESULT_1_23_port, RESULT_1_24_port, RESULT_1_25_port, RESULT_1_26_port, 
      RESULT_1_27_port, RESULT_1_28_port, RESULT_1_29_port, RESULT_1_30_port, 
      RESULT_1_31_port, RESULT_1_32_port, RESULT_1_33_port, RESULT_1_34_port, 
      RESULT_1_35_port, RESULT_1_36_port, RESULT_1_37_port, RESULT_1_38_port, 
      RESULT_1_39_port, RESULT_1_40_port, RESULT_1_41_port, RESULT_1_42_port, 
      RESULT_1_43_port, RESULT_1_44_port, RESULT_1_45_port, RESULT_1_46_port, 
      RESULT_1_47_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, RESULT_1_47_port, RESULT_1_46_port, 
      RESULT_1_45_port, RESULT_1_44_port, RESULT_1_43_port, RESULT_1_42_port, 
      RESULT_1_41_port, RESULT_1_40_port, RESULT_1_39_port, RESULT_1_38_port, 
      RESULT_1_37_port, RESULT_1_36_port, RESULT_1_35_port, RESULT_1_34_port, 
      RESULT_1_33_port, RESULT_1_32_port, RESULT_1_31_port, RESULT_1_30_port, 
      RESULT_1_29_port, RESULT_1_28_port, RESULT_1_27_port, RESULT_1_26_port, 
      RESULT_1_25_port, RESULT_1_24_port, RESULT_1_23_port, RESULT_1_22_port, 
      RESULT_1_21_port, RESULT_1_20_port, RESULT_1_19_port, RESULT_1_18_port, 
      RESULT_1_17_port, RESULT_1_16_port, TO_SHIFT(13), TO_SHIFT(12), 
      TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), TO_SHIFT(7), 
      TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), TO_SHIFT(2), 
      TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, TO_SHIFT(62), 
      TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), TO_SHIFT(57), 
      TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), TO_SHIFT(52), 
      TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), TO_SHIFT(47), 
      RESULT_1_48_port, RESULT_1_47_port, RESULT_1_46_port, RESULT_1_45_port, 
      RESULT_1_44_port, RESULT_1_43_port, RESULT_1_42_port, RESULT_1_41_port, 
      RESULT_1_40_port, RESULT_1_39_port, RESULT_1_38_port, RESULT_1_37_port, 
      RESULT_1_36_port, RESULT_1_35_port, RESULT_1_34_port, RESULT_1_33_port, 
      RESULT_1_32_port, RESULT_1_31_port, RESULT_1_30_port, RESULT_1_29_port, 
      RESULT_1_28_port, RESULT_1_27_port, RESULT_1_26_port, RESULT_1_25_port, 
      RESULT_1_24_port, RESULT_1_23_port, RESULT_1_22_port, RESULT_1_21_port, 
      RESULT_1_20_port, RESULT_1_19_port, RESULT_1_18_port, RESULT_1_17_port, 
      RESULT_1_16_port, TO_SHIFT(13), TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10),
      TO_SHIFT(9), TO_SHIFT(8), TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), 
      TO_SHIFT(4), TO_SHIFT(3), TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : CLKBUF_X1 port map( A => TO_SHIFT(14), Z => RESULT_1_16_port);
   U3 : CLKBUF_X1 port map( A => TO_SHIFT(19), Z => RESULT_1_21_port);
   U4 : CLKBUF_X1 port map( A => TO_SHIFT(20), Z => RESULT_1_22_port);
   U5 : CLKBUF_X1 port map( A => TO_SHIFT(21), Z => RESULT_1_23_port);
   U6 : CLKBUF_X1 port map( A => TO_SHIFT(22), Z => RESULT_1_24_port);
   U7 : CLKBUF_X1 port map( A => TO_SHIFT(23), Z => RESULT_1_25_port);
   U8 : CLKBUF_X1 port map( A => TO_SHIFT(27), Z => RESULT_1_29_port);
   U9 : CLKBUF_X1 port map( A => TO_SHIFT(28), Z => RESULT_1_30_port);
   U10 : CLKBUF_X1 port map( A => TO_SHIFT(17), Z => RESULT_1_19_port);
   U11 : CLKBUF_X1 port map( A => TO_SHIFT(18), Z => RESULT_1_20_port);
   U12 : CLKBUF_X1 port map( A => TO_SHIFT(16), Z => RESULT_1_18_port);
   U13 : CLKBUF_X1 port map( A => TO_SHIFT(15), Z => RESULT_1_17_port);
   U14 : CLKBUF_X1 port map( A => TO_SHIFT(24), Z => RESULT_1_26_port);
   U15 : CLKBUF_X1 port map( A => TO_SHIFT(29), Z => RESULT_1_31_port);
   U16 : CLKBUF_X1 port map( A => TO_SHIFT(30), Z => RESULT_1_32_port);
   U17 : BUF_X1 port map( A => TO_SHIFT(40), Z => RESULT_1_42_port);
   U18 : BUF_X1 port map( A => TO_SHIFT(31), Z => RESULT_1_33_port);
   U19 : BUF_X1 port map( A => TO_SHIFT(32), Z => RESULT_1_34_port);
   U20 : BUF_X1 port map( A => TO_SHIFT(33), Z => RESULT_1_35_port);
   U21 : BUF_X1 port map( A => TO_SHIFT(34), Z => RESULT_1_36_port);
   U22 : BUF_X1 port map( A => TO_SHIFT(35), Z => RESULT_1_37_port);
   U23 : BUF_X1 port map( A => TO_SHIFT(36), Z => RESULT_1_38_port);
   U24 : BUF_X1 port map( A => TO_SHIFT(37), Z => RESULT_1_39_port);
   U25 : BUF_X1 port map( A => TO_SHIFT(38), Z => RESULT_1_40_port);
   U26 : BUF_X1 port map( A => TO_SHIFT(39), Z => RESULT_1_41_port);
   U27 : BUF_X1 port map( A => TO_SHIFT(41), Z => RESULT_1_43_port);
   U28 : BUF_X1 port map( A => TO_SHIFT(44), Z => RESULT_1_46_port);
   U29 : BUF_X1 port map( A => TO_SHIFT(45), Z => RESULT_1_47_port);
   U30 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);
   U31 : BUF_X1 port map( A => TO_SHIFT(42), Z => RESULT_1_44_port);
   U32 : BUF_X1 port map( A => TO_SHIFT(43), Z => RESULT_1_45_port);
   U33 : CLKBUF_X1 port map( A => TO_SHIFT(25), Z => RESULT_1_27_port);
   U34 : CLKBUF_X1 port map( A => TO_SHIFT(26), Z => RESULT_1_28_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_24 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_24;

architecture SYN_Behavior of Shifter_NBIT64_24 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_23 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_23;

architecture SYN_Behavior of Shifter_NBIT64_23 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_22 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_22;

architecture SYN_Behavior of Shifter_NBIT64_22 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_21 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_21;

architecture SYN_Behavior of Shifter_NBIT64_21 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_20 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_20;

architecture SYN_Behavior of Shifter_NBIT64_20 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_19 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_19;

architecture SYN_Behavior of Shifter_NBIT64_19 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_18 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_18;

architecture SYN_Behavior of Shifter_NBIT64_18 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_17 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_17;

architecture SYN_Behavior of Shifter_NBIT64_17 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_13 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_13;

architecture SYN_Behavior of Shifter_NBIT64_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_12 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_12;

architecture SYN_Behavior of Shifter_NBIT64_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_11 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_11;

architecture SYN_Behavior of Shifter_NBIT64_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_10 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_10;

architecture SYN_Behavior of Shifter_NBIT64_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_9 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_9;

architecture SYN_Behavior of Shifter_NBIT64_9 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_16_port, RESULT_1_17_port, RESULT_1_18_port, 
      RESULT_1_19_port, RESULT_1_20_port, RESULT_1_21_port, RESULT_1_22_port, 
      RESULT_1_23_port, RESULT_1_24_port, RESULT_1_25_port, RESULT_1_26_port, 
      RESULT_1_27_port, RESULT_1_28_port, RESULT_1_29_port, RESULT_1_30_port, 
      RESULT_1_31_port, RESULT_1_32_port, RESULT_1_33_port, RESULT_1_34_port, 
      RESULT_1_35_port, RESULT_1_36_port, RESULT_1_37_port, RESULT_1_38_port, 
      RESULT_1_39_port, RESULT_1_40_port, RESULT_1_41_port, RESULT_1_42_port, 
      RESULT_1_43_port, RESULT_1_44_port, RESULT_1_45_port, RESULT_1_46_port, 
      RESULT_1_47_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, RESULT_1_47_port, RESULT_1_46_port, 
      RESULT_1_45_port, RESULT_1_44_port, RESULT_1_43_port, RESULT_1_42_port, 
      RESULT_1_41_port, RESULT_1_40_port, RESULT_1_39_port, RESULT_1_38_port, 
      RESULT_1_37_port, RESULT_1_36_port, RESULT_1_35_port, RESULT_1_34_port, 
      RESULT_1_33_port, RESULT_1_32_port, RESULT_1_31_port, RESULT_1_30_port, 
      RESULT_1_29_port, RESULT_1_28_port, RESULT_1_27_port, RESULT_1_26_port, 
      RESULT_1_25_port, RESULT_1_24_port, RESULT_1_23_port, RESULT_1_22_port, 
      RESULT_1_21_port, RESULT_1_20_port, RESULT_1_19_port, RESULT_1_18_port, 
      RESULT_1_17_port, RESULT_1_16_port, TO_SHIFT(13), TO_SHIFT(12), 
      TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), TO_SHIFT(7), 
      TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), TO_SHIFT(2), 
      TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, TO_SHIFT(62), 
      TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), TO_SHIFT(57), 
      TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), TO_SHIFT(52), 
      TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), TO_SHIFT(47), 
      RESULT_1_48_port, RESULT_1_47_port, RESULT_1_46_port, RESULT_1_45_port, 
      RESULT_1_44_port, RESULT_1_43_port, RESULT_1_42_port, RESULT_1_41_port, 
      RESULT_1_40_port, RESULT_1_39_port, RESULT_1_38_port, RESULT_1_37_port, 
      RESULT_1_36_port, RESULT_1_35_port, RESULT_1_34_port, RESULT_1_33_port, 
      RESULT_1_32_port, RESULT_1_31_port, RESULT_1_30_port, RESULT_1_29_port, 
      RESULT_1_28_port, RESULT_1_27_port, RESULT_1_26_port, RESULT_1_25_port, 
      RESULT_1_24_port, RESULT_1_23_port, RESULT_1_22_port, RESULT_1_21_port, 
      RESULT_1_20_port, RESULT_1_19_port, RESULT_1_18_port, RESULT_1_17_port, 
      RESULT_1_16_port, TO_SHIFT(13), TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10),
      TO_SHIFT(9), TO_SHIFT(8), TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), 
      TO_SHIFT(4), TO_SHIFT(3), TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : CLKBUF_X1 port map( A => TO_SHIFT(23), Z => RESULT_1_25_port);
   U3 : CLKBUF_X1 port map( A => TO_SHIFT(24), Z => RESULT_1_26_port);
   U4 : CLKBUF_X1 port map( A => TO_SHIFT(25), Z => RESULT_1_27_port);
   U5 : CLKBUF_X1 port map( A => TO_SHIFT(26), Z => RESULT_1_28_port);
   U6 : CLKBUF_X1 port map( A => TO_SHIFT(27), Z => RESULT_1_29_port);
   U7 : CLKBUF_X1 port map( A => TO_SHIFT(28), Z => RESULT_1_30_port);
   U8 : CLKBUF_X1 port map( A => TO_SHIFT(37), Z => RESULT_1_39_port);
   U9 : CLKBUF_X1 port map( A => TO_SHIFT(39), Z => RESULT_1_41_port);
   U10 : CLKBUF_X1 port map( A => TO_SHIFT(41), Z => RESULT_1_43_port);
   U11 : CLKBUF_X1 port map( A => TO_SHIFT(43), Z => RESULT_1_45_port);
   U12 : CLKBUF_X1 port map( A => TO_SHIFT(29), Z => RESULT_1_31_port);
   U13 : CLKBUF_X1 port map( A => TO_SHIFT(30), Z => RESULT_1_32_port);
   U14 : CLKBUF_X1 port map( A => TO_SHIFT(31), Z => RESULT_1_33_port);
   U15 : CLKBUF_X1 port map( A => TO_SHIFT(32), Z => RESULT_1_34_port);
   U16 : CLKBUF_X1 port map( A => TO_SHIFT(33), Z => RESULT_1_35_port);
   U17 : CLKBUF_X1 port map( A => TO_SHIFT(34), Z => RESULT_1_36_port);
   U18 : CLKBUF_X1 port map( A => TO_SHIFT(35), Z => RESULT_1_37_port);
   U19 : CLKBUF_X1 port map( A => TO_SHIFT(36), Z => RESULT_1_38_port);
   U20 : CLKBUF_X1 port map( A => TO_SHIFT(38), Z => RESULT_1_40_port);
   U21 : CLKBUF_X1 port map( A => TO_SHIFT(40), Z => RESULT_1_42_port);
   U22 : CLKBUF_X1 port map( A => TO_SHIFT(42), Z => RESULT_1_44_port);
   U23 : CLKBUF_X1 port map( A => TO_SHIFT(44), Z => RESULT_1_46_port);
   U24 : CLKBUF_X1 port map( A => TO_SHIFT(45), Z => RESULT_1_47_port);
   U25 : CLKBUF_X1 port map( A => TO_SHIFT(15), Z => RESULT_1_17_port);
   U26 : CLKBUF_X1 port map( A => TO_SHIFT(17), Z => RESULT_1_19_port);
   U27 : CLKBUF_X1 port map( A => TO_SHIFT(18), Z => RESULT_1_20_port);
   U28 : CLKBUF_X1 port map( A => TO_SHIFT(19), Z => RESULT_1_21_port);
   U29 : CLKBUF_X1 port map( A => TO_SHIFT(20), Z => RESULT_1_22_port);
   U30 : CLKBUF_X1 port map( A => TO_SHIFT(21), Z => RESULT_1_23_port);
   U31 : CLKBUF_X1 port map( A => TO_SHIFT(22), Z => RESULT_1_24_port);
   U32 : CLKBUF_X1 port map( A => TO_SHIFT(16), Z => RESULT_1_18_port);
   U33 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);
   U34 : CLKBUF_X1 port map( A => TO_SHIFT(14), Z => RESULT_1_16_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_8 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_8;

architecture SYN_Behavior of Shifter_NBIT64_8 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_7 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_7;

architecture SYN_Behavior of Shifter_NBIT64_7 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_6 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_6;

architecture SYN_Behavior of Shifter_NBIT64_6 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_5 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_5;

architecture SYN_Behavior of Shifter_NBIT64_5 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_4 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_4;

architecture SYN_Behavior of Shifter_NBIT64_4 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_3 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_3;

architecture SYN_Behavior of Shifter_NBIT64_3 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_2 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_2;

architecture SYN_Behavior of Shifter_NBIT64_2 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_1 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_1;

architecture SYN_Behavior of Shifter_NBIT64_1 is

signal X_Logic0_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), TO_SHIFT(46), TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43), 
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_15 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_15;

architecture SYN_Behavior of Booth_Encoder_15 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n11, n12 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n5);
   U2 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n6);
   U3 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n8, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n8);
   U5 : INV_X1 port map( A => B(2), ZN => n9);
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n11);
   U7 : OAI22_X1 port map( A1 => n7, A2 => n9, B1 => B(2), B2 => n5, ZN => 
                           OUT_TO_MUX(1));
   U8 : AND3_X1 port map( A1 => B(2), A2 => n8, A3 => n7, ZN => OUT_TO_MUX(2));
   U9 : AOI21_X1 port map( B1 => n12, B2 => n6, A => B(2), ZN => OUT_TO_MUX(0))
                           ;
   U10 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n11, ZN => n12);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_14 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_14;

architecture SYN_Behavior of Booth_Encoder_14 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U2 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U3 : INV_X1 port map( A => B(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);
   U6 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_13 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_13;

architecture SYN_Behavior of Booth_Encoder_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U2 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U3 : INV_X1 port map( A => B(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_12 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_12;

architecture SYN_Behavior of Booth_Encoder_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U2 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U3 : INV_X1 port map( A => B(2), ZN => n5);
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_11 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_11;

architecture SYN_Behavior of Booth_Encoder_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_10 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_10;

architecture SYN_Behavior of Booth_Encoder_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_9 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_9;

architecture SYN_Behavior of Booth_Encoder_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_8 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_8;

architecture SYN_Behavior of Booth_Encoder_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_7 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_7;

architecture SYN_Behavior of Booth_Encoder_7 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U2 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U3 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);
   U4 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U5 : INV_X1 port map( A => B(2), ZN => n5);
   U6 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_6 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_6;

architecture SYN_Behavior of Booth_Encoder_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_5 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_5;

architecture SYN_Behavior of Booth_Encoder_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_4 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_4;

architecture SYN_Behavior of Booth_Encoder_4 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);
   U6 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_3 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_3;

architecture SYN_Behavior of Booth_Encoder_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_2 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_2;

architecture SYN_Behavior of Booth_Encoder_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));
   U6 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_1 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_1;

architecture SYN_Behavior of Booth_Encoder_1 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           OUT_TO_MUX(1));
   U2 : INV_X1 port map( A => B(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => B(2), ZN => OUT_TO_MUX(0));
   U4 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n7, ZN => n8);
   U5 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n7);
   U6 : AND3_X1 port map( A1 => B(2), A2 => n7, A3 => n8, ZN => OUT_TO_MUX(2));

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_1_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_1_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_1_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_34_port, carry_33_port, carry_32_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, net25644, net25636, net25623, net25602, 
      net25575, net25574, net25571, net25566, net25478, net25448, net25573, 
      net25572, net47167, net47226, net47230, net25560, net49388, net49501, 
      net51391, net49514, net25606, net61027, net61048, net68328, net70121, 
      net70219, net70303, net70406, net75030, net25463, net25461, net47224, 
      net25614, net25468, net25467, net84851, net25570, net25568, net70449, 
      net25625, net25605, net25601, net25600, net25564, net25563, net25474, 
      net25473, net25472, net25471, net25466, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206 : std_logic;

begin
   
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1 : CLKBUF_X1 port map( A => n55, Z => n1);
   U2 : NAND2_X1 port map( A1 => B(56), A2 => n55, ZN => n2);
   U3 : NAND2_X1 port map( A1 => B(56), A2 => n55, ZN => n3);
   U4 : CLKBUF_X1 port map( A => n23, Z => n4);
   U5 : CLKBUF_X1 port map( A => A(61), Z => net70406);
   U6 : INV_X1 port map( A => A(41), ZN => n90);
   U7 : INV_X1 port map( A => A(44), ZN => n101);
   U8 : INV_X1 port map( A => B(63), ZN => net25568);
   U9 : XNOR2_X1 port map( A => n186, B => n67, ZN => SUM(35));
   U10 : INV_X1 port map( A => B(35), ZN => n151);
   U11 : XNOR2_X1 port map( A => n185, B => n71, ZN => SUM(36));
   U12 : INV_X1 port map( A => B(36), ZN => n152);
   U13 : INV_X1 port map( A => B(37), ZN => n153);
   U14 : INV_X1 port map( A => B(40), ZN => n154);
   U15 : XNOR2_X1 port map( A => n180, B => n90, ZN => SUM(41));
   U16 : INV_X1 port map( A => B(41), ZN => n155);
   U17 : XNOR2_X1 port map( A => A(42), B => n179, ZN => SUM(42));
   U18 : XNOR2_X1 port map( A => n177, B => n101, ZN => SUM(44));
   U19 : INV_X1 port map( A => B(44), ZN => n156);
   U20 : INV_X1 port map( A => B(45), ZN => n157);
   U21 : XNOR2_X1 port map( A => A(46), B => n175, ZN => SUM(46));
   U22 : INV_X1 port map( A => B(48), ZN => n158);
   U23 : XNOR2_X1 port map( A => n61, B => n159, ZN => n172);
   U24 : INV_X1 port map( A => B(49), ZN => n159);
   U25 : INV_X1 port map( A => B(52), ZN => n160);
   U26 : INV_X1 port map( A => B(53), ZN => n161);
   U27 : XNOR2_X1 port map( A => B(54), B => n188, ZN => n167);
   U28 : INV_X1 port map( A => B(56), ZN => n162);
   U29 : INV_X1 port map( A => B(57), ZN => n163);
   U30 : XNOR2_X1 port map( A => B(59), B => n22, ZN => net25574);
   U31 : INV_X1 port map( A => B(61), ZN => net25560);
   U32 : NAND2_X1 port map( A1 => B(63), A2 => net49388, ZN => net25478);
   U33 : NAND2_X1 port map( A1 => net25478, A2 => n150, ZN => SUM(64));
   U34 : XNOR2_X1 port map( A => n164, B => n148, ZN => SUM(57));
   U35 : BUF_X1 port map( A => net84851, Z => net51391);
   U36 : BUF_X1 port map( A => net25625, Z => net49514);
   U37 : NOR2_X1 port map( A1 => n111, A2 => B(48), ZN => n5);
   U38 : NOR2_X1 port map( A1 => n133, A2 => B(54), ZN => n6);
   U39 : OAI211_X1 port map( C1 => n19, C2 => net75030, A => n20, B => n7, ZN 
                           => n8);
   U40 : INV_X1 port map( A => B(59), ZN => n7);
   U41 : INV_X1 port map( A => n8, ZN => net25461);
   U42 : OAI21_X1 port map( B1 => net25473, B2 => net25472, A => net25474, ZN 
                           => net25471);
   U43 : NOR2_X1 port map( A1 => net25471, A2 => B(62), ZN => net25563);
   U44 : NOR2_X1 port map( A1 => B(61), A2 => net25466, ZN => net25472);
   U45 : INV_X1 port map( A => A(61), ZN => net25473);
   U46 : OAI21_X1 port map( B1 => net25473, B2 => net25625, A => net25474, ZN 
                           => net25605);
   U47 : NAND2_X1 port map( A1 => net25466, A2 => B(61), ZN => net25474);
   U48 : CLKBUF_X1 port map( A => net25474, Z => net70121);
   U49 : NOR2_X1 port map( A1 => B(61), A2 => net84851, ZN => net25625);
   U50 : NAND2_X1 port map( A1 => net25467, A2 => net25468, ZN => net25466);
   U51 : NAND2_X1 port map( A1 => net25468, A2 => net25467, ZN => net84851);
   U52 : OAI21_X1 port map( B1 => net25563, B2 => net25564, A => net25600, ZN 
                           => net25601);
   U53 : XNOR2_X1 port map( A => net25601, B => net25568, ZN => net25570);
   U54 : INV_X1 port map( A => A(62), ZN => net25564);
   U55 : CLKBUF_X1 port map( A => net25564, Z => net25644);
   U56 : CLKBUF_X1 port map( A => net25563, Z => net70449);
   U57 : NAND2_X1 port map( A1 => net25605, A2 => B(62), ZN => net25600);
   U58 : OAI21_X1 port map( B1 => net70303, B2 => net70449, A => net25600, ZN 
                           => net70219);
   U59 : XNOR2_X1 port map( A => net25606, B => B(62), ZN => net25571);
   U60 : XNOR2_X1 port map( A => net25570, B => net47226, ZN => SUM(63));
   U61 : NAND2_X1 port map( A1 => net25566, A2 => net25568, ZN => net25602);
   U62 : CLKBUF_X1 port map( A => n144, Z => n12);
   U63 : OAI21_X1 port map( B1 => n5, B2 => n116, A => n117, ZN => n9);
   U64 : NOR2_X1 port map( A1 => n81, A2 => B(40), ZN => n10);
   U65 : XNOR2_X1 port map( A => n172, B => n120, ZN => SUM(49));
   U66 : OAI21_X1 port map( B1 => n10, B2 => n86, A => n87, ZN => n11);
   U67 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n84);
   U68 : CLKBUF_X1 port map( A => A(34), Z => n13);
   U69 : XNOR2_X1 port map( A => n176, B => n105, ZN => SUM(45));
   U70 : NOR2_X1 port map( A1 => n73, A2 => B(38), ZN => n14);
   U71 : OAI21_X1 port map( B1 => n137, B2 => B(55), A => A(55), ZN => n15);
   U72 : CLKBUF_X1 port map( A => n200, Z => n16);
   U73 : OAI21_X1 port map( B1 => n17, B2 => B(60), A => A(60), ZN => net25468)
                           ;
   U74 : OAI21_X1 port map( B1 => net25461, B2 => n18, A => net25463, ZN => n17
                           );
   U75 : INV_X1 port map( A => A(59), ZN => n18);
   U76 : CLKBUF_X1 port map( A => n18, Z => net68328);
   U77 : OAI21_X1 port map( B1 => net25461, B2 => n18, A => net25463, ZN => 
                           net25614);
   U78 : NAND2_X1 port map( A1 => net25614, A2 => B(60), ZN => net25467);
   U79 : XNOR2_X1 port map( A => B(60), B => net47224, ZN => net25573);
   U80 : CLKBUF_X1 port map( A => A(60), Z => net47167);
   U81 : CLKBUF_X1 port map( A => net25614, Z => net47224);
   U82 : OAI21_X1 port map( B1 => n23, B2 => net75030, A => n20, ZN => n21);
   U83 : NOR2_X1 port map( A1 => B(58), A2 => net25448, ZN => n19);
   U84 : NAND2_X1 port map( A1 => B(59), A2 => n21, ZN => net25463);
   U85 : CLKBUF_X1 port map( A => n20, Z => n24);
   U86 : INV_X1 port map( A => A(58), ZN => net75030);
   U87 : NAND2_X1 port map( A1 => net25448, A2 => B(58), ZN => n20);
   U88 : XNOR2_X1 port map( A => B(58), B => net25623, ZN => net25575);
   U89 : NOR2_X1 port map( A1 => B(58), A2 => net61027, ZN => n23);
   U90 : OAI21_X1 port map( B1 => net75030, B2 => n4, A => n24, ZN => n22);
   U91 : NOR2_X1 port map( A1 => B(44), A2 => n96, ZN => n25);
   U92 : CLKBUF_X1 port map( A => n99, Z => n26);
   U93 : CLKBUF_X1 port map( A => n196, Z => n27);
   U94 : NOR2_X1 port map( A1 => B(50), A2 => n118, ZN => n28);
   U95 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n2, ZN => n29);
   U96 : CLKBUF_X1 port map( A => n195, Z => n30);
   U97 : NOR2_X1 port map( A1 => B(36), A2 => n65, ZN => n31);
   U98 : BUF_X1 port map( A => n201, Z => n32);
   U99 : OAI21_X1 port map( B1 => n31, B2 => n71, A => n72, ZN => n33);
   U100 : XNOR2_X1 port map( A => n169, B => n131, ZN => SUM(52));
   U101 : CLKBUF_X1 port map( A => n111, Z => n34);
   U102 : CLKBUF_X1 port map( A => n192, Z => n35);
   U103 : CLKBUF_X1 port map( A => n103, Z => n36);
   U104 : CLKBUF_X1 port map( A => n197, Z => n37);
   U105 : CLKBUF_X1 port map( A => n193, Z => n38);
   U106 : XNOR2_X1 port map( A => A(38), B => n183, ZN => SUM(38));
   U107 : XNOR2_X1 port map( A => n173, B => n116, ZN => SUM(48));
   U108 : XNOR2_X1 port map( A => n181, B => n86, ZN => SUM(40));
   U109 : XNOR2_X1 port map( A => net25571, B => net25636, ZN => SUM(62));
   U110 : CLKBUF_X1 port map( A => n81, Z => n39);
   U111 : NOR2_X1 port map( A1 => n88, A2 => B(42), ZN => n40);
   U112 : NOR2_X1 port map( A1 => n204, A2 => B(45), ZN => n41);
   U113 : NOR2_X1 port map( A1 => n141, A2 => B(56), ZN => n42);
   U114 : OAI21_X1 port map( B1 => n122, B2 => B(51), A => A(51), ZN => n43);
   U115 : CLKBUF_X1 port map( A => n190, Z => n44);
   U116 : INV_X1 port map( A => A(45), ZN => n105);
   U117 : XNOR2_X1 port map( A => n165, B => n146, ZN => SUM(56));
   U118 : XNOR2_X1 port map( A => A(39), B => n182, ZN => SUM(39));
   U119 : XNOR2_X1 port map( A => n168, B => n135, ZN => SUM(53));
   U120 : INV_X1 port map( A => A(53), ZN => n135);
   U121 : INV_X1 port map( A => A(48), ZN => n116);
   U122 : NAND2_X1 port map( A1 => B(56), A2 => n55, ZN => n45);
   U123 : INV_X1 port map( A => n139, ZN => n46);
   U124 : CLKBUF_X1 port map( A => A(55), Z => n47);
   U125 : INV_X1 port map( A => A(36), ZN => n71);
   U126 : INV_X1 port map( A => A(52), ZN => n131);
   U127 : NAND2_X1 port map( A1 => n127, A2 => n43, ZN => n48);
   U128 : CLKBUF_X1 port map( A => A(47), Z => n49);
   U129 : INV_X1 port map( A => A(49), ZN => n120);
   U130 : INV_X1 port map( A => A(38), ZN => n79);
   U131 : CLKBUF_X1 port map( A => A(51), Z => n50);
   U132 : CLKBUF_X1 port map( A => n136, Z => n51);
   U133 : CLKBUF_X1 port map( A => n96, Z => n52);
   U134 : NOR2_X1 port map( A1 => n33, A2 => B(37), ZN => n53);
   U135 : NOR2_X1 port map( A1 => B(35), A2 => n62, ZN => n54);
   U136 : CLKBUF_X1 port map( A => net25644, Z => net70303);
   U137 : XNOR2_X1 port map( A => B(50), B => n44, ZN => n171);
   U138 : NAND2_X1 port map( A1 => n142, A2 => n15, ZN => n55);
   U139 : NOR2_X1 port map( A1 => B(46), A2 => n191, ZN => n56);
   U140 : NOR2_X1 port map( A1 => n84, A2 => B(41), ZN => n57);
   U141 : NOR2_X1 port map( A1 => B(52), A2 => n48, ZN => n58);
   U142 : NOR2_X1 port map( A1 => n144, A2 => B(57), ZN => n59);
   U143 : CLKBUF_X1 port map( A => n62, Z => n60);
   U144 : XNOR2_X1 port map( A => n39, B => n154, ZN => n181);
   U145 : XNOR2_X1 port map( A => B(34), B => carry_34_port, ZN => n187);
   U146 : XNOR2_X1 port map( A => n184, B => n75, ZN => SUM(37));
   U147 : XNOR2_X1 port map( A => n60, B => n151, ZN => n186);
   U148 : INV_X1 port map( A => A(35), ZN => n67);
   U149 : XNOR2_X1 port map( A => n48, B => n160, ZN => n169);
   U150 : NAND2_X1 port map( A1 => B(52), A2 => n126, ZN => n132);
   U151 : INV_X1 port map( A => A(37), ZN => n75);
   U152 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => n126);
   U153 : INV_X1 port map( A => A(46), ZN => n109);
   U154 : INV_X1 port map( A => net68328, ZN => net61048);
   U155 : CLKBUF_X1 port map( A => n9, Z => n61);
   U156 : INV_X1 port map( A => A(42), ZN => n94);
   U157 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => n63);
   U158 : OAI21_X1 port map( B1 => A(34), B2 => B(34), A => carry_34_port, ZN 
                           => n64);
   U159 : XNOR2_X1 port map( A => n13, B => n187, ZN => SUM(34));
   U160 : XNOR2_X1 port map( A => A(43), B => n178, ZN => SUM(43));
   U161 : OAI21_X1 port map( B1 => n59, B2 => n148, A => n149, ZN => net61027);
   U162 : XNOR2_X1 port map( A => n50, B => n170, ZN => SUM(51));
   U163 : XNOR2_X1 port map( A => n34, B => n158, ZN => n173);
   U164 : NAND2_X1 port map( A1 => B(48), A2 => n111, ZN => n117);
   U165 : INV_X1 port map( A => A(56), ZN => n146);
   U166 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n111);
   U167 : OAI21_X1 port map( B1 => net47230, B2 => net49514, A => net70121, ZN 
                           => net25606);
   U168 : INV_X1 port map( A => net70406, ZN => net47230);
   U169 : XNOR2_X1 port map( A => net61048, B => net25574, ZN => SUM(59));
   U170 : INV_X1 port map( A => net75030, ZN => net49501);
   U171 : XNOR2_X1 port map( A => n49, B => n174, ZN => SUM(47));
   U172 : NAND2_X1 port map( A1 => B(44), A2 => n96, ZN => n102);
   U173 : XNOR2_X1 port map( A => n52, B => n156, ZN => n177);
   U174 : XNOR2_X1 port map( A => n46, B => n167, ZN => SUM(54));
   U175 : INV_X1 port map( A => A(54), ZN => n139);
   U176 : XNOR2_X1 port map( A => n1, B => n162, ZN => n165);
   U177 : XNOR2_X1 port map( A => net49501, B => net25575, ZN => SUM(58));
   U178 : CLKBUF_X1 port map( A => A(63), Z => net49388);
   U179 : INV_X1 port map( A => A(57), ZN => n148);
   U180 : XNOR2_X1 port map( A => A(50), B => n171, ZN => SUM(50));
   U181 : XNOR2_X1 port map( A => n202, B => n161, ZN => n168);
   U182 : NAND2_X1 port map( A1 => n142, A2 => n143, ZN => n141);
   U183 : INV_X1 port map( A => A(50), ZN => n124);
   U184 : XNOR2_X1 port map( A => net51391, B => net25560, ZN => net25572);
   U185 : OAI21_X1 port map( B1 => n122, B2 => B(51), A => A(51), ZN => n128);
   U186 : INV_X1 port map( A => A(63), ZN => net47226);
   U187 : NAND2_X1 port map( A1 => n195, A2 => B(51), ZN => n127);
   U188 : XNOR2_X1 port map( A => B(51), B => n30, ZN => n170);
   U189 : XNOR2_X1 port map( A => net25572, B => net47230, ZN => SUM(61));
   U190 : XNOR2_X1 port map( A => n47, B => n166, ZN => SUM(55));
   U191 : OAI21_X1 port map( B1 => n194, B2 => B(55), A => A(55), ZN => n143);
   U192 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n62);
   U193 : NAND2_X1 port map( A1 => B(54), A2 => n189, ZN => n140);
   U194 : NAND2_X1 port map( A1 => n190, A2 => B(50), ZN => n125);
   U195 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => n96);
   U196 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => n81);
   U197 : XNOR2_X1 port map( A => net47167, B => net25573, ZN => SUM(60));
   U198 : NOR2_X1 port map( A1 => n202, A2 => B(53), ZN => n134);
   U199 : OAI21_X1 port map( B1 => n135, B2 => n134, A => n136, ZN => n133);
   U200 : OAI21_X1 port map( B1 => n32, B2 => n135, A => n51, ZN => n188);
   U201 : OAI21_X1 port map( B1 => n201, B2 => n135, A => n136, ZN => n189);
   U202 : NOR2_X1 port map( A1 => n114, A2 => B(49), ZN => n119);
   U203 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n118);
   U204 : OAI21_X1 port map( B1 => n203, B2 => n120, A => n121, ZN => n190);
   U205 : OAI21_X1 port map( B1 => n41, B2 => n105, A => n106, ZN => n103);
   U206 : NAND2_X1 port map( A1 => n191, A2 => B(46), ZN => n110);
   U207 : XNOR2_X1 port map( A => B(46), B => n36, ZN => n175);
   U208 : NOR2_X1 port map( A1 => n103, A2 => B(46), ZN => n108);
   U209 : NOR2_X1 port map( A1 => n204, A2 => B(45), ZN => n104);
   U210 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n191);
   U211 : OAI21_X1 port map( B1 => n57, B2 => n90, A => n91, ZN => n88);
   U212 : NAND2_X1 port map( A1 => B(42), A2 => n192, ZN => n95);
   U213 : XNOR2_X1 port map( A => B(42), B => n35, ZN => n179);
   U214 : NOR2_X1 port map( A1 => n88, A2 => B(42), ZN => n93);
   U215 : NOR2_X1 port map( A1 => n84, A2 => B(41), ZN => n89);
   U216 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n192);
   U217 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n73);
   U218 : NAND2_X1 port map( A1 => n193, A2 => B(38), ZN => n80);
   U219 : XNOR2_X1 port map( A => B(38), B => n38, ZN => n183);
   U220 : NOR2_X1 port map( A1 => n73, A2 => B(38), ZN => n78);
   U221 : NOR2_X1 port map( A1 => n69, A2 => B(37), ZN => n74);
   U222 : OAI21_X1 port map( B1 => n53, B2 => n75, A => n76, ZN => n193);
   U223 : NOR2_X1 port map( A1 => n133, A2 => B(54), ZN => n138);
   U224 : OAI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n137);
   U225 : OAI21_X1 port map( B1 => n6, B2 => n139, A => n140, ZN => n194);
   U226 : NOR2_X1 port map( A1 => n118, A2 => B(50), ZN => n123);
   U227 : OAI21_X1 port map( B1 => n124, B2 => n123, A => n125, ZN => n122);
   U228 : OAI21_X1 port map( B1 => n28, B2 => n124, A => n125, ZN => n195);
   U229 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n107);
   U230 : NAND2_X1 port map( A1 => B(47), A2 => n196, ZN => n112);
   U231 : OAI21_X1 port map( B1 => n107, B2 => B(47), A => A(47), ZN => n113);
   U232 : XNOR2_X1 port map( A => B(47), B => n27, ZN => n174);
   U233 : OAI21_X1 port map( B1 => n56, B2 => n109, A => n110, ZN => n196);
   U234 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n92);
   U235 : NAND2_X1 port map( A1 => B(43), A2 => n197, ZN => n97);
   U236 : OAI21_X1 port map( B1 => n92, B2 => B(43), A => A(43), ZN => n98);
   U237 : XNOR2_X1 port map( A => B(43), B => n37, ZN => n178);
   U238 : OAI21_X1 port map( B1 => n40, B2 => n94, A => n95, ZN => n197);
   U239 : OAI21_X1 port map( B1 => n14, B2 => n79, A => n80, ZN => n77);
   U240 : NAND2_X1 port map( A1 => B(39), A2 => n198, ZN => n82);
   U241 : OAI21_X1 port map( B1 => n77, B2 => B(39), A => A(39), ZN => n83);
   U242 : XNOR2_X1 port map( A => B(39), B => n198, ZN => n182);
   U243 : OAI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n198);
   U244 : OAI21_X1 port map( B1 => n42, B2 => n146, A => n45, ZN => n144);
   U245 : XNOR2_X1 port map( A => n12, B => n163, ZN => n164);
   U246 : NAND2_X1 port map( A1 => n29, A2 => B(57), ZN => n149);
   U247 : NOR2_X1 port map( A1 => n199, A2 => B(57), ZN => n147);
   U248 : NOR2_X1 port map( A1 => n141, A2 => B(56), ZN => n145);
   U249 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n3, ZN => n199);
   U250 : OAI21_X1 port map( B1 => n54, B2 => n67, A => n68, ZN => n65);
   U251 : XNOR2_X1 port map( A => n16, B => n152, ZN => n185);
   U252 : NAND2_X1 port map( A1 => n200, A2 => B(36), ZN => n72);
   U253 : NOR2_X1 port map( A1 => n65, A2 => B(36), ZN => n70);
   U254 : NOR2_X1 port map( A1 => B(35), A2 => n62, ZN => n66);
   U255 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n200);
   U256 : OAI21_X1 port map( B1 => n147, B2 => n148, A => n149, ZN => net25448)
                           ;
   U257 : CLKBUF_X1 port map( A => net61027, Z => net25623);
   U258 : NOR2_X1 port map( A1 => n129, A2 => B(53), ZN => n201);
   U259 : NOR2_X1 port map( A1 => B(52), A2 => n126, ZN => n130);
   U260 : OAI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => n129);
   U261 : OAI21_X1 port map( B1 => n58, B2 => n131, A => n132, ZN => n202);
   U262 : NAND2_X1 port map( A1 => n129, A2 => B(53), ZN => n136);
   U263 : NOR2_X1 port map( A1 => B(49), A2 => n9, ZN => n203);
   U264 : NOR2_X1 port map( A1 => n111, A2 => B(48), ZN => n115);
   U265 : OAI21_X1 port map( B1 => n115, B2 => n116, A => n117, ZN => n114);
   U266 : NAND2_X1 port map( A1 => n114, A2 => B(49), ZN => n121);
   U267 : OAI21_X1 port map( B1 => n25, B2 => n101, A => n102, ZN => n99);
   U268 : XNOR2_X1 port map( A => n26, B => n157, ZN => n176);
   U269 : NAND2_X1 port map( A1 => n99, A2 => B(45), ZN => n106);
   U270 : NOR2_X1 port map( A1 => B(44), A2 => n96, ZN => n100);
   U271 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n204);
   U272 : XNOR2_X1 port map( A => n205, B => n155, ZN => n180);
   U273 : NAND2_X1 port map( A1 => n11, A2 => B(41), ZN => n91);
   U274 : NOR2_X1 port map( A1 => n81, A2 => B(40), ZN => n85);
   U275 : CLKBUF_X1 port map( A => n11, Z => n205);
   U276 : NAND2_X1 port map( A1 => B(40), A2 => n81, ZN => n87);
   U277 : INV_X1 port map( A => A(40), ZN => n86);
   U278 : XNOR2_X1 port map( A => n194, B => B(55), ZN => n166);
   U279 : NAND2_X1 port map( A1 => n137, A2 => B(55), ZN => n142);
   U280 : OAI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n69);
   U281 : XNOR2_X1 port map( A => n206, B => n153, ZN => n184);
   U282 : NAND2_X1 port map( A1 => n69, A2 => B(37), ZN => n76);
   U283 : CLKBUF_X1 port map( A => n33, Z => n206);
   U284 : NAND2_X1 port map( A1 => net25602, A2 => net70219, ZN => n150);
   U285 : INV_X1 port map( A => net25644, ZN => net25636);
   U286 : NAND2_X1 port map( A1 => B(35), A2 => n62, ZN => n68);
   U287 : INV_X1 port map( A => net49388, ZN => net25566);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_2_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_2_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_2_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_34_port, carry_33_port, carry_32_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, net47136, net47122, net47106, net47105, 
      net47104, net47103, net47102, net47100, net47098, net47097, net47096, 
      net47095, net47094, net47075, net47068, net47065, net46998, net46993, 
      net46964, net46962, net46941, net46939, net46930, net46905, net47165, 
      net47221, net49454, net49484, net49498, net47125, net46994, net46992, 
      net46991, net47120, net47091, net47084, net47083, net75234, net75475, 
      net75502, net75551, net75553, net51394, net47093, net84237, net84812, 
      net75546, net46911, net46957, net84827, net47139, net47072, net46971, 
      net46969, net46965, net49516, net47228, net47092, net47080, net46986, 
      net75542, net74792, net47146, net46942, net47144, net46970, net46968, 
      net70134, net47134, net47099, net46959, net46958, net46954, net46953, 
      net46952, net46951, net46934, net47148, net46916, net47141, net47124, 
      net47123, net46977, net46974, net75162, net47127, net47126, net46948, 
      net46947, net46946, net46945, net47147, net47129, net47061, net46925, 
      net46924, net46923, net46922, net47232, net47135, net46935, net46931, 
      net46928, net74790, net47158, net46988, net46987, net46983, net46982, 
      net46981, net46980, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129 : std_logic;

begin
   
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1 : INV_X1 port map( A => A(44), ZN => n1);
   U2 : NAND2_X1 port map( A1 => n127, A2 => B(36), ZN => n2);
   U3 : CLKBUF_X1 port map( A => A(51), Z => net75551);
   U4 : BUF_X1 port map( A => n129, Z => n3);
   U5 : NAND2_X1 port map( A1 => n123, A2 => B(42), ZN => n4);
   U6 : NAND2_X1 port map( A1 => n124, A2 => B(38), ZN => n5);
   U7 : INV_X1 port map( A => A(58), ZN => n6);
   U8 : CLKBUF_X1 port map( A => net46970, Z => n7);
   U9 : INV_X1 port map( A => B(61), ZN => net47080);
   U10 : INV_X1 port map( A => B(35), ZN => n101);
   U11 : INV_X1 port map( A => B(36), ZN => n102);
   U12 : INV_X1 port map( A => B(37), ZN => n103);
   U13 : INV_X1 port map( A => B(41), ZN => n105);
   U14 : INV_X1 port map( A => B(57), ZN => net47075);
   U15 : INV_X1 port map( A => B(40), ZN => n104);
   U16 : INV_X1 port map( A => B(44), ZN => n106);
   U17 : INV_X1 port map( A => B(48), ZN => n17);
   U18 : INV_X1 port map( A => B(49), ZN => net47061);
   U19 : INV_X1 port map( A => B(63), ZN => n40);
   U20 : NAND2_X1 port map( A1 => net46998, A2 => n100, ZN => SUM(64));
   U21 : INV_X1 port map( A => B(52), ZN => net47065);
   U22 : INV_X1 port map( A => B(45), ZN => n107);
   U23 : INV_X1 port map( A => B(56), ZN => net47072);
   U24 : INV_X1 port map( A => B(53), ZN => net47068);
   U25 : AND3_X1 port map( A1 => net46935, A2 => n11, A3 => net47065, ZN => n19
                           );
   U26 : NAND2_X1 port map( A1 => net47158, A2 => B(60), ZN => net46987);
   U27 : NAND2_X1 port map( A1 => net46987, A2 => net46988, ZN => net46986);
   U28 : NAND2_X1 port map( A1 => net46988, A2 => net46987, ZN => net47232);
   U29 : OAI21_X1 port map( B1 => net74790, B2 => net46982, A => net46983, ZN 
                           => net47158);
   U30 : OAI21_X1 port map( B1 => net47158, B2 => B(60), A => A(60), ZN => 
                           net46988);
   U31 : INV_X1 port map( A => A(59), ZN => net46982);
   U32 : INV_X1 port map( A => net46982, ZN => net47165);
   U33 : OAI21_X1 port map( B1 => net46981, B2 => net46982, A => net46983, ZN 
                           => net46980);
   U34 : NOR2_X1 port map( A1 => net46974, A2 => B(59), ZN => net74790);
   U35 : XNOR2_X1 port map( A => net46980, B => B(60), ZN => net47093);
   U36 : NOR2_X1 port map( A1 => net46974, A2 => B(59), ZN => net46981);
   U37 : NAND2_X1 port map( A1 => net47123, A2 => B(59), ZN => net46983);
   U38 : XNOR2_X1 port map( A => net47124, B => B(59), ZN => net47094);
   U39 : NAND2_X1 port map( A1 => net47135, A2 => B(51), ZN => net46935);
   U40 : NAND2_X1 port map( A1 => net46935, A2 => n9, ZN => net75502);
   U41 : NAND2_X1 port map( A1 => net46935, A2 => n11, ZN => net46934);
   U42 : OAI21_X1 port map( B1 => net46930, B2 => n10, A => net46931, ZN => 
                           net47135);
   U43 : XNOR2_X1 port map( A => net47135, B => B(51), ZN => net47102);
   U44 : NOR2_X1 port map( A1 => net46922, A2 => B(50), ZN => n10);
   U45 : OAI21_X1 port map( B1 => net46928, B2 => B(51), A => A(51), ZN => n11)
                           ;
   U46 : OAI21_X1 port map( B1 => net46928, B2 => B(51), A => A(51), ZN => n9);
   U47 : OAI21_X1 port map( B1 => n8, B2 => net46930, A => net46931, ZN => 
                           net46928);
   U48 : NOR2_X1 port map( A1 => net46922, A2 => B(50), ZN => n8);
   U49 : XNOR2_X1 port map( A => net47129, B => B(50), ZN => net47103);
   U50 : NAND2_X1 port map( A1 => net47129, A2 => B(50), ZN => net46931);
   U51 : INV_X1 port map( A => A(50), ZN => net46930);
   U52 : NAND2_X1 port map( A1 => net47232, A2 => B(61), ZN => net46994);
   U53 : XNOR2_X1 port map( A => net47232, B => net47080, ZN => net47092);
   U54 : CLKBUF_X1 port map( A => A(60), Z => net51394);
   U55 : OAI21_X1 port map( B1 => net47147, B2 => net46924, A => net46925, ZN 
                           => net47129);
   U56 : INV_X1 port map( A => A(49), ZN => net46924);
   U57 : CLKBUF_X1 port map( A => net46924, Z => net84812);
   U58 : OAI21_X1 port map( B1 => net46923, B2 => net46924, A => net46925, ZN 
                           => net46922);
   U59 : NOR2_X1 port map( A1 => net46916, A2 => B(49), ZN => net47147);
   U60 : XNOR2_X1 port map( A => net46916, B => net47061, ZN => net47104);
   U61 : NAND2_X1 port map( A1 => net47148, A2 => B(49), ZN => net46925);
   U62 : NOR2_X1 port map( A1 => net47148, A2 => B(49), ZN => net46923);
   U63 : NOR2_X1 port map( A1 => net46945, A2 => B(54), ZN => net75162);
   U64 : OAI21_X1 port map( B1 => net75162, B2 => net46953, A => net46954, ZN 
                           => net47134);
   U65 : OAI21_X1 port map( B1 => net46947, B2 => net46946, A => net46948, ZN 
                           => net46945);
   U66 : NOR2_X1 port map( A1 => net46945, A2 => B(54), ZN => net46952);
   U67 : INV_X1 port map( A => A(53), ZN => net46947);
   U68 : XNOR2_X1 port map( A => net47100, B => net46947, ZN => SUM(53));
   U69 : OAI21_X1 port map( B1 => n12, B2 => net46947, A => net46948, ZN => 
                           net47126);
   U70 : OAI21_X1 port map( B1 => n12, B2 => net46947, A => net46948, ZN => 
                           net47127);
   U71 : NOR2_X1 port map( A1 => B(53), A2 => net47146, ZN => net46946);
   U72 : NAND2_X1 port map( A1 => net47126, A2 => B(54), ZN => net46954);
   U73 : XNOR2_X1 port map( A => B(54), B => net47127, ZN => net47099);
   U74 : NAND2_X1 port map( A1 => net47146, A2 => B(53), ZN => net46948);
   U75 : NOR2_X1 port map( A1 => net46939, A2 => B(53), ZN => n12);
   U76 : OAI21_X1 port map( B1 => n6, B2 => n13, A => net46977, ZN => net46974)
                           ;
   U77 : NOR2_X1 port map( A1 => B(58), A2 => net47144, ZN => n13);
   U78 : OAI21_X1 port map( B1 => net47141, B2 => n6, A => net46977, ZN => 
                           net47123);
   U79 : OAI21_X1 port map( B1 => n6, B2 => net47141, A => net46977, ZN => 
                           net47124);
   U80 : NOR2_X1 port map( A1 => B(58), A2 => net46968, ZN => net47141);
   U81 : NAND2_X1 port map( A1 => net46968, A2 => B(58), ZN => net46977);
   U82 : XNOR2_X1 port map( A => net47144, B => B(58), ZN => net47095);
   U83 : CLKBUF_X1 port map( A => A(58), Z => net49498);
   U84 : OAI21_X1 port map( B1 => n18, B2 => n15, A => n16, ZN => net46916);
   U85 : INV_X1 port map( A => A(48), ZN => n15);
   U86 : CLKBUF_X1 port map( A => n15, Z => net84237);
   U87 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => net47148);
   U88 : NOR2_X1 port map( A1 => net75546, A2 => B(48), ZN => n18);
   U89 : XNOR2_X1 port map( A => net75546, B => n17, ZN => net47105);
   U90 : NAND2_X1 port map( A1 => net46911, A2 => B(48), ZN => n16);
   U91 : NOR2_X1 port map( A1 => net46911, A2 => B(48), ZN => n14);
   U92 : OAI21_X1 port map( B1 => net75542, B2 => n19, A => net46942, ZN => 
                           net47146);
   U93 : NAND2_X1 port map( A1 => net46934, A2 => B(52), ZN => net46942);
   U94 : NOR2_X1 port map( A1 => net75502, A2 => B(52), ZN => net74792);
   U95 : NAND2_X1 port map( A1 => net46958, A2 => net46959, ZN => net70134);
   U96 : NAND2_X1 port map( A1 => net70134, A2 => B(56), ZN => net84827);
   U97 : XNOR2_X1 port map( A => net70134, B => net47072, ZN => net47097);
   U98 : NAND2_X1 port map( A1 => net70134, A2 => B(56), ZN => net46965);
   U99 : NAND2_X1 port map( A1 => B(55), A2 => net47134, ZN => net46958);
   U100 : NAND2_X1 port map( A1 => net46958, A2 => net46959, ZN => net46957);
   U101 : OAI21_X1 port map( B1 => net46951, B2 => B(55), A => A(55), ZN => 
                           net46959);
   U102 : OAI21_X1 port map( B1 => net46952, B2 => net46953, A => net46954, ZN 
                           => net46951);
   U103 : INV_X1 port map( A => A(54), ZN => net46953);
   U104 : XNOR2_X1 port map( A => net47134, B => B(55), ZN => net47098);
   U105 : CLKBUF_X1 port map( A => A(55), Z => net75553);
   U106 : XNOR2_X1 port map( A => A(54), B => net47099, ZN => SUM(54));
   U107 : OAI21_X1 port map( B1 => net46969, B2 => net46970, A => net46971, ZN 
                           => net46968);
   U108 : INV_X1 port map( A => A(57), ZN => net46970);
   U109 : XNOR2_X1 port map( A => n7, B => net47096, ZN => SUM(57));
   U110 : OAI21_X1 port map( B1 => net46969, B2 => net46970, A => net46971, ZN 
                           => net47144);
   U111 : INV_X1 port map( A => A(52), ZN => net75542);
   U112 : OAI21_X1 port map( B1 => net74792, B2 => net46941, A => net46942, ZN 
                           => net46939);
   U113 : INV_X1 port map( A => A(52), ZN => net46941);
   U114 : XNOR2_X1 port map( A => net47092, B => net47228, ZN => SUM(61));
   U115 : NOR2_X1 port map( A1 => net46986, A2 => B(61), ZN => net46992);
   U116 : NOR2_X1 port map( A1 => B(61), A2 => net46986, ZN => net49516);
   U117 : INV_X1 port map( A => A(61), ZN => net47228);
   U118 : OAI21_X1 port map( B1 => net49516, B2 => net47228, A => net46994, ZN 
                           => net47125);
   U119 : INV_X1 port map( A => A(61), ZN => net46993);
   U120 : NOR2_X1 port map( A1 => net47139, A2 => B(57), ZN => net46969);
   U121 : OAI21_X1 port map( B1 => n20, B2 => n21, A => net46965, ZN => 
                           net47139);
   U122 : NAND2_X1 port map( A1 => net47139, A2 => B(57), ZN => net46971);
   U123 : INV_X1 port map( A => A(56), ZN => n21);
   U124 : OAI21_X1 port map( B1 => net46964, B2 => n20, A => net84827, ZN => 
                           net46962);
   U125 : NOR2_X1 port map( A1 => net46957, A2 => B(56), ZN => n20);
   U126 : INV_X1 port map( A => A(56), ZN => net46964);
   U127 : NAND2_X1 port map( A1 => n22, A2 => n24, ZN => net75546);
   U128 : OAI21_X1 port map( B1 => net46905, B2 => B(47), A => A(47), ZN => n24
                           );
   U129 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => net46911);
   U130 : OAI21_X1 port map( B1 => net46905, B2 => B(47), A => A(47), ZN => n23
                           );
   U131 : NAND2_X1 port map( A1 => net47136, A2 => B(47), ZN => n22);
   U132 : XNOR2_X1 port map( A => net47136, B => B(47), ZN => net47106);
   U133 : CLKBUF_X1 port map( A => A(47), Z => net75234);
   U134 : OAI21_X1 port map( B1 => n68, B2 => B(39), A => A(39), ZN => n25);
   U135 : CLKBUF_X1 port map( A => n91, Z => n26);
   U136 : INV_X1 port map( A => A(46), ZN => n27);
   U137 : NAND2_X1 port map( A1 => n50, A2 => B(37), ZN => n28);
   U138 : XNOR2_X1 port map( A => net47093, B => net51394, ZN => SUM(60));
   U139 : NAND2_X1 port map( A1 => n25, A2 => n73, ZN => n29);
   U140 : CLKBUF_X1 port map( A => A(34), Z => n30);
   U141 : INV_X1 port map( A => net46930, ZN => net75475);
   U142 : NAND2_X1 port map( A1 => n127, A2 => B(36), ZN => n31);
   U143 : CLKBUF_X1 port map( A => n95, Z => n32);
   U144 : NOR2_X1 port map( A1 => B(42), A2 => n79, ZN => n33);
   U145 : XNOR2_X1 port map( A => n120, B => n59, ZN => SUM(35));
   U146 : INV_X1 port map( A => A(41), ZN => n34);
   U147 : INV_X1 port map( A => A(35), ZN => n59);
   U148 : NOR2_X1 port map( A1 => n93, A2 => B(46), ZN => n35);
   U149 : XNOR2_X1 port map( A => n26, B => n111, ZN => SUM(44));
   U150 : INV_X1 port map( A => A(37), ZN => n66);
   U151 : XNOR2_X1 port map( A => n115, B => n77, ZN => SUM(40));
   U152 : NOR2_X1 port map( A1 => n75, A2 => B(41), ZN => n36);
   U153 : NOR2_X1 port map( A1 => n89, A2 => B(45), ZN => n37);
   U154 : INV_X1 port map( A => A(44), ZN => n91);
   U155 : XNOR2_X1 port map( A => n108, B => net46941, ZN => SUM(52));
   U156 : INV_X1 port map( A => A(45), ZN => n95);
   U157 : NOR2_X1 port map( A1 => n57, A2 => B(36), ZN => n38);
   U158 : XNOR2_X1 port map( A => n119, B => n63, ZN => SUM(36));
   U159 : XNOR2_X1 port map( A => net47105, B => net84237, ZN => SUM(48));
   U160 : INV_X1 port map( A => A(40), ZN => n77);
   U161 : XNOR2_X1 port map( A => n39, B => n41, ZN => SUM(63));
   U162 : XNOR2_X1 port map( A => n42, B => n40, ZN => n41);
   U163 : NAND2_X1 port map( A1 => n40, A2 => net49454, ZN => net47122);
   U164 : OAI21_X1 port map( B1 => net47084, B2 => net47083, A => net47120, ZN 
                           => n42);
   U165 : INV_X1 port map( A => A(62), ZN => net47084);
   U166 : CLKBUF_X1 port map( A => net47084, Z => n43);
   U167 : INV_X1 port map( A => A(63), ZN => n39);
   U168 : CLKBUF_X1 port map( A => n39, Z => net49454);
   U169 : NAND2_X1 port map( A1 => B(63), A2 => net49484, ZN => net46998);
   U170 : NOR2_X1 port map( A1 => net47125, A2 => B(62), ZN => net47083);
   U171 : OAI21_X1 port map( B1 => n43, B2 => net47083, A => net47120, ZN => 
                           net47221);
   U172 : NAND2_X1 port map( A1 => net47125, A2 => B(62), ZN => net47120);
   U173 : XNOR2_X1 port map( A => net47091, B => A(62), ZN => SUM(62));
   U174 : XNOR2_X1 port map( A => net46991, B => B(62), ZN => net47091);
   U175 : NOR2_X1 port map( A1 => B(38), A2 => n64, ZN => n44);
   U176 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => n45);
   U177 : NOR2_X1 port map( A1 => n72, A2 => B(40), ZN => n46);
   U178 : INV_X1 port map( A => A(41), ZN => n81);
   U179 : NOR2_X1 port map( A1 => n45, A2 => B(44), ZN => n47);
   U180 : XNOR2_X1 port map( A => net75502, B => net47065, ZN => n108);
   U181 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n48);
   U182 : XNOR2_X1 port map( A => n114, B => n81, ZN => SUM(41));
   U183 : XNOR2_X1 port map( A => n110, B => n32, ZN => SUM(45));
   U184 : XNOR2_X1 port map( A => n86, B => n106, ZN => n111);
   U185 : NAND2_X1 port map( A1 => n45, A2 => B(44), ZN => n92);
   U186 : XNOR2_X1 port map( A => n29, B => n104, ZN => n115);
   U187 : NAND2_X1 port map( A1 => n72, A2 => B(40), ZN => n78);
   U188 : NOR2_X1 port map( A1 => n61, A2 => B(37), ZN => n49);
   U189 : OAI21_X1 port map( B1 => n38, B2 => n63, A => n2, ZN => n50);
   U190 : INV_X1 port map( A => n98, ZN => n51);
   U191 : INV_X1 port map( A => A(46), ZN => n98);
   U192 : INV_X1 port map( A => A(38), ZN => n70);
   U193 : XNOR2_X1 port map( A => A(38), B => n117, ZN => SUM(38));
   U194 : INV_X1 port map( A => n85, ZN => n52);
   U195 : INV_X1 port map( A => A(42), ZN => n85);
   U196 : NOR2_X1 port map( A1 => n54, A2 => B(35), ZN => n53);
   U197 : INV_X1 port map( A => A(36), ZN => n63);
   U198 : XNOR2_X1 port map( A => net84812, B => net47104, ZN => SUM(49));
   U199 : OAI21_X1 port map( B1 => net46993, B2 => net46992, A => net46994, ZN 
                           => net46991);
   U200 : INV_X1 port map( A => net49454, ZN => net49484);
   U201 : XNOR2_X1 port map( A => net47097, B => net46964, ZN => SUM(56));
   U202 : XNOR2_X1 port map( A => net75475, B => net47103, ZN => SUM(50));
   U203 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => n86);
   U204 : NAND2_X1 port map( A1 => n74, A2 => n73, ZN => n72);
   U205 : XNOR2_X1 port map( A => n48, B => n101, ZN => n120);
   U206 : NAND2_X1 port map( A1 => n54, A2 => B(35), ZN => n60);
   U207 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n93);
   U208 : NAND2_X1 port map( A1 => n122, A2 => B(46), ZN => n99);
   U209 : XNOR2_X1 port map( A => n122, B => B(46), ZN => n109);
   U210 : NOR2_X1 port map( A1 => B(46), A2 => n93, ZN => n97);
   U211 : NOR2_X1 port map( A1 => n89, A2 => B(45), ZN => n94);
   U212 : OAI21_X1 port map( B1 => n37, B2 => n95, A => n96, ZN => n122);
   U213 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => n79);
   U214 : XNOR2_X1 port map( A => n123, B => B(42), ZN => n113);
   U215 : NOR2_X1 port map( A1 => n79, A2 => B(42), ZN => n84);
   U216 : NOR2_X1 port map( A1 => n75, A2 => B(41), ZN => n80);
   U217 : OAI21_X1 port map( B1 => n36, B2 => n34, A => n82, ZN => n123);
   U218 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n28, ZN => n64);
   U219 : NAND2_X1 port map( A1 => n124, A2 => B(38), ZN => n71);
   U220 : XNOR2_X1 port map( A => n124, B => B(38), ZN => n117);
   U221 : NOR2_X1 port map( A1 => n64, A2 => B(38), ZN => n69);
   U222 : NOR2_X1 port map( A1 => n61, A2 => B(37), ZN => n65);
   U223 : OAI21_X1 port map( B1 => n49, B2 => n66, A => n67, ZN => n124);
   U224 : OAI21_X1 port map( B1 => n35, B2 => n98, A => n99, ZN => net46905);
   U225 : OAI21_X1 port map( B1 => n97, B2 => n27, A => n99, ZN => net47136);
   U226 : OAI21_X1 port map( B1 => n85, B2 => n33, A => n4, ZN => n83);
   U227 : NAND2_X1 port map( A1 => n125, A2 => B(43), ZN => n87);
   U228 : OAI21_X1 port map( B1 => n125, B2 => B(43), A => A(43), ZN => n88);
   U229 : XNOR2_X1 port map( A => B(43), B => n83, ZN => n112);
   U230 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n4, ZN => n125);
   U231 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n68);
   U232 : NAND2_X1 port map( A1 => n126, A2 => B(39), ZN => n73);
   U233 : OAI21_X1 port map( B1 => n68, B2 => B(39), A => A(39), ZN => n74);
   U234 : XNOR2_X1 port map( A => n126, B => B(39), ZN => n116);
   U235 : OAI21_X1 port map( B1 => n44, B2 => n70, A => n5, ZN => n126);
   U236 : XNOR2_X1 port map( A => net46962, B => net47075, ZN => net47096);
   U237 : OAI21_X1 port map( B1 => n58, B2 => n59, A => n60, ZN => n57);
   U238 : XNOR2_X1 port map( A => n127, B => n102, ZN => n119);
   U239 : NOR2_X1 port map( A1 => n57, A2 => B(36), ZN => n62);
   U240 : NOR2_X1 port map( A1 => n48, A2 => B(35), ZN => n58);
   U241 : OAI21_X1 port map( B1 => n53, B2 => n59, A => n60, ZN => n127);
   U242 : XNOR2_X1 port map( A => net46939, B => net47068, ZN => net47100);
   U243 : XNOR2_X1 port map( A => net47095, B => net49498, ZN => SUM(58));
   U244 : OAI21_X1 port map( B1 => n90, B2 => n91, A => n92, ZN => n89);
   U245 : XNOR2_X1 port map( A => n128, B => n107, ZN => n110);
   U246 : NAND2_X1 port map( A1 => n128, A2 => B(45), ZN => n96);
   U247 : NOR2_X1 port map( A1 => n86, A2 => B(44), ZN => n90);
   U248 : OAI21_X1 port map( B1 => n47, B2 => n1, A => n92, ZN => n128);
   U249 : OAI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n75);
   U250 : XNOR2_X1 port map( A => n3, B => n105, ZN => n114);
   U251 : NAND2_X1 port map( A1 => n129, A2 => B(41), ZN => n82);
   U252 : NOR2_X1 port map( A1 => n29, A2 => B(40), ZN => n76);
   U253 : OAI21_X1 port map( B1 => n46, B2 => n77, A => n78, ZN => n129);
   U254 : OAI21_X1 port map( B1 => n62, B2 => n63, A => n31, ZN => n61);
   U255 : XNOR2_X1 port map( A => n50, B => n103, ZN => n118);
   U256 : NAND2_X1 port map( A1 => n50, A2 => B(37), ZN => n67);
   U257 : NAND2_X1 port map( A1 => B(34), A2 => A(34), ZN => n55);
   U258 : OAI21_X1 port map( B1 => A(34), B2 => B(34), A => carry_34_port, ZN 
                           => n56);
   U259 : XNOR2_X1 port map( A => n121, B => n30, ZN => SUM(34));
   U260 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n54);
   U261 : XNOR2_X1 port map( A => carry_34_port, B => B(34), ZN => n121);
   U262 : XNOR2_X1 port map( A => net47106, B => net75234, ZN => SUM(47));
   U263 : NAND2_X1 port map( A1 => net47122, A2 => net47221, ZN => n100);
   U264 : XNOR2_X1 port map( A => A(43), B => n112, ZN => SUM(43));
   U265 : XNOR2_X1 port map( A => net47102, B => net75551, ZN => SUM(51));
   U266 : XNOR2_X1 port map( A => n118, B => n66, ZN => SUM(37));
   U267 : XNOR2_X1 port map( A => net47098, B => net75553, ZN => SUM(55));
   U268 : XNOR2_X1 port map( A => A(39), B => n116, ZN => SUM(39));
   U269 : XNOR2_X1 port map( A => net47094, B => net47165, ZN => SUM(59));
   U270 : XNOR2_X1 port map( A => n51, B => n109, ZN => SUM(46));
   U271 : XNOR2_X1 port map( A => n52, B => n113, ZN => SUM(42));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_3_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_3_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_3_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_33_port, carry_32_port, carry_31_port, carry_30_port, 
      carry_29_port, carry_28_port, carry_27_port, carry_26_port, carry_25_port
      , carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, net49365, net49360, net49352, net49347, net49331, net49330,
      net49314, net49309, net49306, net49202, net49201, net49200, net49184, 
      net49183, net49147, net49130, net49500, net49512, net49373, net49316, 
      net61101, net49310, carry_63_port, net49363, net49321, net49301, net49196
      , net49194, net75320, net49397, net49366, net49320, net49195, net49193, 
      net74903, net49322, net49298, net49182, net84553, net75559, net49284, 
      net49136, net49369, net49329, net49287, net49150, net49149, net49148, 
      net49141, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184 : 
      std_logic;

begin
   
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_63 : FA_X1 port map( A => carry_63_port, B => B(63), CI => A(63), CO => 
                           SUM(64), S => SUM(63));
   U1 : CLKBUF_X1 port map( A => n72, Z => n1);
   U2 : INV_X1 port map( A => A(37), ZN => n2);
   U3 : INV_X1 port map( A => A(53), ZN => n3);
   U4 : CLKBUF_X1 port map( A => net49149, Z => n4);
   U5 : BUF_X1 port map( A => A(46), Z => net61101);
   U6 : INV_X1 port map( A => A(44), ZN => n5);
   U7 : INV_X1 port map( A => A(44), ZN => n105);
   U8 : INV_X1 port map( A => B(35), ZN => n138);
   U9 : INV_X1 port map( A => B(36), ZN => n139);
   U10 : INV_X1 port map( A => A(36), ZN => n76);
   U11 : INV_X1 port map( A => B(40), ZN => n141);
   U12 : INV_X1 port map( A => B(52), ZN => n145);
   U13 : INV_X1 port map( A => B(56), ZN => net49301);
   U14 : INV_X1 port map( A => B(34), ZN => n137);
   U15 : INV_X1 port map( A => B(39), ZN => n140);
   U16 : INV_X1 port map( A => B(43), ZN => n142);
   U17 : INV_X1 port map( A => B(44), ZN => n143);
   U18 : INV_X1 port map( A => B(47), ZN => net49284);
   U19 : INV_X1 port map( A => B(60), ZN => net49306);
   U20 : INV_X1 port map( A => B(51), ZN => n144);
   U21 : INV_X1 port map( A => B(48), ZN => net49287);
   U22 : INV_X1 port map( A => B(55), ZN => net49298);
   U23 : XNOR2_X1 port map( A => net49329, B => n4, ZN => SUM(48));
   U24 : INV_X1 port map( A => A(48), ZN => net49149);
   U25 : OAI21_X1 port map( B1 => net49369, B2 => net49149, A => net49150, ZN 
                           => net49352);
   U26 : OAI21_X1 port map( B1 => net49148, B2 => net49149, A => net49150, ZN 
                           => net49147);
   U27 : XNOR2_X1 port map( A => n9, B => net49287, ZN => net49329);
   U28 : OAI21_X1 port map( B1 => n7, B2 => n10, A => n8, ZN => n9);
   U29 : NOR2_X1 port map( A1 => n9, A2 => B(48), ZN => net49369);
   U30 : INV_X1 port map( A => A(47), ZN => n7);
   U31 : CLKBUF_X1 port map( A => n7, Z => net84553);
   U32 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n8, ZN => net49141);
   U33 : NOR2_X1 port map( A1 => net49136, A2 => B(47), ZN => n10);
   U34 : NAND2_X1 port map( A1 => net49141, A2 => B(48), ZN => net49150);
   U35 : NOR2_X1 port map( A1 => net49141, A2 => B(48), ZN => net49148);
   U36 : NOR2_X1 port map( A1 => B(47), A2 => net49136, ZN => n6);
   U37 : NAND2_X1 port map( A1 => B(47), A2 => net75559, ZN => n8);
   U38 : NAND2_X1 port map( A1 => n13, A2 => n11, ZN => net49136);
   U39 : OAI21_X1 port map( B1 => net49360, B2 => B(46), A => A(46), ZN => n13)
                           ;
   U40 : XNOR2_X1 port map( A => net75559, B => net49284, ZN => net49330);
   U41 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => net75559);
   U42 : XNOR2_X1 port map( A => net49360, B => B(46), ZN => net49331);
   U43 : OAI21_X1 port map( B1 => net49130, B2 => B(46), A => A(46), ZN => n12)
                           ;
   U44 : NAND2_X1 port map( A1 => net49130, A2 => B(46), ZN => n11);
   U45 : CLKBUF_X1 port map( A => n90, Z => n14);
   U46 : BUF_X1 port map( A => A(42), Z => n43);
   U47 : NOR2_X1 port map( A1 => net49500, A2 => B(60), ZN => n15);
   U48 : NOR2_X1 port map( A1 => n114, A2 => B(51), ZN => n16);
   U49 : CLKBUF_X1 port map( A => n101, Z => n17);
   U50 : OAI21_X1 port map( B1 => n19, B2 => n22, A => n20, ZN => n18);
   U51 : NOR2_X1 port map( A1 => n18, A2 => B(56), ZN => net49194);
   U52 : INV_X1 port map( A => A(55), ZN => n19);
   U53 : XNOR2_X1 port map( A => net49322, B => n19, ZN => SUM(55));
   U54 : NOR2_X1 port map( A1 => net49182, A2 => B(55), ZN => n22);
   U55 : NAND2_X1 port map( A1 => B(55), A2 => net74903, ZN => n20);
   U56 : OAI21_X1 port map( B1 => n21, B2 => n22, A => n20, ZN => net49363);
   U57 : INV_X1 port map( A => A(55), ZN => n21);
   U58 : NAND2_X1 port map( A1 => net49184, A2 => net49183, ZN => net49182);
   U59 : XNOR2_X1 port map( A => net74903, B => net49298, ZN => net49322);
   U60 : NAND2_X1 port map( A1 => net49184, A2 => net49183, ZN => net74903);
   U61 : XNOR2_X1 port map( A => net49320, B => net49397, ZN => SUM(57));
   U62 : INV_X1 port map( A => net75320, ZN => net49397);
   U63 : INV_X1 port map( A => A(57), ZN => net75320);
   U64 : OAI21_X1 port map( B1 => net49201, B2 => net49365, A => net49202, ZN 
                           => net49347);
   U65 : XNOR2_X1 port map( A => net49366, B => B(57), ZN => net49320);
   U66 : INV_X1 port map( A => A(57), ZN => net49201);
   U67 : OAI21_X1 port map( B1 => net49194, B2 => net49195, A => net49196, ZN 
                           => net49366);
   U68 : NOR2_X1 port map( A1 => B(57), A2 => net49193, ZN => net49200);
   U69 : INV_X1 port map( A => A(56), ZN => net49195);
   U70 : XNOR2_X1 port map( A => net49321, B => net49195, ZN => SUM(56));
   U71 : OAI21_X1 port map( B1 => net49194, B2 => net49195, A => net49196, ZN 
                           => net49193);
   U72 : NAND2_X1 port map( A1 => net49366, A2 => B(57), ZN => net49202);
   U73 : NOR2_X1 port map( A1 => net49193, A2 => B(57), ZN => net49365);
   U74 : NAND2_X1 port map( A1 => net49363, A2 => B(56), ZN => net49196);
   U75 : XNOR2_X1 port map( A => net49363, B => net49301, ZN => net49321);
   U76 : INV_X1 port map( A => A(52), ZN => n23);
   U77 : OAI21_X1 port map( B1 => n110, B2 => B(50), A => A(50), ZN => n24);
   U78 : NAND2_X1 port map( A1 => n115, A2 => n24, ZN => n25);
   U79 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n26);
   U80 : CLKBUF_X1 port map( A => A(33), Z => n27);
   U81 : CLKBUF_X1 port map( A => A(49), Z => n28);
   U82 : CLKBUF_X1 port map( A => A(50), Z => n29);
   U83 : NOR2_X1 port map( A1 => net49147, A2 => B(49), ZN => n30);
   U84 : NOR2_X1 port map( A1 => n70, A2 => B(36), ZN => n31);
   U85 : INV_X1 port map( A => A(40), ZN => n90);
   U86 : CLKBUF_X1 port map( A => A(59), Z => n62);
   U87 : CLKBUF_X1 port map( A => A(38), Z => n32);
   U88 : NOR2_X1 port map( A1 => B(41), A2 => n51, ZN => n33);
   U89 : INV_X1 port map( A => n94, ZN => n34);
   U90 : NOR2_X1 port map( A1 => net49500, A2 => B(60), ZN => n35);
   U91 : INV_X1 port map( A => n80, ZN => n36);
   U92 : INV_X1 port map( A => A(35), ZN => n72);
   U93 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => n37);
   U94 : OAI21_X1 port map( B1 => n78, B2 => B(38), A => A(38), ZN => n38);
   U95 : INV_X1 port map( A => A(34), ZN => n68);
   U96 : XNOR2_X1 port map( A => net84553, B => net49330, ZN => SUM(47));
   U97 : INV_X1 port map( A => n108, ZN => n39);
   U98 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => n40);
   U99 : NOR2_X1 port map( A1 => B(37), A2 => n74, ZN => n41);
   U100 : INV_X1 port map( A => A(43), ZN => n101);
   U101 : NOR2_X1 port map( A1 => B(53), A2 => n121, ZN => n42);
   U102 : XNOR2_X1 port map( A => n166, B => n68, ZN => SUM(34));
   U103 : XNOR2_X1 port map( A => n87, B => n161, ZN => SUM(39));
   U104 : XNOR2_X1 port map( A => n165, B => n1, ZN => SUM(35));
   U105 : INV_X1 port map( A => A(39), ZN => n87);
   U106 : XNOR2_X1 port map( A => n157, B => n17, ZN => SUM(43));
   U107 : NOR2_X1 port map( A1 => B(58), A2 => n129, ZN => n44);
   U108 : OAI21_X1 port map( B1 => n45, B2 => n46, A => n47, ZN => 
                           carry_63_port);
   U109 : NAND2_X1 port map( A1 => B(62), A2 => n50, ZN => n47);
   U110 : NOR2_X1 port map( A1 => B(62), A2 => n50, ZN => n46);
   U111 : INV_X1 port map( A => A(62), ZN => n45);
   U112 : XNOR2_X1 port map( A => n48, B => B(62), ZN => n49);
   U113 : OAI21_X1 port map( B1 => net49309, B2 => net49310, A => net49314, ZN 
                           => n50);
   U114 : INV_X1 port map( A => A(61), ZN => net49310);
   U115 : OAI21_X1 port map( B1 => net49310, B2 => net49309, A => net49314, ZN 
                           => n48);
   U116 : XNOR2_X1 port map( A => n49, B => A(62), ZN => SUM(62));
   U117 : BUF_X1 port map( A => A(61), Z => net49512);
   U118 : OAI21_X1 port map( B1 => n90, B2 => n89, A => n91, ZN => n51);
   U119 : INV_X1 port map( A => n127, ZN => n52);
   U120 : NOR2_X1 port map( A1 => n96, A2 => B(43), ZN => n53);
   U121 : NOR2_X1 port map( A1 => n40, A2 => B(39), ZN => n54);
   U122 : NOR2_X1 port map( A1 => B(34), A2 => n63, ZN => n55);
   U123 : NOR2_X1 port map( A1 => n66, A2 => B(35), ZN => n56);
   U124 : XNOR2_X1 port map( A => n164, B => n76, ZN => SUM(36));
   U125 : XNOR2_X1 port map( A => n26, B => n142, ZN => n157);
   U126 : NAND2_X1 port map( A1 => n115, A2 => n116, ZN => n114);
   U127 : XNOR2_X1 port map( A => n160, B => n14, ZN => SUM(40));
   U128 : XNOR2_X1 port map( A => n156, B => n105, ZN => SUM(44));
   U129 : XNOR2_X1 port map( A => n163, B => n36, ZN => SUM(37));
   U130 : OAI21_X1 port map( B1 => n110, B2 => B(50), A => A(50), ZN => n116);
   U131 : CLKBUF_X1 port map( A => A(54), Z => n57);
   U132 : INV_X1 port map( A => n132, ZN => n58);
   U133 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => n96);
   U134 : XNOR2_X1 port map( A => n40, B => n140, ZN => n161);
   U135 : NAND2_X1 port map( A1 => B(39), A2 => n82, ZN => n88);
   U136 : NAND2_X1 port map( A1 => B(43), A2 => n26, ZN => n102);
   U137 : NAND2_X1 port map( A1 => n38, A2 => n83, ZN => n82);
   U138 : OAI21_X1 port map( B1 => n61, B2 => n35, A => n60, ZN => n59);
   U139 : XNOR2_X1 port map( A => n59, B => B(61), ZN => net49316);
   U140 : INV_X1 port map( A => A(60), ZN => n61);
   U141 : OAI21_X1 port map( B1 => n61, B2 => n15, A => n60, ZN => net49373);
   U142 : NAND2_X1 port map( A1 => net49500, A2 => B(60), ZN => n60);
   U143 : XNOR2_X1 port map( A => net49316, B => net49512, ZN => SUM(61));
   U144 : NAND2_X1 port map( A1 => B(61), A2 => net49373, ZN => net49314);
   U145 : NOR2_X1 port map( A1 => net49373, A2 => B(61), ZN => net49309);
   U146 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => net49500);
   U147 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => n134);
   U148 : OAI21_X1 port map( B1 => n125, B2 => B(54), A => A(54), ZN => 
                           net49184);
   U149 : OAI21_X1 port map( B1 => n173, B2 => B(59), A => A(59), ZN => n136);
   U150 : INV_X1 port map( A => A(51), ZN => n119);
   U151 : XNOR2_X1 port map( A => n151, B => n123, ZN => SUM(52));
   U152 : OAI21_X1 port map( B1 => net49200, B2 => net75320, A => net49202, ZN 
                           => n129);
   U153 : OAI21_X1 port map( B1 => net49365, B2 => net49201, A => net49202, ZN 
                           => n168);
   U154 : NOR2_X1 port map( A1 => n117, A2 => B(52), ZN => n122);
   U155 : OAI21_X1 port map( B1 => n123, B2 => n122, A => n124, ZN => n121);
   U156 : OAI21_X1 port map( B1 => n179, B2 => n23, A => n124, ZN => n169);
   U157 : NOR2_X1 port map( A1 => n182, A2 => B(44), ZN => n104);
   U158 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n103);
   U159 : OAI21_X1 port map( B1 => n181, B2 => n5, A => n106, ZN => n170);
   U160 : NAND2_X1 port map( A1 => n171, A2 => B(41), ZN => n95);
   U161 : XNOR2_X1 port map( A => n51, B => B(41), ZN => n159);
   U162 : NOR2_X1 port map( A1 => n171, A2 => B(41), ZN => n93);
   U163 : NOR2_X1 port map( A1 => n85, A2 => B(40), ZN => n89);
   U164 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n171);
   U165 : OAI21_X1 port map( B1 => n31, B2 => n76, A => n77, ZN => n74);
   U166 : NAND2_X1 port map( A1 => n172, A2 => B(37), ZN => n81);
   U167 : XNOR2_X1 port map( A => n172, B => B(37), ZN => n163);
   U168 : NOR2_X1 port map( A1 => n74, A2 => B(37), ZN => n79);
   U169 : NOR2_X1 port map( A1 => n70, A2 => B(36), ZN => n75);
   U170 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => n172);
   U171 : NOR2_X1 port map( A1 => B(58), A2 => n129, ZN => n131);
   U172 : OAI21_X1 port map( B1 => n132, B2 => n131, A => n133, ZN => n130);
   U173 : OAI21_X1 port map( B1 => n44, B2 => n132, A => n133, ZN => n173);
   U174 : NOR2_X1 port map( A1 => n121, A2 => B(53), ZN => n126);
   U175 : OAI21_X1 port map( B1 => n126, B2 => n3, A => n128, ZN => n125);
   U176 : OAI21_X1 port map( B1 => n42, B2 => n127, A => n128, ZN => n174);
   U177 : NOR2_X1 port map( A1 => net49147, A2 => B(49), ZN => n111);
   U178 : OAI21_X1 port map( B1 => n30, B2 => n112, A => n113, ZN => n110);
   U179 : OAI21_X1 port map( B1 => n112, B2 => n111, A => n113, ZN => n175);
   U180 : NOR2_X1 port map( A1 => n103, A2 => B(45), ZN => n107);
   U181 : OAI21_X1 port map( B1 => n108, B2 => n107, A => n109, ZN => net49130)
                           ;
   U182 : OAI21_X1 port map( B1 => n108, B2 => n107, A => n109, ZN => net49360)
                           ;
   U183 : OAI21_X1 port map( B1 => n94, B2 => n33, A => n95, ZN => n92);
   U184 : NAND2_X1 port map( A1 => n176, A2 => B(42), ZN => n97);
   U185 : OAI21_X1 port map( B1 => n176, B2 => B(42), A => A(42), ZN => n98);
   U186 : XNOR2_X1 port map( A => B(42), B => n92, ZN => n158);
   U187 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n176);
   U188 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U189 : NAND2_X1 port map( A1 => n177, A2 => B(38), ZN => n83);
   U190 : OAI21_X1 port map( B1 => n78, B2 => B(38), A => A(38), ZN => n84);
   U191 : XNOR2_X1 port map( A => n177, B => B(38), ZN => n162);
   U192 : OAI21_X1 port map( B1 => n41, B2 => n2, A => n81, ZN => n177);
   U193 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => n66);
   U194 : XNOR2_X1 port map( A => n178, B => n138, ZN => n165);
   U195 : NAND2_X1 port map( A1 => n178, A2 => B(35), ZN => n73);
   U196 : NOR2_X1 port map( A1 => B(35), A2 => n66, ZN => n71);
   U197 : NOR2_X1 port map( A1 => n37, A2 => B(34), ZN => n67);
   U198 : OAI21_X1 port map( B1 => n55, B2 => n68, A => n69, ZN => n178);
   U199 : NOR2_X1 port map( A1 => n180, A2 => B(52), ZN => n179);
   U200 : NOR2_X1 port map( A1 => n114, A2 => B(51), ZN => n118);
   U201 : OAI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n117);
   U202 : OAI21_X1 port map( B1 => n16, B2 => n119, A => n120, ZN => n180);
   U203 : NAND2_X1 port map( A1 => n180, A2 => B(52), ZN => n124);
   U204 : NOR2_X1 port map( A1 => n99, A2 => B(44), ZN => n181);
   U205 : OAI21_X1 port map( B1 => n101, B2 => n100, A => n102, ZN => n99);
   U206 : XNOR2_X1 port map( A => n182, B => n143, ZN => n156);
   U207 : NAND2_X1 port map( A1 => n99, A2 => B(44), ZN => n106);
   U208 : NOR2_X1 port map( A1 => B(43), A2 => n96, ZN => n100);
   U209 : OAI21_X1 port map( B1 => n101, B2 => n53, A => n102, ZN => n182);
   U210 : NAND2_X1 port map( A1 => B(58), A2 => net49347, ZN => n133);
   U211 : XNOR2_X1 port map( A => n130, B => B(59), ZN => n147);
   U212 : NAND2_X1 port map( A1 => n173, A2 => B(59), ZN => n135);
   U213 : XNOR2_X1 port map( A => n168, B => B(58), ZN => n148);
   U214 : NAND2_X1 port map( A1 => n169, A2 => B(53), ZN => n128);
   U215 : XNOR2_X1 port map( A => n174, B => B(54), ZN => n149);
   U216 : NAND2_X1 port map( A1 => n125, A2 => B(54), ZN => net49183);
   U217 : XNOR2_X1 port map( A => n117, B => n145, ZN => n151);
   U218 : XNOR2_X1 port map( A => n169, B => B(53), ZN => n150);
   U219 : XNOR2_X1 port map( A => net49352, B => B(49), ZN => n154);
   U220 : XNOR2_X1 port map( A => n175, B => B(50), ZN => n153);
   U221 : NAND2_X1 port map( A1 => n175, A2 => B(50), ZN => n115);
   U222 : NAND2_X1 port map( A1 => B(45), A2 => n170, ZN => n109);
   U223 : INV_X1 port map( A => A(45), ZN => n108);
   U224 : XNOR2_X1 port map( A => n147, B => n62, ZN => SUM(59));
   U225 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n85);
   U226 : XNOR2_X1 port map( A => n183, B => n141, ZN => n160);
   U227 : NAND2_X1 port map( A1 => n183, A2 => B(40), ZN => n91);
   U228 : NOR2_X1 port map( A1 => B(39), A2 => n82, ZN => n86);
   U229 : OAI21_X1 port map( B1 => n87, B2 => n54, A => n88, ZN => n183);
   U230 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n70);
   U231 : XNOR2_X1 port map( A => n184, B => n139, ZN => n164);
   U232 : NAND2_X1 port map( A1 => n184, A2 => B(36), ZN => n77);
   U233 : XNOR2_X1 port map( A => carry_33_port, B => B(33), ZN => n167);
   U234 : OAI21_X1 port map( B1 => A(33), B2 => B(33), A => carry_33_port, ZN 
                           => n65);
   U235 : OAI21_X1 port map( B1 => n72, B2 => n56, A => n73, ZN => n184);
   U236 : NAND2_X1 port map( A1 => n25, A2 => B(51), ZN => n120);
   U237 : NAND2_X1 port map( A1 => B(33), A2 => A(33), ZN => n64);
   U238 : XNOR2_X1 port map( A => n167, B => n27, ZN => SUM(33));
   U239 : XNOR2_X1 port map( A => n43, B => n158, ZN => SUM(42));
   U240 : XNOR2_X1 port map( A => n149, B => n57, ZN => SUM(54));
   U241 : XNOR2_X1 port map( A => n170, B => B(45), ZN => n155);
   U242 : XNOR2_X1 port map( A => n153, B => n29, ZN => SUM(50));
   U243 : INV_X1 port map( A => A(58), ZN => n132);
   U244 : XNOR2_X1 port map( A => n150, B => n52, ZN => SUM(53));
   U245 : XNOR2_X1 port map( A => net49331, B => net61101, ZN => SUM(46));
   U246 : XNOR2_X1 port map( A => n134, B => net49306, ZN => n146);
   U247 : XNOR2_X1 port map( A => n146, B => n61, ZN => SUM(60));
   U248 : XNOR2_X1 port map( A => n162, B => n32, ZN => SUM(38));
   U249 : INV_X1 port map( A => A(41), ZN => n94);
   U250 : XNOR2_X1 port map( A => n148, B => n58, ZN => SUM(58));
   U251 : NAND2_X1 port map( A1 => net49352, A2 => B(49), ZN => n113);
   U252 : INV_X1 port map( A => A(49), ZN => n112);
   U253 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => n63);
   U254 : INV_X1 port map( A => A(53), ZN => n127);
   U255 : XNOR2_X1 port map( A => n159, B => n34, ZN => SUM(41));
   U256 : XNOR2_X1 port map( A => n37, B => n137, ZN => n166);
   U257 : NAND2_X1 port map( A1 => B(34), A2 => n63, ZN => n69);
   U258 : XNOR2_X1 port map( A => n155, B => n39, ZN => SUM(45));
   U259 : INV_X1 port map( A => A(52), ZN => n123);
   U260 : XNOR2_X1 port map( A => n154, B => n28, ZN => SUM(49));
   U261 : XNOR2_X1 port map( A => n25, B => n144, ZN => n152);
   U262 : XNOR2_X1 port map( A => n119, B => n152, ZN => SUM(51));
   U263 : INV_X1 port map( A => A(37), ZN => n80);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_4_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_4_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_4_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_30_port, carry_29_port, carry_28_port, carry_27_port, 
      carry_26_port, carry_25_port, carry_24_port, carry_23_port, carry_22_port
      , carry_21_port, carry_20_port, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_15_port, carry_14_port, carry_13_port
      , carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port
      , carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, net60892, net60885, net60871, net60859, 
      net60847, net60848, net60830, net60829, net60828, net60827, net60826, 
      net60825, net60817, net60812, net60811, net60806, net60777, net60702, 
      net60698, net60658, net60657, net60652, net60615, net61029, net61044, 
      carry_63_port, carry_62_port, carry_61_port, carry_60_port, net75572, 
      net74645, net60903, net60705, net60704, net60849, net60816, net60696, 
      net84712, net84833, net75501, net60781, net60635, net60634, net60908, 
      net60856, net60824, net60650, net60633, net84440, net60870, net60641, 
      net60640, net60638, net74646, net60852, net60784, net60653, net60647, 
      net60646, net60645, net60644, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178 : std_logic;

begin
   
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1 : CLKBUF_X1 port map( A => n89, Z => n1);
   U2 : INV_X1 port map( A => A(46), ZN => n2);
   U3 : INV_X1 port map( A => A(38), ZN => n3);
   U4 : CLKBUF_X1 port map( A => n118, Z => n26);
   U5 : INV_X1 port map( A => A(41), ZN => n4);
   U6 : INV_X1 port map( A => A(45), ZN => n5);
   U7 : XOR2_X1 port map( A => A(24), B => B(24), Z => n6);
   U8 : XOR2_X1 port map( A => carry_24_port, B => n6, Z => SUM(24));
   U9 : NAND2_X1 port map( A1 => carry_24_port, A2 => A(24), ZN => n7);
   U10 : NAND2_X1 port map( A1 => carry_24_port, A2 => B(24), ZN => n8);
   U11 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n9);
   U12 : NAND3_X1 port map( A1 => n7, A2 => n8, A3 => n9, ZN => carry_25_port);
   U13 : CLKBUF_X1 port map( A => A(30), Z => n10);
   U14 : NOR2_X1 port map( A1 => net60644, A2 => B(46), ZN => n11);
   U15 : AND2_X1 port map( A1 => n82, A2 => n46, ZN => n84);
   U16 : INV_X1 port map( A => B(52), ZN => n138);
   U17 : INV_X1 port map( A => B(33), ZN => n132);
   U18 : INV_X1 port map( A => B(40), ZN => n135);
   U19 : INV_X1 port map( A => B(41), ZN => net60777);
   U20 : INV_X1 port map( A => B(57), ZN => n140);
   U21 : INV_X1 port map( A => B(31), ZN => n130);
   U22 : INV_X1 port map( A => B(32), ZN => n131);
   U23 : INV_X1 port map( A => B(37), ZN => n134);
   U24 : INV_X1 port map( A => B(48), ZN => n136);
   U25 : INV_X1 port map( A => B(49), ZN => n137);
   U26 : INV_X1 port map( A => B(53), ZN => n139);
   U27 : INV_X1 port map( A => B(36), ZN => n133);
   U28 : INV_X1 port map( A => B(45), ZN => net60784);
   U29 : INV_X1 port map( A => B(44), ZN => net60781);
   U30 : NAND2_X1 port map( A1 => net60852, A2 => B(46), ZN => net60653);
   U31 : OAI21_X1 port map( B1 => n2, B2 => n11, A => net60653, ZN => net60856)
                           ;
   U32 : OAI21_X1 port map( B1 => n11, B2 => net60652, A => net60653, ZN => 
                           net60650);
   U33 : OAI21_X1 port map( B1 => net74646, B2 => n5, A => net60647, ZN => 
                           net60852);
   U34 : XNOR2_X1 port map( A => net60852, B => B(46), ZN => net60825);
   U35 : INV_X1 port map( A => A(45), ZN => net60646);
   U36 : CLKBUF_X1 port map( A => net60646, Z => net84833);
   U37 : OAI21_X1 port map( B1 => net60645, B2 => net60646, A => net60647, ZN 
                           => net60644);
   U38 : NOR2_X1 port map( A1 => net60638, A2 => B(45), ZN => net74646);
   U39 : XNOR2_X1 port map( A => net60870, B => net60784, ZN => net60826);
   U40 : NAND2_X1 port map( A1 => net60638, A2 => B(45), ZN => net60647);
   U41 : NOR2_X1 port map( A1 => net60870, A2 => B(45), ZN => net60645);
   U42 : OAI21_X1 port map( B1 => net84440, B2 => net60640, A => net60641, ZN 
                           => net60870);
   U43 : INV_X1 port map( A => A(44), ZN => net60640);
   U44 : CLKBUF_X1 port map( A => net60640, Z => net84712);
   U45 : OAI21_X1 port map( B1 => net84440, B2 => net60640, A => net60641, ZN 
                           => net60638);
   U46 : NOR2_X1 port map( A1 => net60633, A2 => B(44), ZN => net84440);
   U47 : NAND2_X1 port map( A1 => net75501, A2 => B(44), ZN => net60641);
   U48 : NAND2_X1 port map( A1 => net60634, A2 => net60635, ZN => net60633);
   U49 : NAND2_X1 port map( A1 => net60635, A2 => net60634, ZN => net75501);
   U50 : XNOR2_X1 port map( A => net60824, B => net60908, ZN => SUM(47));
   U51 : CLKBUF_X1 port map( A => A(47), Z => net60908);
   U52 : XNOR2_X1 port map( A => net60856, B => B(47), ZN => net60824);
   U53 : OAI21_X1 port map( B1 => B(47), B2 => net60650, A => A(47), ZN => 
                           net75572);
   U54 : OAI21_X1 port map( B1 => net60650, B2 => B(47), A => A(47), ZN => 
                           net60658);
   U55 : NAND2_X1 port map( A1 => net60856, A2 => B(47), ZN => net60657);
   U56 : INV_X1 port map( A => A(46), ZN => net60652);
   U57 : OAI21_X1 port map( B1 => n21, B2 => B(43), A => A(43), ZN => net60635)
                           ;
   U58 : OAI21_X1 port map( B1 => n17, B2 => n18, A => n19, ZN => n21);
   U59 : INV_X1 port map( A => A(42), ZN => n18);
   U60 : OAI21_X1 port map( B1 => n18, B2 => n17, A => n19, ZN => n16);
   U61 : XNOR2_X1 port map( A => n16, B => B(43), ZN => net60828);
   U62 : NAND2_X1 port map( A1 => n16, A2 => B(43), ZN => net60634);
   U63 : CLKBUF_X1 port map( A => A(43), Z => net60892);
   U64 : NOR2_X1 port map( A1 => n12, A2 => B(42), ZN => n17);
   U65 : OAI21_X1 port map( B1 => n22, B2 => n14, A => n15, ZN => n12);
   U66 : INV_X1 port map( A => A(41), ZN => n14);
   U67 : XNOR2_X1 port map( A => net60830, B => n14, ZN => SUM(41));
   U68 : OAI21_X1 port map( B1 => n13, B2 => n4, A => n15, ZN => n20);
   U69 : NOR2_X1 port map( A1 => net60615, A2 => B(41), ZN => n22);
   U70 : NAND2_X1 port map( A1 => n20, A2 => B(42), ZN => n19);
   U71 : XNOR2_X1 port map( A => n20, B => B(42), ZN => net60829);
   U72 : NOR2_X1 port map( A1 => B(41), A2 => net60615, ZN => n13);
   U73 : NAND2_X1 port map( A1 => net60871, A2 => B(41), ZN => n15);
   U74 : XNOR2_X1 port map( A => net75501, B => net60781, ZN => net60827);
   U75 : NOR2_X1 port map( A1 => net60696, A2 => B(55), ZN => n23);
   U76 : CLKBUF_X1 port map( A => n99, Z => n24);
   U77 : CLKBUF_X1 port map( A => A(51), Z => n176);
   U78 : OAI21_X1 port map( B1 => n91, B2 => B(39), A => A(39), ZN => n25);
   U79 : CLKBUF_X1 port map( A => n108, Z => n44);
   U80 : INV_X1 port map( A => A(31), ZN => n66);
   U81 : OAI21_X1 port map( B1 => n38, B2 => n37, A => n36, ZN => n27);
   U82 : XOR2_X1 port map( A => A(25), B => B(25), Z => n28);
   U83 : XOR2_X1 port map( A => carry_25_port, B => n28, Z => SUM(25));
   U84 : NAND2_X1 port map( A1 => carry_25_port, A2 => A(25), ZN => n29);
   U85 : NAND2_X1 port map( A1 => carry_25_port, A2 => B(25), ZN => n30);
   U86 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n31);
   U87 : NAND3_X1 port map( A1 => n29, A2 => n30, A3 => n31, ZN => 
                           carry_26_port);
   U88 : NAND2_X1 port map( A1 => B(58), A2 => n163, ZN => net60811);
   U89 : INV_X1 port map( A => A(58), ZN => n32);
   U90 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n33);
   U91 : OAI21_X1 port map( B1 => n170, B2 => n74, A => n75, ZN => n34);
   U92 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n68);
   U93 : XNOR2_X1 port map( A => n27, B => B(55), ZN => net60816);
   U94 : INV_X1 port map( A => A(54), ZN => n38);
   U95 : OAI21_X1 port map( B1 => n37, B2 => net60698, A => n36, ZN => net60849
                           );
   U96 : NOR2_X1 port map( A1 => net60848, A2 => B(54), ZN => n37);
   U97 : NAND2_X1 port map( A1 => net60848, A2 => B(54), ZN => n36);
   U98 : OAI21_X1 port map( B1 => net60698, B2 => n35, A => n36, ZN => net60696
                           );
   U99 : INV_X1 port map( A => A(54), ZN => net60698);
   U100 : NOR2_X1 port map( A1 => net60847, A2 => B(54), ZN => n35);
   U101 : XNOR2_X1 port map( A => net60847, B => B(54), ZN => net60817);
   U102 : XNOR2_X1 port map( A => net60816, B => net60903, ZN => SUM(55));
   U103 : NAND2_X1 port map( A1 => B(55), A2 => net60849, ZN => net60705);
   U104 : NOR2_X1 port map( A1 => net60696, A2 => B(55), ZN => net74645);
   U105 : INV_X1 port map( A => net60704, ZN => net60903);
   U106 : INV_X1 port map( A => A(55), ZN => net60704);
   U107 : OAI21_X1 port map( B1 => net74645, B2 => net60704, A => net60705, ZN 
                           => net60702);
   U108 : OAI21_X1 port map( B1 => n23, B2 => net60704, A => net60705, ZN => 
                           net60859);
   U109 : OAI21_X1 port map( B1 => n85, B2 => n84, A => n86, ZN => n39);
   U110 : OAI21_X1 port map( B1 => n85, B2 => n84, A => n86, ZN => n174);
   U111 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => n40);
   U112 : NOR2_X1 port map( A1 => n95, A2 => B(40), ZN => n41);
   U113 : NAND2_X1 port map( A1 => net75572, A2 => net60657, ZN => n42);
   U114 : CLKBUF_X1 port map( A => A(34), Z => n43);
   U115 : BUF_X1 port map( A => A(56), Z => n175);
   U116 : INV_X1 port map( A => A(33), ZN => n45);
   U117 : AND2_X1 port map( A1 => n81, A2 => n133, ZN => n46);
   U118 : XNOR2_X1 port map( A => n154, B => n85, ZN => SUM(36));
   U119 : INV_X1 port map( A => A(36), ZN => n85);
   U120 : XNOR2_X1 port map( A => n42, B => n136, ZN => n149);
   U121 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => n47);
   U122 : NOR2_X1 port map( A1 => n172, A2 => B(53), ZN => n48);
   U123 : NOR2_X1 port map( A1 => n114, A2 => B(52), ZN => n49);
   U124 : INV_X1 port map( A => A(57), ZN => n128);
   U125 : NOR2_X1 port map( A1 => B(50), A2 => n164, ZN => n50);
   U126 : CLKBUF_X1 port map( A => A(35), Z => n51);
   U127 : OAI21_X1 port map( B1 => n52, B2 => n53, A => n54, ZN => 
                           carry_60_port);
   U128 : NAND2_X1 port map( A1 => B(59), A2 => n55, ZN => n54);
   U129 : NOR2_X1 port map( A1 => n55, A2 => B(59), ZN => n53);
   U130 : INV_X1 port map( A => A(59), ZN => n52);
   U131 : XNOR2_X1 port map( A => n56, B => B(59), ZN => net60812);
   U132 : OAI21_X1 port map( B1 => net60806, B2 => n32, A => net60811, ZN => 
                           n55);
   U133 : INV_X1 port map( A => n32, ZN => net61044);
   U134 : OAI21_X1 port map( B1 => n32, B2 => net60806, A => net60811, ZN => 
                           n56);
   U135 : XNOR2_X1 port map( A => n24, B => n150, ZN => SUM(40));
   U136 : NOR2_X1 port map( A1 => n165, A2 => B(38), ZN => n57);
   U137 : NOR2_X1 port map( A1 => n102, A2 => B(49), ZN => n58);
   U138 : XNOR2_X1 port map( A => n159, B => n66, ZN => SUM(31));
   U139 : NAND2_X1 port map( A1 => B(36), A2 => n80, ZN => n86);
   U140 : XNOR2_X1 port map( A => n153, B => n1, ZN => SUM(37));
   U141 : XNOR2_X1 port map( A => net60827, B => net84712, ZN => SUM(44));
   U142 : XNOR2_X1 port map( A => net60826, B => net84833, ZN => SUM(45));
   U143 : XNOR2_X1 port map( A => n149, B => n104, ZN => SUM(48));
   U144 : XNOR2_X1 port map( A => n40, B => n135, ZN => n150);
   U145 : NAND2_X1 port map( A1 => n95, A2 => B(40), ZN => n100);
   U146 : NAND2_X1 port map( A1 => n123, A2 => B(57), ZN => n129);
   U147 : XNOR2_X1 port map( A => n144, B => n121, ZN => SUM(53));
   U148 : XNOR2_X1 port map( A => n151, B => n177, ZN => SUM(39));
   U149 : NAND2_X1 port map( A1 => net60658, A2 => net60657, ZN => n101);
   U150 : INV_X1 port map( A => A(33), ZN => n74);
   U151 : INV_X1 port map( A => n93, ZN => n59);
   U152 : INV_X1 port map( A => A(38), ZN => n93);
   U153 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => n60);
   U154 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => n123);
   U155 : INV_X1 port map( A => net60652, ZN => net61029);
   U156 : XNOR2_X1 port map( A => n145, B => n26, ZN => SUM(52));
   U157 : XNOR2_X1 port map( A => n148, B => n44, ZN => SUM(49));
   U158 : INV_X1 port map( A => A(48), ZN => n104);
   U159 : NAND2_X1 port map( A1 => n96, A2 => n25, ZN => n95);
   U160 : NAND2_X1 port map( A1 => n42, A2 => B(48), ZN => n105);
   U161 : INV_X1 port map( A => A(52), ZN => n118);
   U162 : XNOR2_X1 port map( A => n80, B => n133, ZN => n154);
   U163 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n80);
   U164 : NOR2_X1 port map( A1 => B(33), A2 => n68, ZN => n73);
   U165 : OAI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n72);
   U166 : OAI21_X1 port map( B1 => n170, B2 => n45, A => n75, ZN => n161);
   U167 : NOR2_X1 port map( A1 => B(57), A2 => n123, ZN => n127);
   U168 : OAI21_X1 port map( B1 => n171, B2 => n128, A => n129, ZN => n126);
   U169 : OAI21_X1 port map( B1 => n127, B2 => n128, A => n129, ZN => n162);
   U170 : OAI21_X1 port map( B1 => n128, B2 => n127, A => n129, ZN => n163);
   U171 : NOR2_X1 port map( A1 => B(58), A2 => n126, ZN => net60806);
   U172 : NOR2_X1 port map( A1 => B(53), A2 => n117, ZN => n120);
   U173 : OAI21_X1 port map( B1 => n121, B2 => n48, A => n122, ZN => net60848);
   U174 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => net60847)
                           ;
   U175 : OAI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n106);
   U176 : NAND2_X1 port map( A1 => n106, A2 => B(50), ZN => n113);
   U177 : XNOR2_X1 port map( A => n106, B => B(50), ZN => n147);
   U178 : NOR2_X1 port map( A1 => n164, A2 => B(50), ZN => n111);
   U179 : NOR2_X1 port map( A1 => n173, A2 => B(49), ZN => n107);
   U180 : OAI21_X1 port map( B1 => n58, B2 => n108, A => n109, ZN => n164);
   U181 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n87);
   U182 : NAND2_X1 port map( A1 => n165, A2 => B(38), ZN => n94);
   U183 : XNOR2_X1 port map( A => n87, B => B(38), ZN => n152);
   U184 : NOR2_X1 port map( A1 => n87, A2 => B(38), ZN => n92);
   U185 : NOR2_X1 port map( A1 => n83, A2 => B(37), ZN => n88);
   U186 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n165);
   U187 : OAI21_X1 port map( B1 => n111, B2 => n112, A => n113, ZN => n110);
   U188 : NAND2_X1 port map( A1 => n110, A2 => B(51), ZN => n115);
   U189 : OAI21_X1 port map( B1 => n110, B2 => B(51), A => A(51), ZN => n116);
   U190 : XNOR2_X1 port map( A => n166, B => B(51), ZN => n146);
   U191 : OAI21_X1 port map( B1 => n50, B2 => n112, A => n113, ZN => n166);
   U192 : OAI21_X1 port map( B1 => n92, B2 => n93, A => n94, ZN => n91);
   U193 : NAND2_X1 port map( A1 => n167, A2 => B(39), ZN => n96);
   U194 : OAI21_X1 port map( B1 => n91, B2 => B(39), A => A(39), ZN => n97);
   U195 : XNOR2_X1 port map( A => n167, B => B(39), ZN => n151);
   U196 : OAI21_X1 port map( B1 => n57, B2 => n3, A => n94, ZN => n167);
   U197 : OAI21_X1 port map( B1 => n78, B2 => n77, A => n79, ZN => n76);
   U198 : NOR2_X1 port map( A1 => n72, A2 => B(34), ZN => n77);
   U199 : OAI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n168);
   U200 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n64);
   U201 : XNOR2_X1 port map( A => n169, B => n131, ZN => n158);
   U202 : NAND2_X1 port map( A1 => n169, A2 => B(32), ZN => n71);
   U203 : NOR2_X1 port map( A1 => B(32), A2 => n64, ZN => n69);
   U204 : NOR2_X1 port map( A1 => n61, A2 => B(31), ZN => n65);
   U205 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n169);
   U206 : NOR2_X1 port map( A1 => n33, A2 => B(33), ZN => n170);
   U207 : XNOR2_X1 port map( A => n33, B => n132, ZN => n157);
   U208 : NAND2_X1 port map( A1 => n68, A2 => B(33), ZN => n75);
   U209 : NOR2_X1 port map( A1 => B(57), A2 => n60, ZN => n171);
   U210 : XNOR2_X1 port map( A => net60817, B => net60885, ZN => SUM(54));
   U211 : XNOR2_X1 port map( A => n162, B => B(58), ZN => n141);
   U212 : XNOR2_X1 port map( A => net60702, B => B(56), ZN => n143);
   U213 : NAND2_X1 port map( A1 => net60859, A2 => B(56), ZN => n124);
   U214 : OAI21_X1 port map( B1 => n49, B2 => n118, A => n119, ZN => n117);
   U215 : OAI21_X1 port map( B1 => n49, B2 => n118, A => n119, ZN => n172);
   U216 : XNOR2_X1 port map( A => n117, B => n139, ZN => n144);
   U217 : NAND2_X1 port map( A1 => n172, A2 => B(53), ZN => n122);
   U218 : XNOR2_X1 port map( A => n147, B => n178, ZN => SUM(50));
   U219 : OAI21_X1 port map( B1 => n104, B2 => n103, A => n105, ZN => n102);
   U220 : XNOR2_X1 port map( A => n102, B => n137, ZN => n148);
   U221 : NAND2_X1 port map( A1 => n173, A2 => B(49), ZN => n109);
   U222 : NOR2_X1 port map( A1 => n101, A2 => B(48), ZN => n103);
   U223 : OAI21_X1 port map( B1 => n104, B2 => n103, A => n105, ZN => n173);
   U224 : XNOR2_X1 port map( A => net60825, B => net61029, ZN => SUM(46));
   U225 : XNOR2_X1 port map( A => net60829, B => A(42), ZN => SUM(42));
   U226 : OAI21_X1 port map( B1 => n41, B2 => n99, A => n100, ZN => net60615);
   U227 : XNOR2_X1 port map( A => net60871, B => net60777, ZN => net60830);
   U228 : XNOR2_X1 port map( A => n168, B => B(35), ZN => n155);
   U229 : NAND2_X1 port map( A1 => n168, A2 => B(35), ZN => n81);
   U230 : NOR2_X1 port map( A1 => n40, A2 => B(40), ZN => n98);
   U231 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => net60871);
   U232 : XNOR2_X1 port map( A => n152, B => n59, ZN => SUM(38));
   U233 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n83);
   U234 : XNOR2_X1 port map( A => n39, B => n134, ZN => n153);
   U235 : NAND2_X1 port map( A1 => B(37), A2 => n174, ZN => n90);
   U236 : XNOR2_X1 port map( A => n157, B => n45, ZN => SUM(33));
   U237 : INV_X1 port map( A => A(32), ZN => n70);
   U238 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n62);
   U239 : OAI21_X1 port map( B1 => A(30), B2 => B(30), A => carry_30_port, ZN 
                           => n63);
   U240 : XNOR2_X1 port map( A => n160, B => n10, ZN => SUM(30));
   U241 : XNOR2_X1 port map( A => n158, B => n70, ZN => SUM(32));
   U242 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n61);
   U243 : OAI21_X1 port map( B1 => net60859, B2 => B(56), A => A(56), ZN => 
                           n125);
   U244 : XNOR2_X1 port map( A => n143, B => n175, ZN => SUM(56));
   U245 : XNOR2_X1 port map( A => n61, B => n130, ZN => n159);
   U246 : NAND2_X1 port map( A1 => B(31), A2 => n61, ZN => n67);
   U247 : XNOR2_X1 port map( A => n156, B => n43, ZN => SUM(34));
   U248 : INV_X1 port map( A => A(34), ZN => n78);
   U249 : XNOR2_X1 port map( A => n155, B => n51, ZN => SUM(35));
   U250 : XNOR2_X1 port map( A => carry_30_port, B => B(30), ZN => n160);
   U251 : XNOR2_X1 port map( A => n146, B => n176, ZN => SUM(51));
   U252 : NAND2_X1 port map( A1 => B(34), A2 => n161, ZN => n79);
   U253 : XNOR2_X1 port map( A => net60828, B => net60892, ZN => SUM(43));
   U254 : INV_X1 port map( A => A(53), ZN => n121);
   U255 : XNOR2_X1 port map( A => net61044, B => n141, ZN => SUM(58));
   U256 : INV_X1 port map( A => n38, ZN => net60885);
   U257 : XNOR2_X1 port map( A => n34, B => B(34), ZN => n156);
   U258 : OAI21_X1 port map( B1 => B(35), B2 => n76, A => A(35), ZN => n82);
   U259 : CLKBUF_X1 port map( A => A(39), Z => n177);
   U260 : XNOR2_X1 port map( A => n60, B => n140, ZN => n142);
   U261 : XNOR2_X1 port map( A => n142, B => n128, ZN => SUM(57));
   U262 : INV_X1 port map( A => A(49), ZN => n108);
   U263 : NAND2_X1 port map( A1 => n115, A2 => n116, ZN => n114);
   U264 : INV_X1 port map( A => A(50), ZN => n112);
   U265 : INV_X1 port map( A => n112, ZN => n178);
   U266 : XNOR2_X1 port map( A => n47, B => n138, ZN => n145);
   U267 : NAND2_X1 port map( A1 => n47, A2 => B(52), ZN => n119);
   U268 : INV_X1 port map( A => A(40), ZN => n99);
   U269 : INV_X1 port map( A => A(37), ZN => n89);
   U270 : XNOR2_X1 port map( A => net60812, B => A(59), ZN => SUM(59));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_5_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_5_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_5_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port,
      carry_1_port, net51234, net51231, net51226, net51215, net51200, net51188,
      net51167, net51160, net51121, net51120, net51119, net51069, net51068, 
      net51067, net51054, net51049, net51005, net51004, net50993, net50985, 
      net50970, carry_9_port, carry_8_port, carry_7_port, carry_23_port, 
      carry_22_port, carry_21_port, carry_20_port, carry_19_port, carry_18_port
      , carry_17_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, net61068, 
      net61034, net51265, net51206, net51106, net68356, net51115, net51114, 
      net51113, net74679, net75138, net75523, net75556, net51257, net68330, 
      net51214, net51060, net51284, net51233, net51154, net50959, net50951, 
      net50950, net61040, net75358, net51230, net50977, net51228, net84534, 
      net75472, net74817, net50975, net50971, net50968, net50952, carry_34_port
      , carry_33_port, carry_32_port, carry_31_port, carry_30_port, 
      carry_29_port, carry_28_port, carry_27_port, carry_26_port, carry_25_port
      , carry_24_port, net75305, net51249, net51225, net50999, net50997, 
      net51232, net50969, net50965, net50964, net50963, net50962, net51260, 
      net50987, net68359, net51253, net51157, net50956, net84442, net74818, 
      net68267, net51242, net51000, net50998, net50994, net50992, net50991, 
      net51164, net50988, net50980, net84709, net84699, net75357, net51250, 
      net50982, net50981, net50976, net50974, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146 : std_logic;

begin
   
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1 : INV_X1 port map( A => net50976, ZN => n1);
   U2 : CLKBUF_X1 port map( A => net51114, Z => n2);
   U3 : INV_X1 port map( A => A(59), ZN => n3);
   U4 : INV_X1 port map( A => B(52), ZN => n28);
   U5 : INV_X1 port map( A => B(57), ZN => n118);
   U6 : INV_X1 port map( A => B(36), ZN => net51157);
   U7 : INV_X1 port map( A => B(37), ZN => net51160);
   U8 : INV_X1 port map( A => B(40), ZN => net51164);
   U9 : INV_X1 port map( A => B(53), ZN => net51188);
   U10 : INV_X1 port map( A => A(35), ZN => n8);
   U11 : INV_X1 port map( A => B(48), ZN => n115);
   U12 : INV_X1 port map( A => B(49), ZN => n116);
   U13 : INV_X1 port map( A => B(58), ZN => n44);
   U14 : INV_X1 port map( A => B(61), ZN => net51200);
   U15 : INV_X1 port map( A => B(45), ZN => n114);
   U16 : NAND2_X1 port map( A1 => B(63), A2 => n42, ZN => net51121);
   U17 : NOR2_X1 port map( A1 => B(63), A2 => n42, ZN => net51119);
   U18 : OAI21_X1 port map( B1 => net51119, B2 => net51120, A => net51121, ZN 
                           => SUM(64));
   U19 : INV_X1 port map( A => B(35), ZN => net51154);
   U20 : INV_X1 port map( A => B(56), ZN => n117);
   U21 : OAI21_X1 port map( B1 => net50963, B2 => net50964, A => net50965, ZN 
                           => net61040);
   U22 : INV_X1 port map( A => B(44), ZN => n113);
   U23 : INV_X1 port map( A => B(41), ZN => net51167);
   U24 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n139);
   U25 : NAND2_X1 port map( A1 => net50982, A2 => net50981, ZN => net75357);
   U26 : XNOR2_X1 port map( A => net75357, B => net51164, ZN => net51228);
   U27 : NAND2_X1 port map( A1 => net75357, A2 => B(40), ZN => net50988);
   U28 : OAI21_X1 port map( B1 => net84699, B2 => B(39), A => A(39), ZN => 
                           net50982);
   U29 : NAND2_X1 port map( A1 => net50974, A2 => B(39), ZN => net50981);
   U30 : NAND2_X1 port map( A1 => net84709, A2 => net50981, ZN => net50980);
   U31 : OAI21_X1 port map( B1 => net50976, B2 => net50975, A => net50977, ZN 
                           => net50974);
   U32 : INV_X1 port map( A => A(38), ZN => net50976);
   U33 : OAI21_X1 port map( B1 => net75358, B2 => net50976, A => net50977, ZN 
                           => net51250);
   U34 : OAI21_X1 port map( B1 => net50975, B2 => net50976, A => net50977, ZN 
                           => net84699);
   U35 : OAI21_X1 port map( B1 => net84699, B2 => B(39), A => A(39), ZN => 
                           net84709);
   U36 : XNOR2_X1 port map( A => net51250, B => B(39), ZN => n4);
   U37 : XNOR2_X1 port map( A => n4, B => A(39), ZN => SUM(39));
   U38 : XNOR2_X1 port map( A => net51230, B => n1, ZN => SUM(38));
   U39 : OAI21_X1 port map( B1 => n5, B2 => net50987, A => net50988, ZN => 
                           net51260);
   U40 : OAI21_X1 port map( B1 => n6, B2 => net50987, A => net50988, ZN => 
                           net50985);
   U41 : NOR2_X1 port map( A1 => net50980, A2 => B(40), ZN => n6);
   U42 : NOR2_X1 port map( A1 => net50980, A2 => B(40), ZN => n5);
   U43 : NAND2_X1 port map( A1 => net50991, A2 => B(42), ZN => net51000);
   U44 : OAI21_X1 port map( B1 => net74818, B2 => net50999, A => net51000, ZN 
                           => net51249);
   U45 : OAI21_X1 port map( B1 => net50999, B2 => net50998, A => net51000, ZN 
                           => net50997);
   U46 : OAI21_X1 port map( B1 => net50992, B2 => net84442, A => net50994, ZN 
                           => net50991);
   U47 : NOR2_X1 port map( A1 => net50991, A2 => B(42), ZN => net50998);
   U48 : NOR2_X1 port map( A1 => net50991, A2 => B(42), ZN => net74818);
   U49 : INV_X1 port map( A => A(41), ZN => net84442);
   U50 : NOR2_X1 port map( A1 => net51260, A2 => B(41), ZN => net50992);
   U51 : XNOR2_X1 port map( A => B(42), B => net51242, ZN => net51226);
   U52 : OAI21_X1 port map( B1 => net68267, B2 => net50993, A => net50994, ZN 
                           => net51242);
   U53 : INV_X1 port map( A => A(41), ZN => net50993);
   U54 : NAND2_X1 port map( A1 => net51260, A2 => B(41), ZN => net50994);
   U55 : NOR2_X1 port map( A1 => B(41), A2 => net50985, ZN => net68267);
   U56 : NOR2_X1 port map( A1 => net50956, A2 => B(36), ZN => net68359);
   U57 : OAI21_X1 port map( B1 => net68359, B2 => net50964, A => net50965, ZN 
                           => net50962);
   U58 : OAI21_X1 port map( B1 => n7, B2 => n8, A => net50959, ZN => net50956);
   U59 : XNOR2_X1 port map( A => net50956, B => net51157, ZN => net51232);
   U60 : XNOR2_X1 port map( A => net51233, B => n8, ZN => SUM(35));
   U61 : OAI21_X1 port map( B1 => n9, B2 => n8, A => net50959, ZN => net51253);
   U62 : AND2_X1 port map( A1 => net51284, A2 => net50951, ZN => n7);
   U63 : NOR2_X1 port map( A1 => net51253, A2 => B(36), ZN => net50963);
   U64 : NAND2_X1 port map( A1 => net51253, A2 => B(36), ZN => net50965);
   U65 : AND2_X1 port map( A1 => net51284, A2 => net50951, ZN => n9);
   U66 : NAND2_X1 port map( A1 => net50952, A2 => net50951, ZN => net50950);
   U67 : INV_X1 port map( A => A(40), ZN => net50987);
   U68 : XNOR2_X1 port map( A => net51228, B => net50987, ZN => SUM(40));
   U69 : NOR2_X1 port map( A1 => net50962, A2 => B(37), ZN => net50969);
   U70 : OAI21_X1 port map( B1 => net50969, B2 => net74817, A => net50971, ZN 
                           => net75472);
   U71 : NOR2_X1 port map( A1 => B(37), A2 => net50962, ZN => net84534);
   U72 : INV_X1 port map( A => A(36), ZN => net50964);
   U73 : XNOR2_X1 port map( A => net51232, B => net50964, ZN => SUM(36));
   U74 : XNOR2_X1 port map( A => net50997, B => B(43), ZN => net51225);
   U75 : XNOR2_X1 port map( A => net51225, B => net75305, ZN => SUM(43));
   U76 : NAND2_X1 port map( A1 => net50997, A2 => B(43), ZN => net51004);
   U77 : INV_X1 port map( A => A(42), ZN => net50999);
   U78 : INV_X1 port map( A => net50999, ZN => net75556);
   U79 : OAI21_X1 port map( B1 => net51249, B2 => B(43), A => A(43), ZN => 
                           net75138);
   U80 : OAI21_X1 port map( B1 => net51249, B2 => B(43), A => A(43), ZN => 
                           net51005);
   U81 : CLKBUF_X1 port map( A => A(43), Z => net75305);
   U82 : OAI21_X1 port map( B1 => A(34), B2 => B(34), A => carry_34_port, ZN =>
                           net50952);
   U83 : AND2_X1 port map( A1 => net50952, A2 => net51154, ZN => net51284);
   U84 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => net50951);
   U85 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => net51234);
   U86 : CLKBUF_X1 port map( A => carry_34_port, Z => net74679);
   U87 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => 
                           carry_24_port);
   U88 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n13);
   U89 : NAND2_X1 port map( A1 => carry_23_port, A2 => B(23), ZN => n12);
   U90 : NAND2_X1 port map( A1 => carry_23_port, A2 => A(23), ZN => n11);
   U91 : XOR2_X1 port map( A => A(23), B => B(23), Z => n10);
   U92 : XOR2_X1 port map( A => carry_23_port, B => n10, Z => SUM(23));
   U93 : NOR2_X1 port map( A1 => net75472, A2 => B(38), ZN => net50975);
   U94 : NOR2_X1 port map( A1 => B(38), A2 => net75472, ZN => net75358);
   U95 : NAND2_X1 port map( A1 => net61040, A2 => B(37), ZN => net50971);
   U96 : INV_X1 port map( A => A(37), ZN => net74817);
   U97 : OAI21_X1 port map( B1 => net84534, B2 => net74817, A => net50971, ZN 
                           => net50968);
   U98 : NAND2_X1 port map( A1 => B(38), A2 => net50968, ZN => net50977);
   U99 : XNOR2_X1 port map( A => net50968, B => B(38), ZN => net51230);
   U100 : XNOR2_X1 port map( A => net61040, B => net51160, ZN => net51231);
   U101 : INV_X1 port map( A => A(37), ZN => net50970);
   U102 : NAND2_X1 port map( A1 => B(35), A2 => net50950, ZN => net50959);
   U103 : XNOR2_X1 port map( A => net50950, B => net51154, ZN => net51233);
   U104 : CLKBUF_X1 port map( A => A(62), Z => net61034);
   U105 : OAI21_X1 port map( B1 => n26, B2 => n25, A => n27, ZN => n14);
   U106 : OAI21_X1 port map( B1 => n47, B2 => n66, A => n67, ZN => n15);
   U107 : OAI21_X1 port map( B1 => n26, B2 => n25, A => n27, ZN => net51054);
   U108 : NOR2_X1 port map( A1 => n32, A2 => B(48), ZN => n16);
   U109 : NOR2_X1 port map( A1 => n145, A2 => B(46), ZN => n17);
   U110 : CLKBUF_X1 port map( A => n79, Z => n18);
   U111 : OAI21_X1 port map( B1 => n24, B2 => n21, A => n22, ZN => n19);
   U112 : XNOR2_X1 port map( A => n19, B => B(54), ZN => net51214);
   U113 : XNOR2_X1 port map( A => net51214, B => net68330, ZN => SUM(54));
   U114 : OAI21_X1 port map( B1 => n24, B2 => n21, A => n22, ZN => n23);
   U115 : NAND2_X1 port map( A1 => n23, A2 => B(54), ZN => net51069);
   U116 : INV_X1 port map( A => A(53), ZN => n21);
   U117 : XNOR2_X1 port map( A => net51215, B => n21, ZN => SUM(53));
   U118 : OAI21_X1 port map( B1 => n20, B2 => n21, A => n22, ZN => net51060);
   U119 : NOR2_X1 port map( A1 => B(53), A2 => net51257, ZN => n24);
   U120 : NOR2_X1 port map( A1 => net51060, A2 => B(54), ZN => net68356);
   U121 : NOR2_X1 port map( A1 => net51060, A2 => B(54), ZN => net51067);
   U122 : NAND2_X1 port map( A1 => net51257, A2 => B(53), ZN => n22);
   U123 : NOR2_X1 port map( A1 => n14, A2 => B(53), ZN => n20);
   U124 : CLKBUF_X1 port map( A => A(54), Z => net68330);
   U125 : INV_X1 port map( A => A(54), ZN => net51068);
   U126 : OAI21_X1 port map( B1 => n30, B2 => n26, A => n27, ZN => net51257);
   U127 : INV_X1 port map( A => A(52), ZN => n26);
   U128 : XNOR2_X1 port map( A => n29, B => n26, ZN => SUM(52));
   U129 : NOR2_X1 port map( A1 => B(52), A2 => net75523, ZN => n30);
   U130 : NAND2_X1 port map( A1 => net51049, A2 => B(52), ZN => n27);
   U131 : NOR2_X1 port map( A1 => B(52), A2 => net51049, ZN => n25);
   U132 : XNOR2_X1 port map( A => net75523, B => n28, ZN => n29);
   U133 : OAI21_X1 port map( B1 => B(51), B2 => n85, A => A(51), ZN => n31);
   U134 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => n32);
   U135 : NAND2_X1 port map( A1 => n89, A2 => n31, ZN => net75523);
   U136 : AND2_X1 port map( A1 => n33, A2 => n94, ZN => n96);
   U137 : AND2_X1 port map( A1 => n93, A2 => n117, ZN => n33);
   U138 : CLKBUF_X1 port map( A => A(55), Z => n34);
   U139 : NAND2_X1 port map( A1 => net51004, A2 => net75138, ZN => n35);
   U140 : INV_X1 port map( A => n87, ZN => n36);
   U141 : NOR2_X1 port map( A1 => n64, A2 => B(45), ZN => n37);
   U142 : OAI21_X1 port map( B1 => n68, B2 => n69, A => n70, ZN => n38);
   U143 : NOR2_X1 port map( A1 => B(61), A2 => net61068, ZN => n39);
   U144 : XNOR2_X1 port map( A => n41, B => A(63), ZN => SUM(63));
   U145 : XNOR2_X1 port map( A => n40, B => B(63), ZN => n41);
   U146 : OAI21_X1 port map( B1 => net51114, B2 => net51113, A => net51115, ZN 
                           => n40);
   U147 : INV_X1 port map( A => A(62), ZN => net51114);
   U148 : NOR2_X1 port map( A1 => net51265, A2 => B(62), ZN => net51113);
   U149 : OAI21_X1 port map( B1 => net51113, B2 => n2, A => net51115, ZN => n42
                           );
   U150 : NAND2_X1 port map( A1 => net51265, A2 => B(62), ZN => net51115);
   U151 : XNOR2_X1 port map( A => net51106, B => B(62), ZN => net51206);
   U152 : CLKBUF_X1 port map( A => A(47), Z => n43);
   U153 : BUF_X1 port map( A => A(60), Z => n60);
   U154 : XNOR2_X1 port map( A => n142, B => n44, ZN => n45);
   U155 : XNOR2_X1 port map( A => n45, B => n56, ZN => SUM(58));
   U156 : NOR2_X1 port map( A1 => n81, A2 => B(50), ZN => n46);
   U157 : NOR2_X1 port map( A1 => n63, A2 => B(44), ZN => n47);
   U158 : NAND2_X1 port map( A1 => n134, A2 => B(59), ZN => n48);
   U159 : INV_X1 port map( A => A(49), ZN => n83);
   U160 : OAI21_X1 port map( B1 => n104, B2 => n56, A => n105, ZN => n49);
   U161 : OAI21_X1 port map( B1 => n59, B2 => n141, A => n105, ZN => n103);
   U162 : INV_X1 port map( A => A(63), ZN => net51120);
   U163 : CLKBUF_X1 port map( A => A(51), Z => n50);
   U164 : INV_X1 port map( A => A(48), ZN => n79);
   U165 : XNOR2_X1 port map( A => net61034, B => net51206, ZN => SUM(62));
   U166 : OAI21_X1 port map( B1 => n39, B2 => n52, A => n53, ZN => net51106);
   U167 : INV_X1 port map( A => A(61), ZN => n52);
   U168 : OAI21_X1 port map( B1 => n52, B2 => n51, A => n53, ZN => net51265);
   U169 : NOR2_X1 port map( A1 => B(61), A2 => net61068, ZN => n51);
   U170 : NAND2_X1 port map( A1 => B(61), A2 => net61068, ZN => n53);
   U171 : NOR2_X1 port map( A1 => n49, A2 => B(59), ZN => n54);
   U172 : INV_X1 port map( A => A(57), ZN => n55);
   U173 : INV_X1 port map( A => A(58), ZN => n56);
   U174 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => net61068);
   U175 : OAI21_X1 port map( B1 => n17, B2 => n72, A => n73, ZN => n57);
   U176 : OAI21_X1 port map( B1 => n72, B2 => n17, A => n73, ZN => n71);
   U177 : OAI21_X1 port map( B1 => n3, B2 => n54, A => n48, ZN => n58);
   U178 : INV_X1 port map( A => A(58), ZN => n59);
   U179 : NAND2_X1 port map( A1 => n134, A2 => B(59), ZN => n109);
   U180 : NOR2_X1 port map( A1 => n49, A2 => B(59), ZN => n61);
   U181 : XNOR2_X1 port map( A => n92, B => n117, ZN => n123);
   U182 : NAND2_X1 port map( A1 => n63, A2 => B(44), ZN => n67);
   U183 : XNOR2_X1 port map( A => n35, B => n113, ZN => n132);
   U184 : INV_X1 port map( A => A(56), ZN => n97);
   U185 : INV_X1 port map( A => n3, ZN => n62);
   U186 : OAI21_X1 port map( B1 => B(51), B2 => n85, A => A(51), ZN => n90);
   U187 : OAI21_X1 port map( B1 => B(60), B2 => n106, A => A(60), ZN => n112);
   U188 : XNOR2_X1 port map( A => net51234, B => net74679, ZN => SUM(34));
   U189 : XNOR2_X1 port map( A => n123, B => n97, ZN => SUM(56));
   U190 : INV_X1 port map( A => A(57), ZN => n101);
   U191 : XNOR2_X1 port map( A => n119, B => n52, ZN => SUM(61));
   U192 : XNOR2_X1 port map( A => n128, B => n18, ZN => SUM(48));
   U193 : XNOR2_X1 port map( A => net51231, B => net50970, ZN => SUM(37));
   U194 : XNOR2_X1 port map( A => n131, B => n69, ZN => SUM(45));
   U195 : XNOR2_X1 port map( A => n132, B => n66, ZN => SUM(44));
   U196 : NOR2_X1 port map( A1 => B(58), A2 => n99, ZN => n104);
   U197 : OAI21_X1 port map( B1 => n59, B2 => n141, A => n105, ZN => n134);
   U198 : OAI21_X1 port map( B1 => n56, B2 => n104, A => n105, ZN => n135);
   U199 : NOR2_X1 port map( A1 => B(49), A2 => n144, ZN => n82);
   U200 : OAI21_X1 port map( B1 => n82, B2 => n83, A => n84, ZN => n81);
   U201 : OAI21_X1 port map( B1 => n143, B2 => n83, A => n84, ZN => n136);
   U202 : NAND2_X1 port map( A1 => n38, A2 => B(46), ZN => n73);
   U203 : XNOR2_X1 port map( A => n38, B => B(46), ZN => n130);
   U204 : NOR2_X1 port map( A1 => n103, A2 => B(59), ZN => n107);
   U205 : OAI21_X1 port map( B1 => n61, B2 => n108, A => n48, ZN => n106);
   U206 : OAI21_X1 port map( B1 => n108, B2 => n107, A => n109, ZN => n137);
   U207 : XNOR2_X1 port map( A => n137, B => B(60), ZN => n120);
   U208 : NAND2_X1 port map( A1 => B(60), A2 => n58, ZN => n111);
   U209 : OAI21_X1 port map( B1 => net51067, B2 => net51068, A => net51069, ZN 
                           => n91);
   U210 : OAI21_X1 port map( B1 => net68356, B2 => net51068, A => net51069, ZN 
                           => n138);
   U211 : NOR2_X1 port map( A1 => n81, A2 => B(50), ZN => n86);
   U212 : OAI21_X1 port map( B1 => n46, B2 => n87, A => n88, ZN => n85);
   U213 : NAND2_X1 port map( A1 => n71, A2 => B(47), ZN => n75);
   U214 : OAI21_X1 port map( B1 => n57, B2 => B(47), A => A(47), ZN => n76);
   U215 : XNOR2_X1 port map( A => n71, B => B(47), ZN => n129);
   U216 : OAI21_X1 port map( B1 => n97, B2 => n96, A => n98, ZN => n95);
   U217 : XNOR2_X1 port map( A => n95, B => n118, ZN => n122);
   U218 : NAND2_X1 port map( A1 => n140, A2 => B(57), ZN => n102);
   U219 : NOR2_X1 port map( A1 => n140, A2 => B(57), ZN => n100);
   U220 : OAI21_X1 port map( B1 => n96, B2 => n97, A => n98, ZN => n140);
   U221 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n64);
   U222 : XNOR2_X1 port map( A => n15, B => n114, ZN => n131);
   U223 : NAND2_X1 port map( A1 => n15, A2 => B(45), ZN => n70);
   U224 : NOR2_X1 port map( A1 => n64, A2 => B(45), ZN => n68);
   U225 : NOR2_X1 port map( A1 => B(44), A2 => n35, ZN => n65);
   U226 : NOR2_X1 port map( A1 => n99, A2 => B(58), ZN => n141);
   U227 : OAI21_X1 port map( B1 => n101, B2 => n100, A => n102, ZN => n99);
   U228 : NAND2_X1 port map( A1 => n142, A2 => B(58), ZN => n105);
   U229 : OAI21_X1 port map( B1 => n100, B2 => n55, A => n102, ZN => n142);
   U230 : XNOR2_X1 port map( A => n138, B => B(55), ZN => n124);
   U231 : NAND2_X1 port map( A1 => n91, A2 => B(55), ZN => n93);
   U232 : XNOR2_X1 port map( A => net51054, B => net51188, ZN => net51215);
   U233 : NOR2_X1 port map( A1 => n77, A2 => B(49), ZN => n143);
   U234 : OAI21_X1 port map( B1 => n16, B2 => n79, A => n80, ZN => n77);
   U235 : XNOR2_X1 port map( A => n144, B => n116, ZN => n127);
   U236 : NAND2_X1 port map( A1 => n77, A2 => B(49), ZN => n84);
   U237 : NOR2_X1 port map( A1 => n74, A2 => B(48), ZN => n78);
   U238 : OAI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n144);
   U239 : XNOR2_X1 port map( A => n129, B => n43, ZN => SUM(47));
   U240 : XNOR2_X1 port map( A => B(59), B => n135, ZN => n121);
   U241 : XNOR2_X1 port map( A => n139, B => B(51), ZN => n125);
   U242 : NAND2_X1 port map( A1 => n139, A2 => B(51), ZN => n89);
   U243 : XNOR2_X1 port map( A => n136, B => B(50), ZN => n126);
   U244 : XNOR2_X1 port map( A => n121, B => n62, ZN => SUM(59));
   U245 : XNOR2_X1 port map( A => net50985, B => net51167, ZN => n133);
   U246 : NAND2_X1 port map( A1 => net51004, A2 => net51005, ZN => n63);
   U247 : NAND2_X1 port map( A1 => B(56), A2 => n92, ZN => n98);
   U248 : XNOR2_X1 port map( A => n130, B => n146, ZN => SUM(46));
   U249 : INV_X1 port map( A => A(46), ZN => n72);
   U250 : OAI21_X1 port map( B1 => n37, B2 => n69, A => n70, ZN => n145);
   U251 : XNOR2_X1 port map( A => n124, B => n34, ZN => SUM(55));
   U252 : XNOR2_X1 port map( A => n125, B => n50, ZN => SUM(51));
   U253 : XNOR2_X1 port map( A => n122, B => n101, ZN => SUM(57));
   U254 : XNOR2_X1 port map( A => net51226, B => net75556, ZN => SUM(42));
   U255 : XNOR2_X1 port map( A => n120, B => n60, ZN => SUM(60));
   U256 : OAI21_X1 port map( B1 => n91, B2 => B(55), A => A(55), ZN => n94);
   U257 : INV_X1 port map( A => A(45), ZN => n69);
   U258 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => net51049);
   U259 : XNOR2_X1 port map( A => n126, B => n36, ZN => SUM(50));
   U260 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => n110);
   U261 : XNOR2_X1 port map( A => n110, B => net51200, ZN => n119);
   U262 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U263 : INV_X1 port map( A => n72, ZN => n146);
   U264 : NAND2_X1 port map( A1 => n136, A2 => B(50), ZN => n88);
   U265 : INV_X1 port map( A => A(50), ZN => n87);
   U266 : XNOR2_X1 port map( A => n133, B => net50993, ZN => SUM(41));
   U267 : INV_X1 port map( A => A(59), ZN => n108);
   U268 : INV_X1 port map( A => A(44), ZN => n66);
   U269 : XNOR2_X1 port map( A => n127, B => n83, ZN => SUM(49));
   U270 : XNOR2_X1 port map( A => n32, B => n115, ZN => n128);
   U271 : NAND2_X1 port map( A1 => n74, A2 => B(48), ZN => n80);
   U272 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => n92);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_6_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_6_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_6_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port,
      carry_3_port, carry_2_port, carry_1_port, net68161, net68162, net68160, 
      net68157, net68121, net68033, net68026, net67980, net67969, net67872, 
      net67871, net68354, net68398, net68363, net68125, net68123, net68136, 
      net67977, net67975, net68177, net68135, net68103, net67983, net67982, 
      net67981, net67974, net84800, net74815, carry_34_port, carry_33_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347 : std_logic;

begin
   
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1 : INV_X1 port map( A => n204, ZN => n1);
   U2 : OAI21_X1 port map( B1 => B(55), B2 => n253, A => A(55), ZN => n2);
   U3 : BUF_X1 port map( A => carry_34_port, Z => net74815);
   U4 : BUF_X1 port map( A => n144, Z => n138);
   U5 : CLKBUF_X1 port map( A => n41, Z => n3);
   U6 : OAI21_X1 port map( B1 => n202, B2 => B(39), A => A(39), ZN => n4);
   U7 : OAI21_X2 port map( B1 => n63, B2 => n64, A => n65, ZN => n141);
   U8 : NOR2_X2 port map( A1 => B(29), A2 => n66, ZN => n71);
   U9 : NOR2_X2 port map( A1 => B(27), A2 => n59, ZN => n63);
   U10 : NAND2_X1 port map( A1 => B(31), A2 => n134, ZN => n89);
   U11 : NAND2_X1 port map( A1 => B(28), A2 => n142, ZN => n69);
   U12 : INV_X1 port map( A => B(53), ZN => net68103);
   U13 : NAND2_X1 port map( A1 => B(27), A2 => n137, ZN => n65);
   U14 : NAND2_X1 port map( A1 => B(30), A2 => n140, ZN => n77);
   U15 : INV_X1 port map( A => B(44), ZN => n287);
   U16 : INV_X1 port map( A => B(45), ZN => n288);
   U17 : INV_X1 port map( A => B(20), ZN => n40);
   U18 : INV_X1 port map( A => A(23), ZN => n49);
   U19 : INV_X1 port map( A => B(41), ZN => n286);
   U20 : NAND2_X1 port map( A1 => A(9), A2 => n91, ZN => n119);
   U21 : INV_X1 port map( A => n117, ZN => n8);
   U22 : NAND2_X1 port map( A1 => A(19), A2 => n107, ZN => n120);
   U23 : INV_X1 port map( A => B(22), ZN => n45);
   U24 : INV_X1 port map( A => B(36), ZN => n283);
   U25 : INV_X1 port map( A => B(37), ZN => n284);
   U26 : INV_X1 port map( A => B(52), ZN => n158);
   U27 : INV_X1 port map( A => B(56), ZN => n291);
   U28 : XNOR2_X1 port map( A => B(8), B => carry_8_port, ZN => n118);
   U29 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n90);
   U30 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => n91);
   U31 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n122);
   U32 : OAI21_X1 port map( B1 => A(8), B2 => B(8), A => carry_8_port, ZN => 
                           n121);
   U33 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n116);
   U34 : OAI211_X1 port map( C1 => n123, C2 => n80, A => n119, B => n124, ZN =>
                           n117);
   U35 : INV_X1 port map( A => n91, ZN => n123);
   U36 : INV_X1 port map( A => B(9), ZN => n80);
   U37 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n124);
   U38 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n115);
   U39 : OAI221_X1 port map( B1 => n8, B2 => n9, C1 => n8, C2 => n10, A => n11,
                           ZN => n7);
   U40 : INV_X1 port map( A => A(10), ZN => n9);
   U41 : INV_X1 port map( A => B(10), ZN => n10);
   U42 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n11);
   U43 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n114);
   U44 : OAI21_X1 port map( B1 => n13, B2 => n14, A => n15, ZN => n12);
   U45 : INV_X1 port map( A => A(11), ZN => n14);
   U46 : NAND2_X1 port map( A1 => B(11), A2 => n7, ZN => n15);
   U47 : NOR2_X1 port map( A1 => B(11), A2 => n7, ZN => n13);
   U48 : XNOR2_X1 port map( A => B(13), B => A(13), ZN => n113);
   U49 : OAI21_X1 port map( B1 => n17, B2 => n18, A => n19, ZN => n16);
   U50 : INV_X1 port map( A => A(12), ZN => n18);
   U51 : NAND2_X1 port map( A1 => B(12), A2 => n12, ZN => n19);
   U52 : NOR2_X1 port map( A1 => B(12), A2 => n12, ZN => n17);
   U53 : XNOR2_X1 port map( A => B(14), B => A(14), ZN => n112);
   U54 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => n20);
   U55 : NAND2_X1 port map( A1 => B(13), A2 => n16, ZN => n21);
   U56 : OAI21_X1 port map( B1 => B(13), B2 => n16, A => A(13), ZN => n22);
   U57 : XNOR2_X1 port map( A => B(15), B => A(15), ZN => n111);
   U58 : OAI21_X1 port map( B1 => n24, B2 => n25, A => n26, ZN => n23);
   U59 : INV_X1 port map( A => A(14), ZN => n25);
   U60 : NAND2_X1 port map( A1 => B(14), A2 => n20, ZN => n26);
   U61 : NOR2_X1 port map( A1 => B(14), A2 => n20, ZN => n24);
   U62 : XNOR2_X1 port map( A => B(16), B => A(16), ZN => n110);
   U63 : OAI21_X1 port map( B1 => n28, B2 => n29, A => n30, ZN => n27);
   U64 : INV_X1 port map( A => A(15), ZN => n29);
   U65 : NAND2_X1 port map( A1 => B(15), A2 => n23, ZN => n30);
   U66 : NOR2_X1 port map( A1 => B(15), A2 => n23, ZN => n28);
   U67 : XNOR2_X1 port map( A => B(17), B => A(17), ZN => n109);
   U68 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U69 : INV_X1 port map( A => A(16), ZN => n33);
   U70 : NAND2_X1 port map( A1 => B(16), A2 => n27, ZN => n34);
   U71 : NOR2_X1 port map( A1 => B(16), A2 => n27, ZN => n32);
   U72 : XNOR2_X1 port map( A => B(18), B => A(18), ZN => n108);
   U73 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n35);
   U74 : NAND2_X1 port map( A1 => B(17), A2 => n31, ZN => n36);
   U75 : OAI21_X1 port map( B1 => B(17), B2 => n31, A => A(17), ZN => n37);
   U76 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => n106);
   U77 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n125, ZN => n107);
   U78 : INV_X1 port map( A => A(18), ZN => n82);
   U79 : NAND2_X1 port map( A1 => B(18), A2 => n35, ZN => n125);
   U80 : NOR2_X1 port map( A1 => B(18), A2 => n35, ZN => n81);
   U81 : XNOR2_X1 port map( A => B(20), B => n131, ZN => n104);
   U82 : OAI211_X1 port map( C1 => n126, C2 => n83, A => n120, B => n127, ZN =>
                           n105);
   U83 : INV_X1 port map( A => n107, ZN => n126);
   U84 : INV_X1 port map( A => B(19), ZN => n83);
   U85 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n127);
   U86 : XNOR2_X1 port map( A => n101, B => n129, ZN => SUM(23));
   U87 : XNOR2_X1 port map( A => B(23), B => A(23), ZN => n101);
   U88 : NAND2_X1 port map( A1 => B(29), A2 => n135, ZN => n73);
   U89 : INV_X1 port map( A => B(35), ZN => n282);
   U90 : INV_X1 port map( A => B(48), ZN => n289);
   U91 : INV_X1 port map( A => B(49), ZN => n290);
   U92 : INV_X1 port map( A => B(61), ZN => n293);
   U93 : XNOR2_X1 port map( A => A(8), B => n118, ZN => SUM(8));
   U94 : XNOR2_X1 port map( A => n90, B => n91, ZN => SUM(9));
   U95 : XNOR2_X1 port map( A => n116, B => n117, ZN => SUM(10));
   U96 : XNOR2_X1 port map( A => n115, B => n7, ZN => SUM(11));
   U97 : XNOR2_X1 port map( A => n114, B => n12, ZN => SUM(12));
   U98 : XNOR2_X1 port map( A => n113, B => n16, ZN => SUM(13));
   U99 : XNOR2_X1 port map( A => n112, B => n20, ZN => SUM(14));
   U100 : XNOR2_X1 port map( A => n111, B => n23, ZN => SUM(15));
   U101 : XNOR2_X1 port map( A => n110, B => n27, ZN => SUM(16));
   U102 : XNOR2_X1 port map( A => n109, B => n31, ZN => SUM(17));
   U103 : XNOR2_X1 port map( A => n108, B => n35, ZN => SUM(18));
   U104 : XNOR2_X1 port map( A => n106, B => n107, ZN => SUM(19));
   U105 : XNOR2_X1 port map( A => n104, B => n105, ZN => SUM(20));
   U106 : XNOR2_X1 port map( A => n93, B => n133, ZN => SUM(31));
   U107 : INV_X1 port map( A => B(63), ZN => net68123);
   U108 : NAND2_X1 port map( A1 => net68033, A2 => n281, ZN => SUM(64));
   U109 : XOR2_X1 port map( A => B(21), B => A(21), Z => n5);
   U110 : XNOR2_X1 port map( A => n102, B => n147, ZN => SUM(22));
   U111 : NAND2_X1 port map( A1 => n207, A2 => n4, ZN => n6);
   U112 : INV_X1 port map( A => B(40), ZN => n285);
   U113 : INV_X1 port map( A => B(57), ZN => n292);
   U114 : XNOR2_X1 port map( A => n94, B => n70, ZN => SUM(30));
   U115 : XNOR2_X1 port map( A => n97, B => n136, ZN => SUM(27));
   U116 : OAI21_X1 port map( B1 => n215, B2 => n171, A => n216, ZN => n213);
   U117 : OAI21_X1 port map( B1 => n156, B2 => net67975, A => net67977, ZN => 
                           net67974);
   U118 : OAI21_X1 port map( B1 => n255, B2 => n254, A => n256, ZN => n330);
   U119 : OAI21_X2 port map( B1 => n52, B2 => n53, A => n54, ZN => n51);
   U120 : OAI21_X2 port map( B1 => n56, B2 => n57, A => n58, ZN => n55);
   U121 : OAI221_X1 port map( B1 => n43, B2 => n44, C1 => n43, C2 => n45, A => 
                           n46, ZN => n42);
   U122 : OAI221_X1 port map( B1 => n44, B2 => n43, C1 => n43, C2 => n45, A => 
                           n46, ZN => n129);
   U123 : OAI221_X1 port map( B1 => n43, B2 => n44, C1 => n43, C2 => n45, A => 
                           n46, ZN => n130);
   U124 : INV_X1 port map( A => A(20), ZN => n41);
   U125 : INV_X1 port map( A => n3, ZN => n131);
   U126 : INV_X1 port map( A => n105, ZN => n39);
   U127 : OAI222_X1 port map( A1 => n39, A2 => n40, B1 => n39, B2 => n41, C1 =>
                           n41, C2 => n40, ZN => n38);
   U128 : OAI222_X1 port map( A1 => n39, A2 => n40, B1 => n39, B2 => n41, C1 =>
                           n41, C2 => n40, ZN => n132);
   U129 : NAND2_X1 port map( A1 => B(21), A2 => n132, ZN => n128);
   U130 : NOR2_X1 port map( A1 => n42, A2 => B(23), ZN => n48);
   U131 : NAND2_X1 port map( A1 => B(23), A2 => n130, ZN => n50);
   U132 : NOR2_X1 port map( A1 => n38, A2 => B(21), ZN => n85);
   U133 : CLKBUF_X1 port map( A => n132, Z => net84800);
   U134 : OAI21_X1 port map( B1 => n143, B2 => n76, A => n77, ZN => n74);
   U135 : NOR2_X1 port map( A1 => B(30), A2 => n140, ZN => n75);
   U136 : OAI21_X1 port map( B1 => n76, B2 => n75, A => n77, ZN => n133);
   U137 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => n134);
   U138 : NOR2_X1 port map( A1 => B(28), A2 => n142, ZN => n67);
   U139 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => n66);
   U140 : OAI21_X1 port map( B1 => n145, B2 => n68, A => n69, ZN => n135);
   U141 : NOR2_X1 port map( A1 => B(26), A2 => n55, ZN => n60);
   U142 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n59);
   U143 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n136);
   U144 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n137);
   U145 : NAND2_X1 port map( A1 => B(25), A2 => n51, ZN => n58);
   U146 : XNOR2_X1 port map( A => n99, B => n51, ZN => SUM(25));
   U147 : NOR2_X1 port map( A1 => B(25), A2 => n51, ZN => n56);
   U148 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => n47);
   U149 : NAND2_X1 port map( A1 => B(24), A2 => n144, ZN => n54);
   U150 : XNOR2_X1 port map( A => n100, B => n138, ZN => SUM(24));
   U151 : NOR2_X1 port map( A1 => n47, A2 => B(24), ZN => n52);
   U152 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n89, ZN => n88);
   U153 : OAI22_X1 port map( A1 => B(32), A2 => n139, B1 => A(32), B2 => n88, 
                           ZN => n79);
   U154 : XNOR2_X1 port map( A => n92, B => n139, ZN => SUM(32));
   U155 : NOR2_X1 port map( A1 => B(31), A2 => n74, ZN => n86);
   U156 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n89, ZN => n139);
   U157 : NOR2_X1 port map( A1 => n79, A2 => n78, ZN => carry_33_port);
   U158 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n70);
   U159 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n140);
   U160 : OAI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n142);
   U161 : NAND2_X1 port map( A1 => B(26), A2 => n55, ZN => n62);
   U162 : XNOR2_X1 port map( A => n98, B => n146, ZN => SUM(26));
   U163 : NOR2_X1 port map( A1 => B(30), A2 => n70, ZN => n143);
   U164 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => n144);
   U165 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n102);
   U166 : NAND2_X1 port map( A1 => A(22), A2 => B(22), ZN => n46);
   U167 : INV_X1 port map( A => A(22), ZN => n44);
   U168 : NOR2_X1 port map( A1 => B(28), A2 => n141, ZN => n145);
   U169 : BUF_X1 port map( A => n55, Z => n146);
   U170 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n128, ZN => n103);
   U171 : CLKBUF_X1 port map( A => n103, Z => n147);
   U172 : XNOR2_X1 port map( A => B(26), B => A(26), ZN => n98);
   U173 : INV_X1 port map( A => A(26), ZN => n61);
   U174 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n95);
   U175 : INV_X1 port map( A => A(29), ZN => n72);
   U176 : XNOR2_X1 port map( A => B(28), B => A(28), ZN => n96);
   U177 : INV_X1 port map( A => A(28), ZN => n68);
   U178 : XNOR2_X1 port map( A => B(27), B => A(27), ZN => n97);
   U179 : INV_X1 port map( A => A(27), ZN => n64);
   U180 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n94);
   U181 : INV_X1 port map( A => A(30), ZN => n76);
   U182 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n93);
   U183 : INV_X1 port map( A => A(31), ZN => n87);
   U184 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n92);
   U185 : NOR2_X1 port map( A1 => B(32), A2 => A(32), ZN => n78);
   U186 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n100);
   U187 : INV_X1 port map( A => A(24), ZN => n53);
   U188 : INV_X1 port map( A => A(21), ZN => n84);
   U189 : INV_X1 port map( A => n103, ZN => n43);
   U190 : XNOR2_X1 port map( A => B(25), B => A(25), ZN => n99);
   U191 : INV_X1 port map( A => A(25), ZN => n57);
   U192 : XNOR2_X1 port map( A => n95, B => n135, ZN => SUM(29));
   U193 : XNOR2_X1 port map( A => n96, B => n141, ZN => SUM(28));
   U194 : OAI21_X1 port map( B1 => B(34), B2 => A(34), A => carry_34_port, ZN 
                           => net67872);
   U195 : XNOR2_X1 port map( A => n148, B => net74815, ZN => SUM(34));
   U196 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n148);
   U197 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => net67871);
   U198 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => n149);
   U199 : NAND2_X1 port map( A1 => n2, A2 => n258, ZN => n150);
   U200 : NOR2_X1 port map( A1 => B(40), A2 => n6, ZN => n151);
   U201 : NOR2_X1 port map( A1 => n199, A2 => B(38), ZN => n152);
   U202 : OAI21_X1 port map( B1 => B(47), B2 => n232, A => A(47), ZN => n153);
   U203 : NAND2_X1 port map( A1 => n164, A2 => B(37), ZN => n154);
   U204 : INV_X1 port map( A => n234, ZN => n155);
   U205 : XNOR2_X1 port map( A => net68135, B => net67982, ZN => SUM(53));
   U206 : INV_X1 port map( A => A(53), ZN => net67982);
   U207 : OAI21_X1 port map( B1 => net67982, B2 => net68177, A => net67983, ZN 
                           => net68162);
   U208 : OAI21_X1 port map( B1 => net68177, B2 => net67982, A => net67983, ZN 
                           => net68161);
   U209 : OAI21_X1 port map( B1 => net67981, B2 => net67982, A => net67983, ZN 
                           => net67980);
   U210 : XNOR2_X1 port map( A => n157, B => net68103, ZN => net68135);
   U211 : OAI21_X1 port map( B1 => n156, B2 => net67975, A => net67977, ZN => 
                           n157);
   U212 : NOR2_X1 port map( A1 => n157, A2 => B(53), ZN => net67981);
   U213 : INV_X1 port map( A => A(52), ZN => n156);
   U214 : XNOR2_X1 port map( A => net68136, B => n156, ZN => SUM(52));
   U215 : NAND2_X1 port map( A1 => net67974, A2 => B(53), ZN => net67983);
   U216 : NOR2_X1 port map( A1 => net67974, A2 => B(53), ZN => net68177);
   U217 : NOR2_X1 port map( A1 => net67969, A2 => B(52), ZN => net67975);
   U218 : NAND2_X1 port map( A1 => n149, A2 => B(52), ZN => net67977);
   U219 : XNOR2_X1 port map( A => n149, B => n158, ZN => net68136);
   U220 : NOR2_X1 port map( A1 => n195, A2 => B(37), ZN => n159);
   U221 : XNOR2_X1 port map( A => n317, B => n197, ZN => SUM(36));
   U222 : NOR2_X1 port map( A1 => B(36), A2 => n191, ZN => n160);
   U223 : INV_X1 port map( A => n219, ZN => n161);
   U224 : OAI21_X1 port map( B1 => n217, B2 => B(43), A => A(43), ZN => n162);
   U225 : OAI21_X1 port map( B1 => n240, B2 => n241, A => n242, ZN => n163);
   U226 : OAI21_X1 port map( B1 => n196, B2 => n197, A => n198, ZN => n164);
   U227 : CLKBUF_X1 port map( A => A(39), Z => n165);
   U228 : NOR2_X1 port map( A1 => net67980, A2 => B(54), ZN => n166);
   U229 : OAI21_X1 port map( B1 => n233, B2 => n234, A => n235, ZN => n167);
   U230 : NOR2_X1 port map( A1 => n239, A2 => B(49), ZN => n168);
   U231 : XNOR2_X1 port map( A => n318, B => n193, ZN => SUM(35));
   U232 : INV_X1 port map( A => A(35), ZN => n193);
   U233 : CLKBUF_X1 port map( A => A(47), Z => n345);
   U234 : NAND2_X1 port map( A1 => n222, A2 => n223, ZN => n169);
   U235 : NOR2_X1 port map( A1 => n321, A2 => B(42), ZN => n170);
   U236 : NOR2_X1 port map( A1 => n209, A2 => B(41), ZN => n171);
   U237 : INV_X1 port map( A => A(44), ZN => n172);
   U238 : XNOR2_X1 port map( A => n313, B => n211, ZN => SUM(40));
   U239 : NOR2_X1 port map( A1 => B(56), A2 => n150, ZN => n173);
   U240 : XNOR2_X1 port map( A => n304, B => n245, ZN => SUM(49));
   U241 : NAND2_X1 port map( A1 => n153, A2 => n237, ZN => n174);
   U242 : NOR2_X1 port map( A1 => B(44), A2 => n221, ZN => n175);
   U243 : INV_X1 port map( A => A(45), ZN => n230);
   U244 : INV_X1 port map( A => A(40), ZN => n211);
   U245 : INV_X1 port map( A => A(42), ZN => n219);
   U246 : INV_X1 port map( A => A(37), ZN => n201);
   U247 : OAI21_X1 port map( B1 => n177, B2 => n176, A => n179, ZN => n180);
   U248 : XNOR2_X1 port map( A => n180, B => net68123, ZN => net68125);
   U249 : INV_X1 port map( A => A(62), ZN => n177);
   U250 : CLKBUF_X1 port map( A => n177, Z => n181);
   U251 : NOR2_X1 port map( A1 => B(62), A2 => net68160, ZN => n176);
   U252 : OAI21_X1 port map( B1 => n181, B2 => n176, A => n179, ZN => net68354)
                           ;
   U253 : NAND2_X1 port map( A1 => B(62), A2 => net68160, ZN => n179);
   U254 : XNOR2_X1 port map( A => n178, B => A(62), ZN => SUM(62));
   U255 : XNOR2_X1 port map( A => net68026, B => B(62), ZN => n178);
   U256 : XNOR2_X1 port map( A => net68125, B => net68363, ZN => SUM(63));
   U257 : NAND2_X1 port map( A1 => net68121, A2 => net68123, ZN => net68157);
   U258 : NAND2_X1 port map( A1 => B(63), A2 => net68398, ZN => net68033);
   U259 : INV_X1 port map( A => A(63), ZN => net68363);
   U260 : CLKBUF_X1 port map( A => A(63), Z => net68398);
   U261 : CLKBUF_X1 port map( A => A(54), Z => n182);
   U262 : NOR2_X1 port map( A1 => n323, A2 => B(58), ZN => n183);
   U263 : NOR2_X1 port map( A1 => n323, A2 => B(58), ZN => n269);
   U264 : OAI21_X1 port map( B1 => n188, B2 => n183, A => n271, ZN => n184);
   U265 : INV_X1 port map( A => A(61), ZN => n185);
   U266 : NAND2_X1 port map( A1 => B(56), A2 => n257, ZN => n263);
   U267 : BUF_X1 port map( A => A(60), Z => n341);
   U268 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => n186);
   U269 : BUF_X1 port map( A => A(59), Z => n187);
   U270 : XNOR2_X1 port map( A => n169, B => n287, ZN => n309);
   U271 : NAND2_X1 port map( A1 => B(44), A2 => n221, ZN => n227);
   U272 : NAND2_X1 port map( A1 => n222, A2 => n162, ZN => n221);
   U273 : INV_X1 port map( A => A(58), ZN => n188);
   U274 : OAI21_X1 port map( B1 => n279, B2 => n185, A => n280, ZN => net68160)
                           ;
   U275 : INV_X1 port map( A => A(57), ZN => n189);
   U276 : NAND2_X1 port map( A1 => B(48), A2 => n236, ZN => n242);
   U277 : NAND2_X1 port map( A1 => n335, A2 => B(49), ZN => n246);
   U278 : XNOR2_X1 port map( A => n305, B => n241, ZN => SUM(48));
   U279 : XNOR2_X1 port map( A => n6, B => n285, ZN => n313);
   U280 : NAND2_X1 port map( A1 => B(40), A2 => n206, ZN => n212);
   U281 : XNOR2_X1 port map( A => n294, B => n185, ZN => SUM(61));
   U282 : XNOR2_X1 port map( A => n215, B => n312, ZN => SUM(41));
   U283 : INV_X1 port map( A => net68398, ZN => net68121);
   U284 : NAND2_X1 port map( A1 => n258, A2 => n259, ZN => n257);
   U285 : XNOR2_X1 port map( A => n309, B => n226, ZN => SUM(44));
   U286 : XNOR2_X1 port map( A => n298, B => n189, ZN => SUM(57));
   U287 : INV_X1 port map( A => A(49), ZN => n245);
   U288 : XNOR2_X1 port map( A => n174, B => n289, ZN => n305);
   U289 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => n236);
   U290 : NAND2_X1 port map( A1 => n207, A2 => n208, ZN => n206);
   U291 : NOR2_X1 port map( A1 => B(61), A2 => n186, ZN => n279);
   U292 : OAI21_X1 port map( B1 => n185, B2 => n279, A => n280, ZN => net68026)
                           ;
   U293 : NOR2_X1 port map( A1 => B(45), A2 => n333, ZN => n229);
   U294 : OAI21_X1 port map( B1 => n230, B2 => n229, A => n231, ZN => n228);
   U295 : OAI21_X1 port map( B1 => n332, B2 => n230, A => n231, ZN => n319);
   U296 : OAI21_X1 port map( B1 => n332, B2 => n230, A => n231, ZN => n320);
   U297 : NAND2_X1 port map( A1 => n213, A2 => B(42), ZN => n220);
   U298 : XNOR2_X1 port map( A => n213, B => B(42), ZN => n311);
   U299 : NOR2_X1 port map( A1 => n321, A2 => B(42), ZN => n218);
   U300 : NOR2_X1 port map( A1 => B(41), A2 => n334, ZN => n214);
   U301 : OAI21_X1 port map( B1 => n214, B2 => n215, A => n216, ZN => n321);
   U302 : OAI21_X1 port map( B1 => n159, B2 => n201, A => n154, ZN => n199);
   U303 : NAND2_X1 port map( A1 => n322, A2 => B(38), ZN => n205);
   U304 : XNOR2_X1 port map( A => n322, B => B(38), ZN => n315);
   U305 : NOR2_X1 port map( A1 => n199, A2 => B(38), ZN => n203);
   U306 : NOR2_X1 port map( A1 => n195, A2 => B(37), ZN => n200);
   U307 : OAI21_X1 port map( B1 => n201, B2 => n200, A => n154, ZN => n322);
   U308 : OAI21_X1 port map( B1 => n266, B2 => n265, A => n267, ZN => n264);
   U309 : NAND2_X1 port map( A1 => B(58), A2 => n340, ZN => n271);
   U310 : XNOR2_X1 port map( A => n264, B => B(58), ZN => n297);
   U311 : NOR2_X1 port map( A1 => n260, A2 => B(57), ZN => n265);
   U312 : OAI21_X1 port map( B1 => n265, B2 => n266, A => n267, ZN => n323);
   U313 : OAI21_X1 port map( B1 => n183, B2 => n270, A => n271, ZN => n268);
   U314 : NAND2_X1 port map( A1 => n184, A2 => B(59), ZN => n275);
   U315 : XNOR2_X1 port map( A => n324, B => B(59), ZN => n296);
   U316 : NOR2_X1 port map( A1 => n268, A2 => B(59), ZN => n273);
   U317 : OAI21_X1 port map( B1 => n188, B2 => n269, A => n271, ZN => n324);
   U318 : OAI21_X1 port map( B1 => n168, B2 => n245, A => n246, ZN => n243);
   U319 : NAND2_X1 port map( A1 => n243, A2 => B(50), ZN => n250);
   U320 : XNOR2_X1 port map( A => B(50), B => n325, ZN => n303);
   U321 : NOR2_X1 port map( A1 => n243, A2 => B(50), ZN => n248);
   U322 : NOR2_X1 port map( A1 => B(49), A2 => n239, ZN => n244);
   U323 : OAI21_X1 port map( B1 => n245, B2 => n244, A => n246, ZN => n325);
   U324 : OAI21_X1 port map( B1 => n273, B2 => n274, A => n275, ZN => n272);
   U325 : NAND2_X1 port map( A1 => n272, A2 => B(60), ZN => n277);
   U326 : OAI21_X1 port map( B1 => n272, B2 => B(60), A => A(60), ZN => n278);
   U327 : XNOR2_X1 port map( A => n326, B => B(60), ZN => n295);
   U328 : OAI21_X1 port map( B1 => n274, B2 => n273, A => n275, ZN => n326);
   U329 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n247);
   U330 : NAND2_X1 port map( A1 => n247, A2 => B(51), ZN => n251);
   U331 : OAI21_X1 port map( B1 => n247, B2 => B(51), A => A(51), ZN => n252);
   U332 : XNOR2_X1 port map( A => n327, B => B(51), ZN => n302);
   U333 : OAI21_X1 port map( B1 => n249, B2 => n248, A => n250, ZN => n327);
   U334 : OAI21_X1 port map( B1 => n218, B2 => n219, A => n220, ZN => n217);
   U335 : NAND2_X1 port map( A1 => n328, A2 => B(43), ZN => n222);
   U336 : OAI21_X1 port map( B1 => n217, B2 => B(43), A => A(43), ZN => n223);
   U337 : XNOR2_X1 port map( A => n328, B => B(43), ZN => n310);
   U338 : OAI21_X1 port map( B1 => n170, B2 => n219, A => n220, ZN => n328);
   U339 : OAI21_X1 port map( B1 => n152, B2 => n204, A => n205, ZN => n202);
   U340 : NAND2_X1 port map( A1 => n329, A2 => B(39), ZN => n207);
   U341 : OAI21_X1 port map( B1 => n202, B2 => B(39), A => A(39), ZN => n208);
   U342 : XNOR2_X1 port map( A => n329, B => B(39), ZN => n314);
   U343 : OAI21_X1 port map( B1 => n204, B2 => n203, A => n205, ZN => n329);
   U344 : NOR2_X1 port map( A1 => B(54), A2 => net67980, ZN => n254);
   U345 : OAI21_X1 port map( B1 => n166, B2 => n255, A => n256, ZN => n253);
   U346 : NOR2_X1 port map( A1 => n228, A2 => B(46), ZN => n233);
   U347 : OAI21_X1 port map( B1 => n233, B2 => n234, A => n235, ZN => n232);
   U348 : OAI21_X1 port map( B1 => n343, B2 => n193, A => n194, ZN => n191);
   U349 : XNOR2_X1 port map( A => n331, B => n283, ZN => n317);
   U350 : NAND2_X1 port map( A1 => n331, A2 => B(36), ZN => n198);
   U351 : NOR2_X1 port map( A1 => n191, A2 => B(36), ZN => n196);
   U352 : NOR2_X1 port map( A1 => B(35), A2 => n347, ZN => n192);
   U353 : OAI21_X1 port map( B1 => n192, B2 => n193, A => n194, ZN => n331);
   U354 : NOR2_X1 port map( A1 => B(45), A2 => n333, ZN => n332);
   U355 : OAI21_X1 port map( B1 => n225, B2 => n172, A => n227, ZN => n224);
   U356 : XNOR2_X1 port map( A => n224, B => n288, ZN => n308);
   U357 : NAND2_X1 port map( A1 => n224, A2 => B(45), ZN => n231);
   U358 : NOR2_X1 port map( A1 => n169, A2 => B(44), ZN => n225);
   U359 : OAI21_X1 port map( B1 => n226, B2 => n175, A => n227, ZN => n333);
   U360 : XNOR2_X1 port map( A => n338, B => n297, ZN => SUM(58));
   U361 : NAND2_X1 port map( A1 => B(54), A2 => net68161, ZN => n256);
   U362 : INV_X1 port map( A => A(54), ZN => n255);
   U363 : XNOR2_X1 port map( A => n330, B => B(55), ZN => n300);
   U364 : NAND2_X1 port map( A1 => n330, A2 => B(55), ZN => n258);
   U365 : XNOR2_X1 port map( A => n296, B => n187, ZN => SUM(59));
   U366 : XNOR2_X1 port map( A => n295, B => n341, ZN => SUM(60));
   U367 : OAI21_X1 port map( B1 => n262, B2 => n261, A => n263, ZN => n260);
   U368 : XNOR2_X1 port map( A => n337, B => n292, ZN => n298);
   U369 : NAND2_X1 port map( A1 => n260, A2 => B(57), ZN => n267);
   U370 : XNOR2_X1 port map( A => B(54), B => net68162, ZN => n301);
   U371 : XNOR2_X1 port map( A => n300, B => n342, ZN => SUM(55));
   U372 : NOR2_X1 port map( A1 => B(56), A2 => n257, ZN => n261);
   U373 : OAI21_X1 port map( B1 => n151, B2 => n211, A => n212, ZN => n209);
   U374 : XNOR2_X1 port map( A => n334, B => n286, ZN => n312);
   U375 : NAND2_X1 port map( A1 => n209, A2 => B(41), ZN => n216);
   U376 : NOR2_X1 port map( A1 => B(40), A2 => n206, ZN => n210);
   U377 : OAI21_X1 port map( B1 => n210, B2 => n211, A => n212, ZN => n334);
   U378 : OAI21_X1 port map( B1 => n160, B2 => n197, A => n198, ZN => n195);
   U379 : XNOR2_X1 port map( A => n164, B => n284, ZN => n316);
   U380 : NAND2_X1 port map( A1 => n320, A2 => B(46), ZN => n235);
   U381 : INV_X1 port map( A => A(46), ZN => n234);
   U382 : XNOR2_X1 port map( A => n232, B => B(47), ZN => n306);
   U383 : NAND2_X1 port map( A1 => n167, A2 => B(47), ZN => n237);
   U384 : NOR2_X1 port map( A1 => B(48), A2 => n236, ZN => n240);
   U385 : OAI21_X1 port map( B1 => n336, B2 => n241, A => n242, ZN => n239);
   U386 : OAI21_X1 port map( B1 => n240, B2 => n241, A => n242, ZN => n335);
   U387 : NOR2_X1 port map( A1 => B(48), A2 => n174, ZN => n336);
   U388 : XNOR2_X1 port map( A => n316, B => n201, ZN => SUM(37));
   U389 : INV_X1 port map( A => A(56), ZN => n262);
   U390 : OAI21_X1 port map( B1 => n262, B2 => n173, A => n263, ZN => n337);
   U391 : XNOR2_X1 port map( A => n339, B => n302, ZN => SUM(51));
   U392 : XNOR2_X1 port map( A => B(46), B => n319, ZN => n307);
   U393 : INV_X1 port map( A => A(38), ZN => n204);
   U394 : OAI21_X1 port map( B1 => n167, B2 => B(47), A => A(47), ZN => n238);
   U395 : XNOR2_X1 port map( A => n306, B => n345, ZN => SUM(47));
   U396 : XNOR2_X1 port map( A => n303, B => n344, ZN => SUM(50));
   U397 : NAND2_X1 port map( A1 => net67872, A2 => net67871, ZN => n190);
   U398 : XNOR2_X1 port map( A => n161, B => n311, ZN => SUM(42));
   U399 : INV_X1 port map( A => A(36), ZN => n197);
   U400 : INV_X1 port map( A => A(58), ZN => n270);
   U401 : INV_X1 port map( A => n270, ZN => n338);
   U402 : CLKBUF_X1 port map( A => A(51), Z => n339);
   U403 : OAI21_X1 port map( B1 => B(55), B2 => n253, A => A(55), ZN => n259);
   U404 : XNOR2_X1 port map( A => n347, B => n282, ZN => n318);
   U405 : NAND2_X1 port map( A1 => n190, A2 => B(35), ZN => n194);
   U406 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => net67969);
   U407 : INV_X1 port map( A => A(57), ZN => n266);
   U408 : OAI21_X1 port map( B1 => n189, B2 => n265, A => n267, ZN => n340);
   U409 : INV_X1 port map( A => A(59), ZN => n274);
   U410 : INV_X1 port map( A => A(44), ZN => n226);
   U411 : CLKBUF_X1 port map( A => A(55), Z => n342);
   U412 : XNOR2_X1 port map( A => n301, B => n182, ZN => SUM(54));
   U413 : NAND2_X1 port map( A1 => net68157, A2 => net68354, ZN => n281);
   U414 : INV_X1 port map( A => A(41), ZN => n215);
   U415 : XNOR2_X1 port map( A => n155, B => n307, ZN => SUM(46));
   U416 : XNOR2_X1 port map( A => n310, B => n346, ZN => SUM(43));
   U417 : INV_X1 port map( A => A(48), ZN => n241);
   U418 : XNOR2_X1 port map( A => n1, B => n315, ZN => SUM(38));
   U419 : NOR2_X1 port map( A1 => B(35), A2 => n190, ZN => n343);
   U420 : XNOR2_X1 port map( A => n308, B => n230, ZN => SUM(45));
   U421 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => n276);
   U422 : XNOR2_X1 port map( A => n314, B => n165, ZN => SUM(39));
   U423 : XNOR2_X1 port map( A => n150, B => n291, ZN => n299);
   U424 : XNOR2_X1 port map( A => n262, B => n299, ZN => SUM(56));
   U425 : XNOR2_X1 port map( A => n276, B => n293, ZN => n294);
   U426 : NAND2_X1 port map( A1 => n186, A2 => B(61), ZN => n280);
   U427 : INV_X1 port map( A => A(50), ZN => n249);
   U428 : INV_X1 port map( A => n249, ZN => n344);
   U429 : XNOR2_X1 port map( A => n163, B => n290, ZN => n304);
   U430 : CLKBUF_X1 port map( A => A(43), Z => n346);
   U431 : NAND2_X1 port map( A1 => net67872, A2 => net67871, ZN => n347);
   U432 : XOR2_X1 port map( A => net84800, B => n5, Z => SUM(21));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_7_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_7_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_7_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_2_port, carry_1_port, net33448, net33446, net33437, net33429, 
      net33424, net33413, net33410, net33388, net33384, net33383, net33382, 
      net33380, net33379, net33376, net33375, net33373, net33370, net33363, 
      net33362, net33360, net33358, net33353, net33345, net33338, net33335, 
      net33331, net33307, net33263, net33252, net33250, net33246, net33245, 
      net33244, net33239, net33231, net33223, net33222, net33221, net33203, 
      net33240, net33238, net33364, net33237, net41434, net41427, net41426, 
      net41410, net41408, net41407, net41397, net41338, net41337, net41336, 
      net41324, net41315, net41314, net41313, net41306, net41304, net47234, 
      net51397, net41307, net41330, net61079, net33400, net33249, net63146, 
      net60938, net47233, net33262, net33255, net70463, net33359, carry_63_port
      , carry_62_port, net74683, net75019, net75434, net33377, net33324, 
      net33374, net33381, net68395, net33385, net33310, net33372, net33402, 
      net33205, net33204, net33199, net33197, net33403, net33130, net33128, 
      net33211, net33210, net33209, net33208, net33125, net33123, net33328, 
      net33188, net33186, net33171, net33169, net33398, net33200, net33198, 
      net33193, net33191, net33397, net33131, net33129, net33124, net33122, 
      net33399, net33147, net33145, net33180, net33412, net33396, net33395, 
      net33368, net33217, net33216, net33215, net33214, net33387, net33378, 
      net33165, net33164, net33163, net33162, net33408, net33119, net33118, 
      net33117, net33116, net33112, net33110, net70416, net33182, net33176, 
      net33174, net33450, net33304, net33113, net33154, net33152, net75571, 
      net75492, net33404, net33321, net33159, net33157, net33153, net33151, 
      net33438, net33194, net33192, net33187, net33416, net33317, net33148, 
      net33141, net33139, net33314, net33142, net33134, net33106, net33105, 
      net33104, net33423, net33177, net33170, net33168, net75032, net33136, 
      net33135, carry_32_port, carry_31_port, net41430, net41425, carry_30_port
      , carry_29_port, carry_28_port, carry_27_port, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174 : std_logic;

begin
   
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => carry_62_port, B => B(62), CI => A(62), CO => 
                           carry_63_port, S => SUM(62));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_27 : FA_X1 port map( A => carry_27_port, B => B(27), CI => A(27), CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1 : NOR2_X1 port map( A1 => net68395, A2 => B(35), ZN => n1);
   U2 : NAND2_X1 port map( A1 => n35, A2 => net33182, ZN => n2);
   U3 : NOR2_X1 port map( A1 => n124, A2 => B(22), ZN => n3);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n129, A => n130, ZN => n4);
   U5 : BUF_X1 port map( A => net33170, Z => n9);
   U6 : INV_X1 port map( A => A(47), ZN => n5);
   U7 : OAI21_X1 port map( B1 => n155, B2 => net33238, A => net33240, ZN => n6)
                           ;
   U8 : BUF_X1 port map( A => A(26), Z => net63146);
   U9 : OAI21_X1 port map( B1 => net33151, B2 => B(41), A => A(41), ZN => n7);
   U10 : INV_X1 port map( A => B(55), ZN => net33345);
   U11 : INV_X1 port map( A => B(47), ZN => net33331);
   U12 : NAND2_X1 port map( A1 => B(18), A2 => n119, ZN => net41306);
   U13 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n85);
   U14 : INV_X1 port map( A => A(8), ZN => n87);
   U15 : NAND2_X1 port map( A1 => B(8), A2 => n82, ZN => n88);
   U16 : NOR2_X1 port map( A1 => B(8), A2 => n82, ZN => n86);
   U17 : OAI21_X1 port map( B1 => n90, B2 => n91, A => n92, ZN => n89);
   U18 : INV_X1 port map( A => A(9), ZN => n91);
   U19 : NAND2_X1 port map( A1 => B(9), A2 => n85, ZN => n92);
   U20 : NOR2_X1 port map( A1 => B(9), A2 => n85, ZN => n90);
   U21 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n93);
   U22 : INV_X1 port map( A => A(10), ZN => n95);
   U23 : NAND2_X1 port map( A1 => B(10), A2 => n89, ZN => n96);
   U24 : NOR2_X1 port map( A1 => B(10), A2 => n89, ZN => n94);
   U25 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => n97);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => n93, ZN => n98);
   U27 : OAI21_X1 port map( B1 => B(11), B2 => n93, A => A(11), ZN => n99);
   U28 : OAI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n100);
   U29 : INV_X1 port map( A => A(12), ZN => n102);
   U30 : NAND2_X1 port map( A1 => B(12), A2 => n97, ZN => n103);
   U31 : NOR2_X1 port map( A1 => B(12), A2 => n97, ZN => n101);
   U32 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n104);
   U33 : INV_X1 port map( A => A(13), ZN => n106);
   U34 : NAND2_X1 port map( A1 => B(13), A2 => n100, ZN => n107);
   U35 : NOR2_X1 port map( A1 => B(13), A2 => n100, ZN => n105);
   U36 : OAI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n108);
   U37 : INV_X1 port map( A => A(14), ZN => n110);
   U38 : NAND2_X1 port map( A1 => B(14), A2 => n104, ZN => n111);
   U39 : NOR2_X1 port map( A1 => B(14), A2 => n104, ZN => n109);
   U40 : NAND2_X1 port map( A1 => n113, A2 => n114, ZN => n112);
   U41 : NAND2_X1 port map( A1 => B(15), A2 => n108, ZN => n113);
   U42 : OAI21_X1 port map( B1 => B(15), B2 => n108, A => A(15), ZN => n114);
   U43 : INV_X1 port map( A => A(16), ZN => n117);
   U44 : OAI21_X1 port map( B1 => n116, B2 => n117, A => n118, ZN => n115);
   U45 : NAND2_X1 port map( A1 => B(16), A2 => n112, ZN => n118);
   U46 : NOR2_X1 port map( A1 => B(16), A2 => n112, ZN => n116);
   U47 : INV_X1 port map( A => A(17), ZN => n121);
   U48 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => n119);
   U49 : NAND2_X1 port map( A1 => B(17), A2 => n115, ZN => n122);
   U50 : NOR2_X1 port map( A1 => B(17), A2 => n115, ZN => n120);
   U51 : INV_X1 port map( A => B(38), ZN => net33314);
   U52 : INV_X1 port map( A => B(39), ZN => net33317);
   U53 : INV_X1 port map( A => B(46), ZN => net33328);
   U54 : XNOR2_X1 port map( A => B(2), B => carry_2_port, ZN => n153);
   U55 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n141);
   U56 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n63);
   U57 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n64);
   U58 : OAI21_X1 port map( B1 => A(2), B2 => B(2), A => carry_2_port, ZN => 
                           n65);
   U59 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n140);
   U60 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => n66);
   U61 : INV_X1 port map( A => A(3), ZN => n68);
   U62 : NAND2_X1 port map( A1 => B(3), A2 => n63, ZN => n69);
   U63 : NOR2_X1 port map( A1 => B(3), A2 => n63, ZN => n67);
   U64 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n139);
   U65 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n70);
   U66 : INV_X1 port map( A => A(4), ZN => n72);
   U67 : NAND2_X1 port map( A1 => B(4), A2 => n66, ZN => n73);
   U68 : NOR2_X1 port map( A1 => B(4), A2 => n66, ZN => n71);
   U69 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n138);
   U70 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => n74);
   U71 : INV_X1 port map( A => A(5), ZN => n76);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n70, ZN => n77);
   U73 : NOR2_X1 port map( A1 => B(5), A2 => n70, ZN => n75);
   U74 : XNOR2_X1 port map( A => B(7), B => A(7), ZN => n137);
   U75 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U76 : INV_X1 port map( A => A(6), ZN => n80);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n74, ZN => n81);
   U78 : NOR2_X1 port map( A1 => B(6), A2 => n74, ZN => n79);
   U79 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => n82);
   U80 : NAND2_X1 port map( A1 => B(7), A2 => n78, ZN => n83);
   U81 : OAI21_X1 port map( B1 => B(7), B2 => n78, A => A(7), ZN => n84);
   U82 : XNOR2_X1 port map( A => n135, B => n85, ZN => SUM(9));
   U83 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n135);
   U84 : XNOR2_X1 port map( A => n152, B => n89, ZN => SUM(10));
   U85 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n152);
   U86 : XNOR2_X1 port map( A => n151, B => n93, ZN => SUM(11));
   U87 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n151);
   U88 : XNOR2_X1 port map( A => n150, B => n97, ZN => SUM(12));
   U89 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n150);
   U90 : XNOR2_X1 port map( A => n149, B => n100, ZN => SUM(13));
   U91 : XNOR2_X1 port map( A => B(13), B => A(13), ZN => n149);
   U92 : XNOR2_X1 port map( A => A(14), B => n148, ZN => SUM(14));
   U93 : XNOR2_X1 port map( A => B(14), B => n104, ZN => n148);
   U94 : XNOR2_X1 port map( A => A(15), B => n147, ZN => SUM(15));
   U95 : XNOR2_X1 port map( A => B(15), B => n108, ZN => n147);
   U96 : XNOR2_X1 port map( A => n146, B => n117, ZN => SUM(16));
   U97 : XNOR2_X1 port map( A => n112, B => n132, ZN => n146);
   U98 : INV_X1 port map( A => B(16), ZN => n132);
   U99 : XNOR2_X1 port map( A => n145, B => n121, ZN => SUM(17));
   U100 : XNOR2_X1 port map( A => n115, B => n133, ZN => n145);
   U101 : INV_X1 port map( A => B(17), ZN => n133);
   U102 : XNOR2_X1 port map( A => n144, B => n119, ZN => SUM(18));
   U103 : XNOR2_X1 port map( A => B(18), B => net41427, ZN => n144);
   U104 : INV_X1 port map( A => B(59), ZN => n47);
   U105 : XNOR2_X1 port map( A => A(2), B => n153, ZN => SUM(2));
   U106 : XNOR2_X1 port map( A => n141, B => n63, ZN => SUM(3));
   U107 : XNOR2_X1 port map( A => n140, B => n66, ZN => SUM(4));
   U108 : XNOR2_X1 port map( A => n139, B => n70, ZN => SUM(5));
   U109 : XNOR2_X1 port map( A => n138, B => n74, ZN => SUM(6));
   U110 : XNOR2_X1 port map( A => n137, B => n78, ZN => SUM(7));
   U111 : XNOR2_X1 port map( A => n136, B => n82, ZN => SUM(8));
   U112 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n136);
   U113 : OAI21_X1 port map( B1 => n37, B2 => n38, A => n39, ZN => 
                           carry_62_port);
   U114 : INV_X1 port map( A => B(54), ZN => n165);
   U115 : INV_X1 port map( A => A(33), ZN => n8);
   U116 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n10);
   U117 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n124);
   U118 : INV_X1 port map( A => B(43), ZN => net33324);
   U119 : INV_X1 port map( A => B(42), ZN => net33321);
   U120 : INV_X1 port map( A => B(50), ZN => net33335);
   U121 : INV_X1 port map( A => B(35), ZN => net33310);
   U122 : INV_X1 port map( A => B(25), ZN => n134);
   U123 : INV_X1 port map( A => B(34), ZN => net33307);
   U124 : INV_X1 port map( A => B(33), ZN => net33304);
   U125 : INV_X1 port map( A => B(51), ZN => net33338);
   U126 : BUF_X1 port map( A => n4, Z => net41434);
   U127 : OAI21_X1 port map( B1 => net33112, B2 => n33, A => n22, ZN => 
                           net51397);
   U128 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => 
                           carry_27_port);
   U129 : NAND2_X1 port map( A1 => net41430, A2 => B(26), ZN => n13);
   U130 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n12);
   U131 : NAND2_X1 port map( A1 => A(26), A2 => net41430, ZN => n11);
   U132 : OAI21_X1 port map( B1 => net41397, B2 => n14, A => net41426, ZN => 
                           net41430);
   U133 : INV_X1 port map( A => A(25), ZN => n14);
   U134 : XNOR2_X1 port map( A => net41408, B => n14, ZN => SUM(25));
   U135 : OAI21_X1 port map( B1 => net41397, B2 => n14, A => net41426, ZN => 
                           net41425);
   U136 : XNOR2_X1 port map( A => net41425, B => B(26), ZN => net41407);
   U137 : NAND2_X1 port map( A1 => n31, A2 => net33159, ZN => n15);
   U138 : INV_X1 port map( A => A(39), ZN => n16);
   U139 : NOR2_X1 port map( A1 => B(52), A2 => net33214, ZN => n17);
   U140 : CLKBUF_X1 port map( A => n123, Z => n18);
   U141 : NOR2_X1 port map( A1 => net33145, A2 => B(40), ZN => n19);
   U142 : NOR2_X1 port map( A1 => net33162, A2 => B(43), ZN => n20);
   U143 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => net41307);
   U144 : CLKBUF_X1 port map( A => n55, Z => n21);
   U145 : NAND2_X1 port map( A1 => net33104, A2 => B(33), ZN => n22);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => net41307, ZN => net41315);
   U147 : NOR2_X1 port map( A1 => net33180, A2 => B(46), ZN => n23);
   U148 : OAI21_X1 port map( B1 => A(32), B2 => B(32), A => carry_32_port, ZN 
                           => net33106);
   U149 : CLKBUF_X1 port map( A => carry_32_port, Z => net74683);
   U150 : NAND2_X1 port map( A1 => net33136, A2 => net33135, ZN => net75032);
   U151 : XNOR2_X1 port map( A => net75032, B => net33314, ZN => net33382);
   U152 : NAND2_X1 port map( A1 => net75032, A2 => B(38), ZN => net33142);
   U153 : OAI21_X1 port map( B1 => net33128, B2 => B(37), A => A(37), ZN => 
                           net33136);
   U154 : NAND2_X1 port map( A1 => net33136, A2 => net33135, ZN => net33134);
   U155 : NAND2_X1 port map( A1 => net33128, A2 => B(37), ZN => net33135);
   U156 : XNOR2_X1 port map( A => B(37), B => net33403, ZN => net33383);
   U157 : CLKBUF_X1 port map( A => A(37), Z => net33446);
   U158 : NAND2_X1 port map( A1 => net33423, A2 => B(44), ZN => net33177);
   U159 : OAI21_X1 port map( B1 => n24, B2 => net33176, A => net33177, ZN => 
                           net70416);
   U160 : OAI21_X1 port map( B1 => n25, B2 => net33176, A => net33177, ZN => 
                           net33174);
   U161 : OAI21_X1 port map( B1 => net33170, B2 => net33169, A => net33171, ZN 
                           => net33423);
   U162 : XNOR2_X1 port map( A => net33423, B => B(44), ZN => net33376);
   U163 : INV_X1 port map( A => A(43), ZN => net33170);
   U164 : XNOR2_X1 port map( A => net33377, B => n9, ZN => SUM(43));
   U165 : OAI21_X1 port map( B1 => n20, B2 => net33170, A => net33171, ZN => 
                           net33168);
   U166 : NOR2_X1 port map( A1 => net33168, A2 => B(44), ZN => n25);
   U167 : NOR2_X1 port map( A1 => B(44), A2 => net33168, ZN => n24);
   U168 : NAND2_X1 port map( A1 => net33106, A2 => net33105, ZN => net33104);
   U169 : XNOR2_X1 port map( A => net33104, B => net33304, ZN => net33387);
   U170 : NAND2_X1 port map( A1 => net33104, A2 => B(33), ZN => net33113);
   U171 : NAND2_X1 port map( A1 => A(32), A2 => B(32), ZN => net33105);
   U172 : NAND2_X1 port map( A1 => net33106, A2 => net33105, ZN => net33450);
   U173 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => net33388);
   U174 : OAI21_X1 port map( B1 => n27, B2 => net33141, A => net33142, ZN => 
                           net33139);
   U175 : OAI21_X1 port map( B1 => n26, B2 => net33141, A => net33142, ZN => 
                           net33416);
   U176 : NOR2_X1 port map( A1 => net33134, A2 => B(38), ZN => n26);
   U177 : NOR2_X1 port map( A1 => net33134, A2 => B(38), ZN => n27);
   U178 : NAND2_X1 port map( A1 => net33416, A2 => B(39), ZN => net33148);
   U179 : OAI21_X1 port map( B1 => net33147, B2 => n28, A => net33148, ZN => 
                           net33399);
   U180 : OAI21_X1 port map( B1 => n29, B2 => n16, A => net33148, ZN => 
                           net33145);
   U181 : XNOR2_X1 port map( A => net33416, B => net33317, ZN => net33381);
   U182 : INV_X1 port map( A => A(38), ZN => net33141);
   U183 : CLKBUF_X1 port map( A => net33141, Z => net75019);
   U184 : NOR2_X1 port map( A1 => net33139, A2 => B(39), ZN => n29);
   U185 : NOR2_X1 port map( A1 => net33139, A2 => B(39), ZN => n28);
   U186 : NAND2_X1 port map( A1 => net33438, A2 => B(47), ZN => net33194);
   U187 : OAI21_X1 port map( B1 => net33193, B2 => n30, A => net33194, ZN => 
                           net33398);
   U188 : OAI21_X1 port map( B1 => net33192, B2 => n5, A => net33194, ZN => 
                           net33191);
   U189 : OAI21_X1 port map( B1 => n23, B2 => net33187, A => net33188, ZN => 
                           net33438);
   U190 : NOR2_X1 port map( A1 => net33438, A2 => B(47), ZN => net33192);
   U191 : INV_X1 port map( A => A(46), ZN => net33187);
   U192 : XNOR2_X1 port map( A => net33374, B => net33187, ZN => SUM(46));
   U193 : OAI21_X1 port map( B1 => net33187, B2 => net33186, A => net33188, ZN 
                           => net33437);
   U194 : NOR2_X1 port map( A1 => B(47), A2 => net33437, ZN => n30);
   U195 : NOR2_X1 port map( A1 => B(42), A2 => net33157, ZN => net75492);
   U196 : OAI21_X1 port map( B1 => net75492, B2 => net33164, A => net33165, ZN 
                           => net33162);
   U197 : NOR2_X1 port map( A1 => n15, A2 => B(42), ZN => net33163);
   U198 : NAND2_X1 port map( A1 => net33157, A2 => B(42), ZN => net33165);
   U199 : NAND2_X1 port map( A1 => n31, A2 => n7, ZN => net33157);
   U200 : XNOR2_X1 port map( A => n15, B => net33321, ZN => net33378);
   U201 : OAI21_X1 port map( B1 => net33151, B2 => B(41), A => A(41), ZN => 
                           net33159);
   U202 : OAI21_X1 port map( B1 => n19, B2 => net33153, A => net33154, ZN => 
                           net33151);
   U203 : INV_X1 port map( A => A(40), ZN => net33153);
   U204 : OAI21_X1 port map( B1 => net33152, B2 => net33153, A => net33154, ZN 
                           => net33404);
   U205 : NAND2_X1 port map( A1 => net33404, A2 => B(41), ZN => n31);
   U206 : XNOR2_X1 port map( A => net33404, B => B(41), ZN => net33379);
   U207 : NOR2_X1 port map( A1 => B(50), A2 => net75571, ZN => n32);
   U208 : OAI21_X1 port map( B1 => n32, B2 => net33210, A => net33211, ZN => 
                           net33208);
   U209 : NAND2_X1 port map( A1 => net75571, A2 => B(50), ZN => net33211);
   U210 : NOR2_X1 port map( A1 => B(50), A2 => net33203, ZN => net33209);
   U211 : NAND2_X1 port map( A1 => net33205, A2 => net33204, ZN => net75571);
   U212 : NAND2_X1 port map( A1 => net33205, A2 => net33204, ZN => net33203);
   U213 : NOR2_X1 port map( A1 => B(40), A2 => net33145, ZN => net33152);
   U214 : NAND2_X1 port map( A1 => net33145, A2 => B(40), ZN => net33154);
   U215 : XNOR2_X1 port map( A => B(40), B => net33399, ZN => net33380);
   U216 : OAI21_X1 port map( B1 => n8, B2 => n33, A => n22, ZN => net33408);
   U217 : OAI21_X1 port map( B1 => n34, B2 => net33112, A => net33113, ZN => 
                           net33110);
   U218 : NOR2_X1 port map( A1 => net33450, A2 => B(33), ZN => n33);
   U219 : NOR2_X1 port map( A1 => B(33), A2 => net33450, ZN => n34);
   U220 : OAI21_X1 port map( B1 => net33174, B2 => B(45), A => A(45), ZN => 
                           net33182);
   U221 : INV_X1 port map( A => A(44), ZN => net33176);
   U222 : CLKBUF_X1 port map( A => A(44), Z => net33429);
   U223 : NAND2_X1 port map( A1 => n35, A2 => net33182, ZN => net33180);
   U224 : XNOR2_X1 port map( A => net70416, B => B(45), ZN => net33375);
   U225 : NAND2_X1 port map( A1 => net70416, A2 => B(45), ZN => n35);
   U226 : CLKBUF_X1 port map( A => A(45), Z => net33448);
   U227 : OAI21_X1 port map( B1 => net33117, B2 => net33118, A => net33119, ZN 
                           => net33116);
   U228 : NOR2_X1 port map( A1 => net68395, A2 => B(35), ZN => net33123);
   U229 : INV_X1 port map( A => A(34), ZN => net33118);
   U230 : OAI21_X1 port map( B1 => net33118, B2 => net33117, A => net33119, ZN 
                           => net68395);
   U231 : NOR2_X1 port map( A1 => net33110, A2 => B(34), ZN => net33117);
   U232 : INV_X1 port map( A => A(33), ZN => net33112);
   U233 : XNOR2_X1 port map( A => net33387, B => n8, ZN => SUM(33));
   U234 : NAND2_X1 port map( A1 => net33408, A2 => B(34), ZN => net33119);
   U235 : NOR2_X1 port map( A1 => net33162, A2 => B(43), ZN => net33169);
   U236 : INV_X1 port map( A => A(42), ZN => net33164);
   U237 : OAI21_X1 port map( B1 => net33163, B2 => net33164, A => net33165, ZN 
                           => net75434);
   U238 : XNOR2_X1 port map( A => net33378, B => net33164, ZN => SUM(42));
   U239 : XNOR2_X1 port map( A => net33368, B => A(52), ZN => SUM(52));
   U240 : XNOR2_X1 port map( A => net33396, B => B(52), ZN => net33368);
   U241 : OAI21_X1 port map( B1 => net33412, B2 => net33216, A => net33217, ZN 
                           => net33396);
   U242 : INV_X1 port map( A => A(51), ZN => net33216);
   U243 : OAI21_X1 port map( B1 => net33215, B2 => net33216, A => net33217, ZN 
                           => net33214);
   U244 : INV_X1 port map( A => A(52), ZN => net33222);
   U245 : NAND2_X1 port map( A1 => net33395, A2 => B(52), ZN => net33223);
   U246 : NOR2_X1 port map( A1 => B(52), A2 => net33214, ZN => net33221);
   U247 : NOR2_X1 port map( A1 => B(51), A2 => net33208, ZN => net33412);
   U248 : OAI21_X1 port map( B1 => net33216, B2 => net33412, A => net33217, ZN 
                           => net33395);
   U249 : NAND2_X1 port map( A1 => net33208, A2 => B(51), ZN => net33217);
   U250 : NOR2_X1 port map( A1 => B(51), A2 => net33413, ZN => net33215);
   U251 : NOR2_X1 port map( A1 => n2, A2 => B(46), ZN => net33186);
   U252 : XNOR2_X1 port map( A => n2, B => net33328, ZN => net33374);
   U253 : NAND2_X1 port map( A1 => B(46), A2 => net33180, ZN => net33188);
   U254 : INV_X1 port map( A => A(39), ZN => net33147);
   U255 : XNOR2_X1 port map( A => net33381, B => net33147, ZN => SUM(39));
   U256 : NOR2_X1 port map( A1 => net33122, A2 => B(36), ZN => net33129);
   U257 : OAI21_X1 port map( B1 => net33129, B2 => net33130, A => net33131, ZN 
                           => net33128);
   U258 : OAI21_X1 port map( B1 => net33130, B2 => net33129, A => net33131, ZN 
                           => net33403);
   U259 : OAI21_X1 port map( B1 => net33123, B2 => net33124, A => net33125, ZN 
                           => net33122);
   U260 : NAND2_X1 port map( A1 => net33122, A2 => B(36), ZN => net33131);
   U261 : INV_X1 port map( A => A(35), ZN => net33124);
   U262 : XNOR2_X1 port map( A => net33385, B => net33124, ZN => SUM(35));
   U263 : XNOR2_X1 port map( A => net33397, B => B(36), ZN => net33384);
   U264 : OAI21_X1 port map( B1 => net33124, B2 => n1, A => net33125, ZN => 
                           net33397);
   U265 : NOR2_X1 port map( A1 => net33191, A2 => B(48), ZN => net33198);
   U266 : OAI21_X1 port map( B1 => net33198, B2 => net33199, A => net33200, ZN 
                           => net33197);
   U267 : OAI21_X1 port map( B1 => net33199, B2 => net33198, A => net33200, ZN 
                           => net33402);
   U268 : NAND2_X1 port map( A1 => net33191, A2 => B(48), ZN => net33200);
   U269 : INV_X1 port map( A => A(47), ZN => net33193);
   U270 : XNOR2_X1 port map( A => net33373, B => net33193, ZN => SUM(47));
   U271 : XNOR2_X1 port map( A => net33398, B => B(48), ZN => net33372);
   U272 : NAND2_X1 port map( A1 => net75434, A2 => B(43), ZN => net33171);
   U273 : NAND2_X1 port map( A1 => net33116, A2 => B(35), ZN => net33125);
   U274 : INV_X1 port map( A => A(50), ZN => net33210);
   U275 : OAI21_X1 port map( B1 => net33209, B2 => net33210, A => net33211, ZN 
                           => net33413);
   U276 : XNOR2_X1 port map( A => net33370, B => net33210, ZN => SUM(50));
   U277 : INV_X1 port map( A => A(36), ZN => net33130);
   U278 : CLKBUF_X1 port map( A => A(36), Z => net47234);
   U279 : OAI21_X1 port map( B1 => net33197, B2 => B(49), A => A(49), ZN => 
                           net33205);
   U280 : NAND2_X1 port map( A1 => net33197, A2 => B(49), ZN => net33204);
   U281 : INV_X1 port map( A => A(48), ZN => net33199);
   U282 : XNOR2_X1 port map( A => net33402, B => B(49), ZN => n36);
   U283 : XNOR2_X1 port map( A => n36, B => A(49), ZN => SUM(49));
   U284 : XNOR2_X1 port map( A => net33372, B => A(48), ZN => SUM(48));
   U285 : XNOR2_X1 port map( A => net33116, B => net33310, ZN => net33385);
   U286 : XNOR2_X1 port map( A => net75434, B => net33324, ZN => net33377);
   U287 : XNOR2_X1 port map( A => n170, B => net33118, ZN => SUM(34));
   U288 : NAND2_X1 port map( A1 => B(61), A2 => n42, ZN => n39);
   U289 : NOR2_X1 port map( A1 => n42, A2 => B(61), ZN => n38);
   U290 : INV_X1 port map( A => A(61), ZN => n37);
   U291 : XNOR2_X1 port map( A => n41, B => B(61), ZN => net33359);
   U292 : OAI21_X1 port map( B1 => net33353, B2 => n40, A => net33358, ZN => 
                           n42);
   U293 : INV_X1 port map( A => A(60), ZN => n40);
   U294 : OAI21_X1 port map( B1 => n40, B2 => net33353, A => net33358, ZN => 
                           n41);
   U295 : XNOR2_X1 port map( A => net33359, B => A(61), ZN => SUM(61));
   U296 : BUF_X1 port map( A => A(60), Z => net70463);
   U297 : CLKBUF_X1 port map( A => A(57), Z => n44);
   U298 : XNOR2_X1 port map( A => net33360, B => net70463, ZN => SUM(60));
   U299 : AND2_X1 port map( A1 => n159, A2 => n43, ZN => n160);
   U300 : AND2_X1 port map( A1 => n158, A2 => n165, ZN => n43);
   U301 : CLKBUF_X1 port map( A => A(56), Z => n62);
   U302 : XNOR2_X1 port map( A => n48, B => net33262, ZN => SUM(59));
   U303 : XNOR2_X1 port map( A => net47233, B => n47, ZN => n48);
   U304 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => net47233);
   U305 : INV_X1 port map( A => A(59), ZN => net33262);
   U306 : OAI21_X1 port map( B1 => net33262, B2 => net60938, A => net33263, ZN 
                           => net33424);
   U307 : NOR2_X1 port map( A1 => B(59), A2 => net33255, ZN => net60938);
   U308 : NAND2_X1 port map( A1 => net33255, A2 => B(59), ZN => net33263);
   U309 : OAI21_X1 port map( B1 => B(58), B2 => net33249, A => A(58), ZN => n46
                           );
   U310 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => net33255);
   U311 : NAND2_X1 port map( A1 => net33249, A2 => B(58), ZN => n45);
   U312 : INV_X1 port map( A => A(59), ZN => net61079);
   U313 : XNOR2_X1 port map( A => net33400, B => B(58), ZN => net33362);
   U314 : NOR2_X1 port map( A1 => B(20), A2 => net41307, ZN => net41313);
   U315 : OAI21_X1 port map( B1 => net41313, B2 => net41314, A => net41315, ZN 
                           => n123);
   U316 : OAI21_X1 port map( B1 => net33250, B2 => n49, A => net33252, ZN => 
                           net33249);
   U317 : INV_X1 port map( A => A(57), ZN => n49);
   U318 : OAI21_X1 port map( B1 => n49, B2 => net33250, A => net33252, ZN => 
                           net33400);
   U319 : XNOR2_X1 port map( A => net33363, B => n44, ZN => SUM(57));
   U320 : CLKBUF_X1 port map( A => A(53), Z => n50);
   U321 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n51);
   U322 : XNOR2_X1 port map( A => n51, B => net41330, ZN => SUM(24));
   U323 : INV_X1 port map( A => A(24), ZN => net41337);
   U324 : NAND2_X1 port map( A1 => B(24), A2 => net41330, ZN => net41338);
   U325 : NOR2_X1 port map( A1 => B(24), A2 => net41330, ZN => net41336);
   U326 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => net41330);
   U327 : OAI21_X1 port map( B1 => net41324, B2 => B(23), A => A(23), ZN => n53
                           );
   U328 : NAND2_X1 port map( A1 => n4, A2 => B(23), ZN => n52);
   U329 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => net41410);
   U330 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n54);
   U331 : XNOR2_X1 port map( A => n54, B => net41307, ZN => SUM(20));
   U332 : INV_X1 port map( A => A(20), ZN => net41314);
   U333 : OAI21_X1 port map( B1 => B(19), B2 => n55, A => A(19), ZN => n58);
   U334 : OAI21_X1 port map( B1 => net41304, B2 => n56, A => net41306, ZN => 
                           n55);
   U335 : INV_X1 port map( A => A(18), ZN => n56);
   U336 : INV_X1 port map( A => n56, ZN => net41427);
   U337 : NAND2_X1 port map( A1 => B(19), A2 => n55, ZN => n57);
   U338 : XNOR2_X1 port map( A => B(19), B => n60, ZN => n59);
   U339 : CLKBUF_X1 port map( A => A(19), Z => n60);
   U340 : XNOR2_X1 port map( A => n59, B => n21, ZN => SUM(19));
   U341 : OAI21_X1 port map( B1 => net41337, B2 => net41336, A => net41338, ZN 
                           => n61);
   U342 : NOR2_X1 port map( A1 => B(25), A2 => n131, ZN => net41397);
   U343 : NAND2_X1 port map( A1 => n123, A2 => B(21), ZN => n127);
   U344 : XNOR2_X1 port map( A => n143, B => n18, ZN => SUM(21));
   U345 : NOR2_X1 port map( A1 => n123, A2 => B(21), ZN => n125);
   U346 : NAND2_X1 port map( A1 => n10, A2 => B(22), ZN => n130);
   U347 : XNOR2_X1 port map( A => n142, B => n10, ZN => SUM(22));
   U348 : NOR2_X1 port map( A1 => n124, A2 => B(22), ZN => n128);
   U349 : NOR2_X1 port map( A1 => B(18), A2 => n119, ZN => net41304);
   U350 : OAI21_X1 port map( B1 => n128, B2 => n129, A => n130, ZN => net41324)
                           ;
   U351 : XNOR2_X1 port map( A => net41410, B => net41434, ZN => SUM(23));
   U352 : XNOR2_X1 port map( A => net63146, B => net41407, ZN => SUM(26));
   U353 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n143);
   U354 : INV_X1 port map( A => A(21), ZN => n126);
   U355 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n142);
   U356 : INV_X1 port map( A => A(22), ZN => n129);
   U357 : OAI21_X1 port map( B1 => net41337, B2 => net41336, A => net41338, ZN 
                           => n131);
   U358 : XNOR2_X1 port map( A => n61, B => n134, ZN => net41408);
   U359 : NAND2_X1 port map( A1 => n61, A2 => B(25), ZN => net41426);
   U360 : XNOR2_X1 port map( A => n154, B => B(56), ZN => net33364);
   U361 : XNOR2_X1 port map( A => net33364, B => n62, ZN => SUM(56));
   U362 : OAI21_X1 port map( B1 => net33238, B2 => n155, A => net33240, ZN => 
                           n154);
   U363 : NOR2_X1 port map( A1 => B(56), A2 => net33237, ZN => net33244);
   U364 : INV_X1 port map( A => A(55), ZN => n155);
   U365 : NAND2_X1 port map( A1 => n6, A2 => B(56), ZN => net33246);
   U366 : NOR2_X1 port map( A1 => B(56), A2 => net33237, ZN => net33410);
   U367 : OAI21_X1 port map( B1 => net33239, B2 => net33238, A => net33240, ZN 
                           => net33237);
   U368 : INV_X1 port map( A => A(55), ZN => net33239);
   U369 : INV_X1 port map( A => A(56), ZN => net33245);
   U370 : NOR2_X1 port map( A1 => net33231, A2 => B(55), ZN => net33238);
   U371 : NAND2_X1 port map( A1 => net33231, A2 => B(55), ZN => net33240);
   U372 : XNOR2_X1 port map( A => n161, B => n167, ZN => SUM(54));
   U373 : XNOR2_X1 port map( A => net33382, B => net75019, ZN => SUM(38));
   U374 : XNOR2_X1 port map( A => n166, B => net33239, ZN => SUM(55));
   U375 : NOR2_X1 port map( A1 => net33424, A2 => B(60), ZN => net33353);
   U376 : OAI21_X1 port map( B1 => net33244, B2 => net33245, A => net33246, ZN 
                           => n163);
   U377 : OAI21_X1 port map( B1 => net33245, B2 => net33410, A => net33246, ZN 
                           => n171);
   U378 : OAI21_X1 port map( B1 => net33410, B2 => net33245, A => net33246, ZN 
                           => n172);
   U379 : NOR2_X1 port map( A1 => B(57), A2 => n163, ZN => net33250);
   U380 : OAI21_X1 port map( B1 => n17, B2 => net33222, A => net33223, ZN => 
                           n156);
   U381 : OAI21_X1 port map( B1 => net33222, B2 => net33221, A => net33223, ZN 
                           => n173);
   U382 : OAI21_X1 port map( B1 => n161, B2 => n160, A => n162, ZN => net33231)
                           ;
   U383 : XNOR2_X1 port map( A => n174, B => net33345, ZN => n166);
   U384 : OAI21_X1 port map( B1 => n161, B2 => n160, A => n162, ZN => n174);
   U385 : XNOR2_X1 port map( A => net51397, B => net33307, ZN => n170);
   U386 : XNOR2_X1 port map( A => net33413, B => net33338, ZN => n169);
   U387 : OAI21_X1 port map( B1 => net61079, B2 => net60938, A => net33263, ZN 
                           => n164);
   U388 : NAND2_X1 port map( A1 => B(60), A2 => net33424, ZN => net33358);
   U389 : XNOR2_X1 port map( A => n164, B => B(60), ZN => net33360);
   U390 : NAND2_X1 port map( A1 => B(57), A2 => n172, ZN => net33252);
   U391 : XNOR2_X1 port map( A => n173, B => B(53), ZN => n168);
   U392 : NAND2_X1 port map( A1 => n156, A2 => B(53), ZN => n158);
   U393 : XNOR2_X1 port map( A => n171, B => B(57), ZN => net33363);
   U394 : XNOR2_X1 port map( A => net33375, B => net33448, ZN => SUM(45));
   U395 : XNOR2_X1 port map( A => net33437, B => net33331, ZN => net33373);
   U396 : XNOR2_X1 port map( A => net33376, B => net33429, ZN => SUM(44));
   U397 : OAI21_X1 port map( B1 => n156, B2 => B(53), A => A(53), ZN => n159);
   U398 : XNOR2_X1 port map( A => n168, B => n50, ZN => SUM(53));
   U399 : XNOR2_X1 port map( A => net33383, B => net33446, ZN => SUM(37));
   U400 : XNOR2_X1 port map( A => net33362, B => A(58), ZN => SUM(58));
   U401 : XNOR2_X1 port map( A => net33380, B => A(40), ZN => SUM(40));
   U402 : XNOR2_X1 port map( A => net33388, B => net74683, ZN => SUM(32));
   U403 : INV_X1 port map( A => A(54), ZN => n161);
   U404 : XNOR2_X1 port map( A => net33384, B => net47234, ZN => SUM(36));
   U405 : NAND2_X1 port map( A1 => n159, A2 => n158, ZN => n157);
   U406 : XNOR2_X1 port map( A => net33379, B => A(41), ZN => SUM(41));
   U407 : XNOR2_X1 port map( A => n157, B => n165, ZN => n167);
   U408 : NAND2_X1 port map( A1 => n157, A2 => B(54), ZN => n162);
   U409 : XNOR2_X1 port map( A => net33203, B => net33335, ZN => net33370);
   U410 : XNOR2_X1 port map( A => n169, B => net33216, ZN => SUM(51));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_8_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_8_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_8_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, net29687, 
      net29686, net29677, net29673, net29670, net29669, net29650, net29648, 
      net29643, net29458, net29435, net29421, net29419, net29409, net29407, 
      net29406, net29402, net29396, net29395, net33514, net33532, net29432, 
      net29430, net29438, net29437, net29436, net33512, net29671, net29607, 
      net29429, net29649, net47239, net49490, net49495, net29408, net29403, 
      net29401, net29676, net29597, net29400, net55491, net29431, net29694, 
      net29418, net55500, net55499, net55492, net29426, net29425, carry_63_port
      , carry_62_port, carry_61_port, carry_60_port, carry_59_port, 
      carry_58_port, carry_57_port, carry_56_port, carry_55_port, carry_54_port
      , carry_53_port, carry_52_port, carry_51_port, carry_50_port, 
      carry_49_port, carry_48_port, net29444, net29442, net29447, net29693, 
      net29449, net29448, net29441, net75184, net29461, net29460, net29459, 
      net29706, net29667, net29614, net74662, net29668, net29611, net29455, 
      net29454, net29453, net29452, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1 : AND2_X1 port map( A1 => n111, A2 => n1, ZN => n113);
   U2 : AND2_X1 port map( A1 => n110, A2 => n2, ZN => n1);
   U3 : INV_X1 port map( A => B(45), ZN => n2);
   U4 : INV_X1 port map( A => n88, ZN => n3);
   U5 : INV_X1 port map( A => A(37), ZN => n4);
   U6 : NOR2_X1 port map( A1 => B(22), A2 => n55, ZN => n5);
   U7 : OAI21_X1 port map( B1 => net29643, B2 => n35, A => net29648, ZN => n6);
   U8 : OAI21_X1 port map( B1 => B(39), B2 => n149, A => A(39), ZN => n7);
   U9 : INV_X1 port map( A => B(24), ZN => net55500);
   U10 : INV_X1 port map( A => B(20), ZN => net29597);
   U11 : INV_X1 port map( A => B(25), ZN => net29607);
   U12 : INV_X1 port map( A => B(19), ZN => n42);
   U13 : INV_X1 port map( A => B(32), ZN => n117);
   U14 : INV_X1 port map( A => B(21), ZN => n116);
   U15 : NOR2_X1 port map( A1 => n77, A2 => B(36), ZN => n8);
   U16 : NOR2_X1 port map( A1 => net29435, A2 => B(26), ZN => n9);
   U17 : INV_X1 port map( A => B(37), ZN => n120);
   U18 : INV_X1 port map( A => B(29), ZN => net29614);
   U19 : INV_X1 port map( A => B(40), ZN => n121);
   U20 : INV_X1 port map( A => B(41), ZN => n122);
   U21 : INV_X1 port map( A => B(33), ZN => n118);
   U22 : INV_X1 port map( A => B(36), ZN => n119);
   U23 : INV_X1 port map( A => B(28), ZN => net29611);
   U24 : INV_X1 port map( A => B(45), ZN => n123);
   U25 : NAND2_X1 port map( A1 => B(45), A2 => n161, ZN => n115);
   U26 : OAI21_X1 port map( B1 => n88, B2 => n87, A => n89, ZN => n149);
   U27 : OAI21_X1 port map( B1 => net29460, B2 => net29459, A => net29461, ZN 
                           => net29686);
   U28 : OAI21_X1 port map( B1 => net29454, B2 => net29453, A => net29455, ZN 
                           => net29452);
   U29 : XNOR2_X1 port map( A => net29452, B => net29614, ZN => net29667);
   U30 : INV_X1 port map( A => A(28), ZN => net29454);
   U31 : XNOR2_X1 port map( A => net29454, B => net29668, ZN => SUM(28));
   U32 : NOR2_X1 port map( A1 => B(28), A2 => net29447, ZN => net29453);
   U33 : OAI21_X1 port map( B1 => net74662, B2 => net29453, A => net29455, ZN 
                           => net29706);
   U34 : NAND2_X1 port map( A1 => net29447, A2 => B(28), ZN => net29455);
   U35 : INV_X1 port map( A => A(28), ZN => net74662);
   U36 : XNOR2_X1 port map( A => net29447, B => net29611, ZN => net29668);
   U37 : XNOR2_X1 port map( A => net29667, B => net29460, ZN => SUM(29));
   U38 : NAND2_X1 port map( A1 => net29706, A2 => B(29), ZN => net29461);
   U39 : NOR2_X1 port map( A1 => net29706, A2 => B(29), ZN => net29459);
   U40 : NOR2_X1 port map( A1 => B(29), A2 => net29706, ZN => net75184);
   U41 : INV_X1 port map( A => A(29), ZN => net29460);
   U42 : OAI21_X1 port map( B1 => net75184, B2 => net29460, A => net29461, ZN 
                           => net29458);
   U43 : NAND2_X1 port map( A1 => n30, A2 => B(36), ZN => n10);
   U44 : CLKBUF_X1 port map( A => A(34), Z => n26);
   U45 : CLKBUF_X1 port map( A => carry_17_port, Z => n11);
   U46 : INV_X1 port map( A => A(41), ZN => n12);
   U47 : NOR2_X1 port map( A1 => n101, A2 => B(43), ZN => n13);
   U48 : OAI21_X1 port map( B1 => n8, B2 => n81, A => n10, ZN => n14);
   U49 : BUF_X1 port map( A => A(22), Z => net33532);
   U50 : AND2_X1 port map( A1 => n64, A2 => n15, ZN => n66);
   U51 : AND2_X1 port map( A1 => n63, A2 => n117, ZN => n15);
   U52 : INV_X1 port map( A => A(25), ZN => n16);
   U53 : NAND2_X1 port map( A1 => n7, A2 => n91, ZN => n17);
   U54 : OAI21_X1 port map( B1 => net29441, B2 => B(27), A => A(27), ZN => 
                           net29449);
   U55 : NAND2_X1 port map( A1 => net29449, A2 => net29448, ZN => net29447);
   U56 : OAI21_X1 port map( B1 => n18, B2 => net29442, A => net29444, ZN => 
                           net29441);
   U57 : NAND2_X1 port map( A1 => net29441, A2 => B(27), ZN => net29448);
   U58 : INV_X1 port map( A => A(26), ZN => n18);
   U59 : OAI21_X1 port map( B1 => n9, B2 => n18, A => net29444, ZN => net29693)
                           ;
   U60 : XNOR2_X1 port map( A => net29693, B => B(27), ZN => net29669);
   U61 : CLKBUF_X1 port map( A => A(27), Z => net49490);
   U62 : CLKBUF_X1 port map( A => A(26), Z => net47239);
   U63 : NOR2_X1 port map( A1 => net29687, A2 => B(26), ZN => net29442);
   U64 : NAND2_X1 port map( A1 => net29687, A2 => B(26), ZN => net29444);
   U65 : XNOR2_X1 port map( A => net29435, B => B(26), ZN => net29670);
   U66 : CLKBUF_X1 port map( A => A(30), Z => n19);
   U67 : NOR2_X1 port map( A1 => n109, A2 => B(45), ZN => n20);
   U68 : CLKBUF_X1 port map( A => A(39), Z => n21);
   U69 : INV_X1 port map( A => A(33), ZN => n22);
   U70 : BUF_X1 port map( A => A(35), Z => n25);
   U71 : NOR2_X1 port map( A1 => B(34), A2 => n69, ZN => n23);
   U72 : NOR2_X1 port map( A1 => n77, A2 => B(36), ZN => n24);
   U73 : NOR2_X1 port map( A1 => B(41), A2 => n93, ZN => n27);
   U74 : INV_X1 port map( A => n35, ZN => n28);
   U75 : NOR2_X1 port map( A1 => B(40), A2 => n90, ZN => n29);
   U76 : NAND2_X1 port map( A1 => n79, A2 => n78, ZN => n30);
   U77 : NOR2_X1 port map( A1 => n82, A2 => B(38), ZN => n31);
   U78 : NOR2_X1 port map( A1 => n82, A2 => B(38), ZN => n87);
   U79 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => carry_48_port
                           );
   U80 : NAND2_X1 port map( A1 => n6, A2 => B(47), ZN => n34);
   U81 : NOR2_X1 port map( A1 => n36, A2 => B(47), ZN => n33);
   U82 : INV_X1 port map( A => A(47), ZN => n32);
   U83 : OAI21_X1 port map( B1 => net29643, B2 => n35, A => net29648, ZN => n36
                           );
   U84 : INV_X1 port map( A => A(46), ZN => n35);
   U85 : XNOR2_X1 port map( A => n6, B => B(47), ZN => net29649);
   U86 : XNOR2_X1 port map( A => net29650, B => n28, ZN => SUM(46));
   U87 : NAND2_X1 port map( A1 => net29426, A2 => net29425, ZN => net55492);
   U88 : NAND2_X1 port map( A1 => net55492, A2 => B(24), ZN => net29432);
   U89 : XNOR2_X1 port map( A => net55492, B => net55500, ZN => net55499);
   U90 : OAI21_X1 port map( B1 => net29418, B2 => B(23), A => A(23), ZN => 
                           net29426);
   U91 : NAND2_X1 port map( A1 => net29418, A2 => B(23), ZN => net29425);
   U92 : AND2_X1 port map( A1 => net55500, A2 => net29425, ZN => net55491);
   U93 : XNOR2_X1 port map( A => net29694, B => B(23), ZN => net29673);
   U94 : XNOR2_X1 port map( A => net55499, B => net29431, ZN => SUM(24));
   U95 : OAI21_X1 port map( B1 => net29419, B2 => n37, A => net29421, ZN => 
                           net29418);
   U96 : INV_X1 port map( A => A(22), ZN => n37);
   U97 : OAI21_X1 port map( B1 => n5, B2 => n37, A => net29421, ZN => net29694)
                           ;
   U98 : INV_X1 port map( A => A(24), ZN => net29431);
   U99 : OAI21_X1 port map( B1 => net29431, B2 => net29430, A => net29432, ZN 
                           => net29429);
   U100 : INV_X1 port map( A => A(24), ZN => net33512);
   U101 : OAI21_X1 port map( B1 => net29401, B2 => n40, A => net29403, ZN => 
                           n38);
   U102 : OAI21_X1 port map( B1 => net33514, B2 => net29407, A => net29409, ZN 
                           => n39);
   U103 : AND2_X1 port map( A1 => net55491, A2 => net29426, ZN => net29430);
   U104 : XNOR2_X1 port map( A => n38, B => net29597, ZN => net29676);
   U105 : XNOR2_X1 port map( A => net29676, B => net33514, ZN => SUM(20));
   U106 : NAND2_X1 port map( A1 => n38, A2 => B(20), ZN => net29409);
   U107 : INV_X1 port map( A => A(19), ZN => n40);
   U108 : NOR2_X1 port map( A1 => B(20), A2 => net29400, ZN => net29407);
   U109 : NOR2_X1 port map( A1 => B(20), A2 => net29400, ZN => net49495);
   U110 : OAI21_X1 port map( B1 => net29402, B2 => net29401, A => net29403, ZN 
                           => net29400);
   U111 : INV_X1 port map( A => A(19), ZN => net29402);
   U112 : AND2_X1 port map( A1 => net29396, A2 => n43, ZN => net29401);
   U113 : AND2_X1 port map( A1 => net29395, A2 => n42, ZN => n43);
   U114 : NAND2_X1 port map( A1 => n41, A2 => B(19), ZN => net29403);
   U115 : NAND2_X1 port map( A1 => net29395, A2 => net29396, ZN => n41);
   U116 : XNOR2_X1 port map( A => n41, B => n42, ZN => net29677);
   U117 : INV_X1 port map( A => A(20), ZN => net29408);
   U118 : OAI21_X1 port map( B1 => net29408, B2 => net49495, A => net29409, ZN 
                           => net29406);
   U119 : INV_X1 port map( A => A(20), ZN => net33514);
   U120 : INV_X1 port map( A => A(45), ZN => n114);
   U121 : XNOR2_X1 port map( A => net29649, B => A(47), ZN => SUM(47));
   U122 : NOR2_X1 port map( A1 => net29406, A2 => B(21), ZN => n44);
   U123 : XNOR2_X1 port map( A => net29429, B => net29607, ZN => net29671);
   U124 : XNOR2_X1 port map( A => net29671, B => net29437, ZN => SUM(25));
   U125 : OAI21_X1 port map( B1 => net33512, B2 => net29430, A => net29432, ZN 
                           => n45);
   U126 : NAND2_X1 port map( A1 => n45, A2 => B(25), ZN => net29438);
   U127 : NOR2_X1 port map( A1 => n45, A2 => B(25), ZN => net29436);
   U128 : INV_X1 port map( A => A(25), ZN => net29437);
   U129 : OAI21_X1 port map( B1 => net29437, B2 => net29436, A => net29438, ZN 
                           => net29687);
   U130 : OAI21_X1 port map( B1 => n16, B2 => net29436, A => net29438, ZN => 
                           net29435);
   U131 : OAI21_X1 port map( B1 => n57, B2 => n56, A => n58, ZN => n46);
   U132 : INV_X1 port map( A => A(42), ZN => n103);
   U133 : CLKBUF_X1 port map( A => A(31), Z => n47);
   U134 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => n48);
   U135 : CLKBUF_X1 port map( A => A(18), Z => n49);
   U136 : INV_X1 port map( A => A(21), ZN => n50);
   U137 : OAI21_X1 port map( B1 => B(39), B2 => n149, A => A(39), ZN => n92);
   U138 : XNOR2_X1 port map( A => n133, B => n81, ZN => SUM(36));
   U139 : INV_X1 port map( A => A(33), ZN => n71);
   U140 : NAND2_X1 port map( A1 => n48, A2 => B(32), ZN => n68);
   U141 : INV_X1 port map( A => A(37), ZN => n84);
   U142 : XOR2_X1 port map( A => n11, B => B(17), Z => n51);
   U143 : XOR2_X1 port map( A => A(17), B => n51, Z => SUM(17));
   U144 : NAND2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => n52);
   U145 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n53);
   U146 : NAND2_X1 port map( A1 => carry_17_port, A2 => B(17), ZN => n54);
   U147 : NAND3_X1 port map( A1 => n52, A2 => n54, A3 => n53, ZN => 
                           carry_18_port);
   U148 : XNOR2_X1 port map( A => net29677, B => net29402, ZN => SUM(19));
   U149 : NOR2_X1 port map( A1 => n159, A2 => B(46), ZN => net29643);
   U150 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U151 : NOR2_X1 port map( A1 => B(42), A2 => n154, ZN => n102);
   U152 : OAI21_X1 port map( B1 => n153, B2 => n103, A => n104, ZN => n143);
   U153 : NOR2_X1 port map( A1 => n156, A2 => B(37), ZN => n83);
   U154 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U155 : OAI21_X1 port map( B1 => n155, B2 => n4, A => n85, ZN => n144);
   U156 : NOR2_X1 port map( A1 => n65, A2 => B(33), ZN => n70);
   U157 : OAI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n69);
   U158 : OAI21_X1 port map( B1 => n157, B2 => n71, A => n72, ZN => n145);
   U159 : OAI21_X1 port map( B1 => n157, B2 => n22, A => n72, ZN => n146);
   U160 : NAND2_X1 port map( A1 => net29686, A2 => B(30), ZN => n62);
   U161 : XNOR2_X1 port map( A => net29458, B => B(30), ZN => n139);
   U162 : NOR2_X1 port map( A1 => net29686, A2 => B(30), ZN => n60);
   U163 : OAI21_X1 port map( B1 => n56, B2 => n50, A => n58, ZN => n55);
   U164 : NAND2_X1 port map( A1 => n46, A2 => B(22), ZN => net29421);
   U165 : XNOR2_X1 port map( A => n147, B => B(22), ZN => n140);
   U166 : NOR2_X1 port map( A1 => B(22), A2 => n55, ZN => net29419);
   U167 : NOR2_X1 port map( A1 => net29406, A2 => B(21), ZN => n56);
   U168 : OAI21_X1 port map( B1 => n44, B2 => n50, A => n58, ZN => n147);
   U169 : OAI21_X1 port map( B1 => n13, B2 => n107, A => n108, ZN => n105);
   U170 : NOR2_X1 port map( A1 => n101, A2 => B(43), ZN => n106);
   U171 : OAI21_X1 port map( B1 => n106, B2 => n107, A => n108, ZN => n148);
   U172 : OAI21_X1 port map( B1 => n31, B2 => n88, A => n89, ZN => n86);
   U173 : OAI21_X1 port map( B1 => n75, B2 => n74, A => n76, ZN => n73);
   U174 : NOR2_X1 port map( A1 => n69, A2 => B(34), ZN => n74);
   U175 : OAI21_X1 port map( B1 => n75, B2 => n23, A => n76, ZN => n150);
   U176 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n59);
   U177 : NAND2_X1 port map( A1 => n59, A2 => B(31), ZN => n63);
   U178 : OAI21_X1 port map( B1 => n59, B2 => B(31), A => A(31), ZN => n64);
   U179 : XNOR2_X1 port map( A => n151, B => B(31), ZN => n138);
   U180 : OAI21_X1 port map( B1 => n61, B2 => n60, A => n62, ZN => n151);
   U181 : OAI21_X1 port map( B1 => n29, B2 => n95, A => n96, ZN => n93);
   U182 : XNOR2_X1 port map( A => n152, B => n122, ZN => n128);
   U183 : NAND2_X1 port map( A1 => n152, A2 => B(41), ZN => n100);
   U184 : NOR2_X1 port map( A1 => n93, A2 => B(41), ZN => n98);
   U185 : NOR2_X1 port map( A1 => n17, A2 => B(40), ZN => n94);
   U186 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n152);
   U187 : NOR2_X1 port map( A1 => B(42), A2 => n154, ZN => n153);
   U188 : OAI21_X1 port map( B1 => n99, B2 => n27, A => n100, ZN => n97);
   U189 : NAND2_X1 port map( A1 => B(42), A2 => n154, ZN => n104);
   U190 : XNOR2_X1 port map( A => n97, B => B(42), ZN => n127);
   U191 : OAI21_X1 port map( B1 => n98, B2 => n12, A => n100, ZN => n154);
   U192 : NOR2_X1 port map( A1 => n14, A2 => B(37), ZN => n155);
   U193 : OAI21_X1 port map( B1 => n8, B2 => n81, A => n10, ZN => n80);
   U194 : XNOR2_X1 port map( A => n156, B => n120, ZN => n132);
   U195 : NAND2_X1 port map( A1 => n80, A2 => B(37), ZN => n85);
   U196 : OAI21_X1 port map( B1 => n24, B2 => n81, A => n10, ZN => n156);
   U197 : NOR2_X1 port map( A1 => n158, A2 => B(33), ZN => n157);
   U198 : OAI21_X1 port map( B1 => n67, B2 => n66, A => n68, ZN => n65);
   U199 : XNOR2_X1 port map( A => n65, B => n118, ZN => n136);
   U200 : NAND2_X1 port map( A1 => n158, A2 => B(33), ZN => n72);
   U201 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n158);
   U202 : OAI21_X1 port map( B1 => n20, B2 => n114, A => n115, ZN => n112);
   U203 : OAI21_X1 port map( B1 => n114, B2 => n113, A => n115, ZN => n159);
   U204 : XNOR2_X1 port map( A => A(42), B => n127, ZN => SUM(42));
   U205 : XNOR2_X1 port map( A => n112, B => B(46), ZN => net29650);
   U206 : NAND2_X1 port map( A1 => n112, A2 => B(46), ZN => net29648);
   U207 : XNOR2_X1 port map( A => n160, B => n116, ZN => n141);
   U208 : NAND2_X1 port map( A1 => n39, A2 => B(21), ZN => n58);
   U209 : OAI21_X1 port map( B1 => net29407, B2 => net29408, A => net29409, ZN 
                           => n160);
   U210 : NAND2_X1 port map( A1 => n144, A2 => B(38), ZN => n89);
   U211 : XNOR2_X1 port map( A => n86, B => B(39), ZN => n130);
   U212 : NAND2_X1 port map( A1 => B(39), A2 => n163, ZN => n91);
   U213 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => net29395);
   U214 : OAI21_X1 port map( B1 => A(18), B2 => B(18), A => carry_18_port, ZN 
                           => net29396);
   U215 : XNOR2_X1 port map( A => n142, B => n49, ZN => SUM(18));
   U216 : XNOR2_X1 port map( A => n105, B => B(44), ZN => n125);
   U217 : NAND2_X1 port map( A1 => n148, A2 => B(44), ZN => n110);
   U218 : NAND2_X1 port map( A1 => B(34), A2 => n146, ZN => n76);
   U219 : INV_X1 port map( A => A(34), ZN => n75);
   U220 : XNOR2_X1 port map( A => B(35), B => n150, ZN => n134);
   U221 : NAND2_X1 port map( A1 => n73, A2 => B(35), ZN => n78);
   U222 : NAND2_X1 port map( A1 => n90, A2 => B(40), ZN => n96);
   U223 : INV_X1 port map( A => A(41), ZN => n99);
   U224 : XNOR2_X1 port map( A => n143, B => B(43), ZN => n126);
   U225 : XNOR2_X1 port map( A => n144, B => B(38), ZN => n131);
   U226 : XNOR2_X1 port map( A => n125, B => A(44), ZN => SUM(44));
   U227 : XNOR2_X1 port map( A => n130, B => n21, ZN => SUM(39));
   U228 : XNOR2_X1 port map( A => n47, B => n138, ZN => SUM(31));
   U229 : XNOR2_X1 port map( A => net29669, B => net49490, ZN => SUM(27));
   U230 : XNOR2_X1 port map( A => net29673, B => A(23), ZN => SUM(23));
   U231 : XNOR2_X1 port map( A => n145, B => B(34), ZN => n135);
   U232 : XNOR2_X1 port map( A => n139, B => n19, ZN => SUM(30));
   U233 : XNOR2_X1 port map( A => net29670, B => net47239, ZN => SUM(26));
   U234 : XNOR2_X1 port map( A => n140, B => net33532, ZN => SUM(22));
   U235 : XNOR2_X1 port map( A => carry_18_port, B => B(18), ZN => n142);
   U236 : OAI21_X1 port map( B1 => n73, B2 => B(35), A => A(35), ZN => n79);
   U237 : XNOR2_X1 port map( A => n134, B => n25, ZN => SUM(35));
   U238 : INV_X1 port map( A => A(43), ZN => n107);
   U239 : INV_X1 port map( A => A(38), ZN => n88);
   U240 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => n109);
   U241 : XNOR2_X1 port map( A => n109, B => n123, ZN => n124);
   U242 : XNOR2_X1 port map( A => n17, B => n121, ZN => n129);
   U243 : XNOR2_X1 port map( A => n129, B => n95, ZN => SUM(40));
   U244 : XNOR2_X1 port map( A => n126, B => A(43), ZN => SUM(43));
   U245 : INV_X1 port map( A => A(30), ZN => n61);
   U246 : INV_X1 port map( A => A(21), ZN => n57);
   U247 : INV_X1 port map( A => A(36), ZN => n81);
   U248 : INV_X1 port map( A => A(32), ZN => n67);
   U249 : XNOR2_X1 port map( A => n131, B => n3, ZN => SUM(38));
   U250 : XNOR2_X1 port map( A => n135, B => n26, ZN => SUM(34));
   U251 : XNOR2_X1 port map( A => n124, B => n114, ZN => SUM(45));
   U252 : NAND2_X1 port map( A1 => n79, A2 => n78, ZN => n77);
   U253 : XNOR2_X1 port map( A => n48, B => n117, ZN => n137);
   U254 : XNOR2_X1 port map( A => n137, B => n67, ZN => SUM(32));
   U255 : XNOR2_X1 port map( A => n30, B => n119, ZN => n133);
   U256 : OAI21_X1 port map( B1 => n105, B2 => B(44), A => A(44), ZN => n111);
   U257 : NAND2_X1 port map( A1 => n110, A2 => n162, ZN => n161);
   U258 : XNOR2_X1 port map( A => n132, B => n84, ZN => SUM(37));
   U259 : NAND2_X1 port map( A1 => n143, A2 => B(43), ZN => n108);
   U260 : OAI21_X1 port map( B1 => n148, B2 => B(44), A => A(44), ZN => n162);
   U261 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => n90);
   U262 : OAI21_X1 port map( B1 => n31, B2 => n88, A => n89, ZN => n163);
   U263 : XNOR2_X1 port map( A => n136, B => n22, ZN => SUM(33));
   U264 : XNOR2_X1 port map( A => n141, B => n57, ZN => SUM(21));
   U265 : XNOR2_X1 port map( A => n128, B => n99, ZN => SUM(41));
   U266 : INV_X1 port map( A => A(40), ZN => n95);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_9_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_9_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_9_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net37361, net37305, net37303, net37298, net37249, net37064, net37062,
      net37057, net37051, net37050, net37049, net54021, net54018, net53926, 
      carry_63_port, carry_62_port, carry_61_port, carry_60_port, carry_59_port
      , carry_58_port, carry_57_port, carry_56_port, net75169, net75432, 
      net37333, net54002, net53998, carry_26_port, carry_25_port, carry_24_port
      , carry_23_port, carry_22_port, carry_21_port, net75549, net37058, 
      net75195, net37063, net37331, net37252, net37055, n1, n2, n3, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311 : 
      std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_56 : FA_X1 port map( A => carry_56_port, B => B(56), CI => A(56), CO => 
                           carry_57_port, S => SUM(56));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_59 : FA_X1 port map( A => carry_59_port, B => B(59), CI => A(59), CO => 
                           carry_60_port, S => SUM(59));
   U1_60 : FA_X1 port map( A => B(60), B => A(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1 : INV_X1 port map( A => A(29), ZN => n1);
   U2 : CLKBUF_X1 port map( A => A(55), Z => n2);
   U3 : BUF_X1 port map( A => n166, Z => n3);
   U4 : BUF_X1 port map( A => net53926, Z => n14);
   U5 : CLKBUF_X1 port map( A => A(39), Z => n4);
   U6 : INV_X1 port map( A => n183, ZN => n5);
   U7 : AND2_X1 port map( A1 => n36, A2 => n39, ZN => n6);
   U8 : AND2_X1 port map( A1 => n36, A2 => n39, ZN => n174);
   U9 : NOR2_X1 port map( A1 => n221, A2 => B(46), ZN => n7);
   U10 : NAND2_X1 port map( A1 => B(16), A2 => n154, ZN => n97);
   U11 : NAND2_X1 port map( A1 => B(51), A2 => n289, ZN => n244);
   U12 : INV_X1 port map( A => A(15), ZN => n93);
   U13 : NOR2_X1 port map( A1 => B(15), A2 => n87, ZN => n92);
   U14 : NAND2_X1 port map( A1 => B(15), A2 => n156, ZN => n94);
   U15 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n144);
   U16 : INV_X1 port map( A => n123, ZN => n145);
   U17 : INV_X1 port map( A => n121, ZN => n147);
   U18 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n150);
   U19 : INV_X1 port map( A => A(6), ZN => n109);
   U20 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n67);
   U21 : NOR2_X1 port map( A1 => B(14), A2 => n84, ZN => n88);
   U22 : NAND2_X1 port map( A1 => B(14), A2 => n84, ZN => n90);
   U23 : INV_X1 port map( A => B(37), ZN => n255);
   U24 : INV_X1 port map( A => B(41), ZN => n257);
   U25 : XNOR2_X1 port map( A => B(0), B => CI, ZN => n136);
   U26 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n142);
   U27 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n126);
   U28 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => n127);
   U29 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n140);
   U30 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => CI, ZN => n139);
   U31 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n122);
   U32 : OAI221_X1 port map( B1 => n143, B2 => n102, C1 => n143, C2 => n101, A 
                           => n144, ZN => n123);
   U33 : INV_X1 port map( A => B(2), ZN => n101);
   U34 : INV_X1 port map( A => A(2), ZN => n102);
   U35 : INV_X1 port map( A => n125, ZN => n143);
   U36 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n120);
   U37 : OAI221_X1 port map( B1 => n145, B2 => n104, C1 => n145, C2 => n103, A 
                           => n146, ZN => n121);
   U38 : INV_X1 port map( A => B(3), ZN => n103);
   U39 : INV_X1 port map( A => A(3), ZN => n104);
   U40 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n146);
   U41 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n118);
   U42 : OAI221_X1 port map( B1 => n147, B2 => n106, C1 => n147, C2 => n105, A 
                           => n148, ZN => n119);
   U43 : INV_X1 port map( A => B(4), ZN => n105);
   U44 : INV_X1 port map( A => A(4), ZN => n106);
   U45 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n148);
   U46 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n116);
   U47 : OAI211_X1 port map( C1 => n149, C2 => n107, A => n138, B => n150, ZN 
                           => n117);
   U48 : INV_X1 port map( A => B(5), ZN => n107);
   U49 : INV_X1 port map( A => n119, ZN => n149);
   U50 : NAND2_X1 port map( A1 => A(5), A2 => n119, ZN => n138);
   U51 : INV_X1 port map( A => n152, ZN => n115);
   U52 : OAI222_X1 port map( A1 => n151, A2 => n108, B1 => n151, B2 => n109, C1
                           => n109, C2 => n108, ZN => n152);
   U53 : INV_X1 port map( A => B(6), ZN => n108);
   U54 : INV_X1 port map( A => n117, ZN => n151);
   U55 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n112);
   U56 : OAI211_X1 port map( C1 => n64, C2 => n65, A => n66, B => n67, ZN => 
                           n63);
   U57 : INV_X1 port map( A => B(8), ZN => n65);
   U58 : INV_X1 port map( A => n114, ZN => n64);
   U59 : NAND2_X1 port map( A1 => A(8), A2 => n114, ZN => n66);
   U60 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n135);
   U61 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n68);
   U62 : INV_X1 port map( A => A(9), ZN => n70);
   U63 : NAND2_X1 port map( A1 => B(9), A2 => n63, ZN => n71);
   U64 : NOR2_X1 port map( A1 => B(9), A2 => n63, ZN => n69);
   U65 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n134);
   U66 : OAI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n72);
   U67 : INV_X1 port map( A => A(10), ZN => n74);
   U68 : NAND2_X1 port map( A1 => B(10), A2 => n68, ZN => n75);
   U69 : NOR2_X1 port map( A1 => B(10), A2 => n68, ZN => n73);
   U70 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n133);
   U71 : OAI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n76);
   U72 : INV_X1 port map( A => A(11), ZN => n78);
   U73 : NAND2_X1 port map( A1 => B(11), A2 => n72, ZN => n79);
   U74 : NOR2_X1 port map( A1 => B(11), A2 => n72, ZN => n77);
   U75 : XNOR2_X1 port map( A => B(13), B => A(13), ZN => n132);
   U76 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n80);
   U77 : NAND2_X1 port map( A1 => B(12), A2 => n76, ZN => n83);
   U78 : INV_X1 port map( A => A(12), ZN => n82);
   U79 : NOR2_X1 port map( A1 => B(12), A2 => n76, ZN => n81);
   U80 : XNOR2_X1 port map( A => B(14), B => A(14), ZN => n131);
   U81 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => n84);
   U82 : NAND2_X1 port map( A1 => B(13), A2 => n80, ZN => n85);
   U83 : OAI21_X1 port map( B1 => B(13), B2 => n80, A => A(13), ZN => n86);
   U84 : XNOR2_X1 port map( A => B(15), B => A(15), ZN => n130);
   U85 : INV_X1 port map( A => B(45), ZN => n259);
   U86 : INV_X1 port map( A => B(48), ZN => n260);
   U87 : INV_X1 port map( A => B(49), ZN => n261);
   U88 : INV_X1 port map( A => B(53), ZN => n262);
   U89 : XNOR2_X1 port map( A => A(0), B => n136, ZN => SUM(0));
   U90 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n124);
   U91 : OAI211_X1 port map( C1 => n141, C2 => n100, A => n137, B => n142, ZN 
                           => n125);
   U92 : INV_X1 port map( A => n127, ZN => n141);
   U93 : INV_X1 port map( A => B(1), ZN => n100);
   U94 : NAND2_X1 port map( A1 => A(1), A2 => n127, ZN => n137);
   U95 : XNOR2_X1 port map( A => n126, B => n127, ZN => SUM(1));
   U96 : XNOR2_X1 port map( A => n122, B => n123, ZN => SUM(3));
   U97 : XNOR2_X1 port map( A => n120, B => n121, ZN => SUM(4));
   U98 : XNOR2_X1 port map( A => n118, B => n119, ZN => SUM(5));
   U99 : XNOR2_X1 port map( A => n116, B => n117, ZN => SUM(6));
   U100 : XNOR2_X1 port map( A => n115, B => n8, ZN => SUM(7));
   U101 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n113);
   U102 : OAI221_X1 port map( B1 => n115, B2 => n111, C1 => n115, C2 => n110, A
                           => n153, ZN => n114);
   U103 : INV_X1 port map( A => B(7), ZN => n110);
   U104 : INV_X1 port map( A => A(7), ZN => n111);
   U105 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n153);
   U106 : XNOR2_X1 port map( A => n112, B => n63, ZN => SUM(9));
   U107 : XNOR2_X1 port map( A => n135, B => n68, ZN => SUM(10));
   U108 : XNOR2_X1 port map( A => n134, B => n72, ZN => SUM(11));
   U109 : XNOR2_X1 port map( A => n133, B => n76, ZN => SUM(12));
   U110 : XNOR2_X1 port map( A => n132, B => n80, ZN => SUM(13));
   U111 : XNOR2_X1 port map( A => n131, B => n84, ZN => SUM(14));
   U112 : XNOR2_X1 port map( A => n130, B => n156, ZN => SUM(15));
   U113 : XNOR2_X1 port map( A => n124, B => n125, ZN => SUM(2));
   U114 : XNOR2_X1 port map( A => n113, B => n114, ZN => SUM(8));
   U115 : INV_X1 port map( A => B(32), ZN => n252);
   U116 : INV_X1 port map( A => B(40), ZN => n256);
   U117 : XOR2_X1 port map( A => B(7), B => A(7), Z => n8);
   U118 : INV_X1 port map( A => B(33), ZN => n253);
   U119 : INV_X1 port map( A => B(36), ZN => n254);
   U120 : INV_X1 port map( A => B(29), ZN => n251);
   U121 : INV_X1 port map( A => B(28), ZN => net37252);
   U122 : INV_X1 port map( A => B(27), ZN => net37249);
   U123 : INV_X1 port map( A => B(44), ZN => n258);
   U124 : OAI21_X1 port map( B1 => n204, B2 => n203, A => n205, ZN => n298);
   U125 : NAND2_X1 port map( A1 => n215, A2 => n216, ZN => n41);
   U126 : XNOR2_X1 port map( A => n9, B => net37252, ZN => net37331);
   U127 : XNOR2_X1 port map( A => net37331, B => net37063, ZN => SUM(28));
   U128 : OAI21_X1 port map( B1 => n10, B2 => net75549, A => net37058, ZN => n9
                           );
   U129 : NAND2_X1 port map( A1 => net37055, A2 => B(28), ZN => net37064);
   U130 : INV_X1 port map( A => A(27), ZN => n10);
   U131 : NOR2_X1 port map( A1 => net37055, A2 => B(28), ZN => net37062);
   U132 : NOR2_X1 port map( A1 => B(28), A2 => n9, ZN => net75195);
   U133 : OAI21_X1 port map( B1 => net37057, B2 => net75549, A => net37058, ZN 
                           => net37055);
   U134 : INV_X1 port map( A => A(27), ZN => net37057);
   U135 : INV_X1 port map( A => A(28), ZN => net37063);
   U136 : OAI21_X1 port map( B1 => net75195, B2 => net37063, A => net37064, ZN 
                           => net37361);
   U137 : INV_X1 port map( A => A(28), ZN => net75169);
   U138 : NOR2_X1 port map( A1 => B(27), A2 => net37049, ZN => net75549);
   U139 : NAND2_X1 port map( A1 => net37049, A2 => B(27), ZN => net37058);
   U140 : NOR2_X1 port map( A1 => B(16), A2 => n91, ZN => n11);
   U141 : OAI21_X1 port map( B1 => n6, B2 => n38, A => n176, ZN => n12);
   U142 : NOR2_X1 port map( A1 => B(36), A2 => n185, ZN => n13);
   U143 : NOR2_X1 port map( A1 => B(29), A2 => n29, ZN => n15);
   U144 : OAI21_X1 port map( B1 => n167, B2 => n168, A => n169, ZN => n16);
   U145 : NAND2_X1 port map( A1 => B(18), A2 => net53926, ZN => n21);
   U146 : NAND2_X1 port map( A1 => B(19), A2 => n26, ZN => net54002);
   U147 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => net53926);
   U148 : NOR2_X1 port map( A1 => n303, A2 => B(37), ZN => n17);
   U149 : XNOR2_X1 port map( A => B(17), B => A(17), ZN => n128);
   U150 : OAI21_X1 port map( B1 => B(17), B2 => n95, A => A(17), ZN => n99);
   U151 : XNOR2_X1 port map( A => carry_26_port, B => B(26), ZN => net37333);
   U152 : OAI21_X1 port map( B1 => A(26), B2 => B(26), A => carry_26_port, ZN 
                           => net37051);
   U153 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => carry_21_port);
   U154 : OAI22_X1 port map( A1 => B(20), A2 => n27, B1 => A(20), B2 => n27, ZN
                           => n23);
   U155 : INV_X1 port map( A => A(19), ZN => n24);
   U156 : OAI21_X1 port map( B1 => net53998, B2 => n24, A => net54002, ZN => 
                           n27);
   U157 : NOR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n22);
   U158 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => net54018);
   U159 : NOR2_X1 port map( A1 => B(19), A2 => n18, ZN => net53998);
   U160 : OAI21_X1 port map( B1 => n28, B2 => n20, A => n21, ZN => n18);
   U161 : INV_X1 port map( A => A(18), ZN => n20);
   U162 : OAI21_X1 port map( B1 => n19, B2 => n20, A => n21, ZN => n26);
   U163 : NOR2_X1 port map( A1 => B(18), A2 => net53926, ZN => n28);
   U164 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => net54021);
   U165 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n25);
   U166 : NOR2_X1 port map( A1 => B(18), A2 => net53926, ZN => n19);
   U167 : XNOR2_X1 port map( A => n25, B => n14, ZN => SUM(18));
   U168 : XNOR2_X1 port map( A => net37333, B => net75432, ZN => SUM(26));
   U169 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => net37050);
   U170 : CLKBUF_X1 port map( A => A(26), Z => net75432);
   U171 : OAI21_X1 port map( B1 => net75169, B2 => net37062, A => net37064, ZN 
                           => n29);
   U172 : NAND2_X1 port map( A1 => net37051, A2 => net37050, ZN => n30);
   U173 : CLKBUF_X1 port map( A => A(47), Z => n53);
   U174 : OAI21_X1 port map( B1 => n181, B2 => B(35), A => A(35), ZN => n31);
   U175 : AND2_X1 port map( A1 => n200, A2 => n40, ZN => n203);
   U176 : CLKBUF_X1 port map( A => n208, Z => n32);
   U177 : OAI21_X1 port map( B1 => B(47), B2 => n225, A => A(47), ZN => n33);
   U178 : OAI21_X1 port map( B1 => n174, B2 => n38, A => n176, ZN => n34);
   U179 : OAI21_X1 port map( B1 => n174, B2 => n175, A => n176, ZN => n304);
   U180 : NAND2_X1 port map( A1 => n186, A2 => n31, ZN => n35);
   U181 : OAI21_X1 port map( B1 => B(31), B2 => n3, A => A(31), ZN => n36);
   U182 : OAI21_X1 port map( B1 => n160, B2 => B(43), A => A(43), ZN => n37);
   U183 : OAI21_X1 port map( B1 => n203, B2 => n204, A => n205, ZN => n202);
   U184 : INV_X1 port map( A => A(32), ZN => n38);
   U185 : AND2_X1 port map( A1 => n171, A2 => n252, ZN => n39);
   U186 : AND2_X1 port map( A1 => n201, A2 => n256, ZN => n40);
   U187 : NAND2_X1 port map( A1 => n35, A2 => B(36), ZN => n191);
   U188 : NOR2_X1 port map( A1 => n291, A2 => B(38), ZN => n42);
   U189 : NOR2_X1 port map( A1 => B(41), A2 => n298, ZN => n43);
   U190 : OAI21_X1 port map( B1 => n44, B2 => n45, A => n46, ZN => 
                           carry_56_port);
   U191 : NAND2_X1 port map( A1 => n48, A2 => B(55), ZN => n46);
   U192 : NOR2_X1 port map( A1 => B(55), A2 => n50, ZN => n45);
   U193 : INV_X1 port map( A => A(55), ZN => n44);
   U194 : XNOR2_X1 port map( A => n48, B => B(55), ZN => n49);
   U195 : OAI21_X1 port map( B1 => net37298, B2 => n47, A => net37303, ZN => 
                           n50);
   U196 : INV_X1 port map( A => A(54), ZN => n47);
   U197 : OAI21_X1 port map( B1 => net37298, B2 => n47, A => net37303, ZN => 
                           n48);
   U198 : XNOR2_X1 port map( A => n2, B => n49, ZN => SUM(55));
   U199 : CLKBUF_X1 port map( A => A(31), Z => n51);
   U200 : INV_X1 port map( A => A(48), ZN => n52);
   U201 : CLKBUF_X1 port map( A => A(52), Z => n57);
   U202 : CLKBUF_X1 port map( A => A(51), Z => n54);
   U203 : CLKBUF_X1 port map( A => A(50), Z => n55);
   U204 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => n56);
   U205 : NOR2_X1 port map( A1 => n177, A2 => B(34), ZN => n58);
   U206 : NOR2_X1 port map( A1 => B(30), A2 => n162, ZN => n59);
   U207 : NOR2_X1 port map( A1 => n214, A2 => B(44), ZN => n60);
   U208 : NOR2_X1 port map( A1 => n173, A2 => B(33), ZN => n61);
   U209 : NAND2_X1 port map( A1 => n290, A2 => B(46), ZN => n228);
   U210 : XNOR2_X1 port map( A => n276, B => n204, ZN => SUM(40));
   U211 : INV_X1 port map( A => A(45), ZN => n223);
   U212 : XNOR2_X1 port map( A => A(54), B => net37305, ZN => SUM(54));
   U213 : NAND2_X1 port map( A1 => n215, A2 => n37, ZN => n214);
   U214 : XNOR2_X1 port map( A => n129, B => n154, ZN => SUM(16));
   U215 : XNOR2_X1 port map( A => n272, B => n219, ZN => SUM(44));
   U216 : XNOR2_X1 port map( A => n41, B => n258, ZN => n272);
   U217 : NAND2_X1 port map( A1 => n170, A2 => B(32), ZN => n176);
   U218 : XNOR2_X1 port map( A => n279, B => n194, ZN => SUM(37));
   U219 : OAI21_X1 port map( B1 => n307, B2 => n235, A => n236, ZN => n62);
   U220 : XNOR2_X1 port map( A => n287, B => n164, ZN => SUM(29));
   U221 : OAI21_X1 port map( B1 => n92, B2 => n93, A => n94, ZN => n91);
   U222 : OAI21_X1 port map( B1 => n92, B2 => n93, A => n94, ZN => n154);
   U223 : OAI21_X1 port map( B1 => n11, B2 => n96, A => n97, ZN => n95);
   U224 : OAI21_X1 port map( B1 => n11, B2 => n96, A => n97, ZN => n155);
   U225 : XNOR2_X1 port map( A => n128, B => n155, ZN => SUM(17));
   U226 : NAND2_X1 port map( A1 => B(17), A2 => n155, ZN => n98);
   U227 : XNOR2_X1 port map( A => net54018, B => n27, ZN => SUM(20));
   U228 : INV_X1 port map( A => A(14), ZN => n89);
   U229 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n87);
   U230 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n156);
   U231 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n129);
   U232 : INV_X1 port map( A => A(16), ZN => n96);
   U233 : XNOR2_X1 port map( A => net54021, B => n26, ZN => SUM(19));
   U234 : XNOR2_X1 port map( A => n283, B => n179, ZN => SUM(33));
   U235 : OAI21_X1 port map( B1 => n52, B2 => n306, A => n234, ZN => n157);
   U236 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => n158);
   U237 : XNOR2_X1 port map( A => n275, B => n32, ZN => SUM(41));
   U238 : INV_X1 port map( A => A(33), ZN => n179);
   U239 : XNOR2_X1 port map( A => n268, B => n52, ZN => SUM(48));
   U240 : XNOR2_X1 port map( A => n284, B => n38, ZN => SUM(32));
   U241 : INV_X1 port map( A => n168, ZN => n159);
   U242 : INV_X1 port map( A => A(53), ZN => n249);
   U243 : NAND2_X1 port map( A1 => n186, A2 => n187, ZN => n185);
   U244 : XNOR2_X1 port map( A => n35, B => n254, ZN => n280);
   U245 : XNOR2_X1 port map( A => n280, B => n190, ZN => SUM(36));
   U246 : XNOR2_X1 port map( A => n271, B => n223, ZN => SUM(45));
   U247 : OAI21_X1 port map( B1 => n211, B2 => n212, A => n213, ZN => n160);
   U248 : XNOR2_X1 port map( A => n229, B => n260, ZN => n268);
   U249 : XNOR2_X1 port map( A => n270, B => A(46), ZN => SUM(46));
   U250 : XNOR2_X1 port map( A => n249, B => n263, ZN => SUM(53));
   U251 : XNOR2_X1 port map( A => n56, B => n262, ZN => n263);
   U252 : NOR2_X1 port map( A1 => n308, A2 => B(54), ZN => net37298);
   U253 : NOR2_X1 port map( A1 => B(50), A2 => n300, ZN => n238);
   U254 : OAI21_X1 port map( B1 => n238, B2 => n239, A => n240, ZN => n237);
   U255 : OAI21_X1 port map( B1 => n299, B2 => n239, A => n240, ZN => n289);
   U256 : NOR2_X1 port map( A1 => n302, A2 => B(45), ZN => n222);
   U257 : OAI21_X1 port map( B1 => n222, B2 => n223, A => n224, ZN => n221);
   U258 : OAI21_X1 port map( B1 => n301, B2 => n223, A => n224, ZN => n290);
   U259 : NAND2_X1 port map( A1 => n206, A2 => B(42), ZN => n213);
   U260 : XNOR2_X1 port map( A => B(42), B => n305, ZN => n274);
   U261 : NOR2_X1 port map( A1 => n206, A2 => B(42), ZN => n211);
   U262 : OAI21_X1 port map( B1 => n17, B2 => n194, A => n195, ZN => n192);
   U263 : NAND2_X1 port map( A1 => n192, A2 => B(38), ZN => n199);
   U264 : XNOR2_X1 port map( A => n291, B => B(38), ZN => n278);
   U265 : NOR2_X1 port map( A1 => B(38), A2 => n192, ZN => n197);
   U266 : NOR2_X1 port map( A1 => n188, A2 => B(37), ZN => n193);
   U267 : OAI21_X1 port map( B1 => n193, B2 => n194, A => n195, ZN => n291);
   U268 : OAI21_X1 port map( B1 => n61, B2 => n179, A => n180, ZN => n177);
   U269 : NAND2_X1 port map( A1 => n292, A2 => B(34), ZN => n184);
   U270 : XNOR2_X1 port map( A => n292, B => B(34), ZN => n282);
   U271 : NOR2_X1 port map( A1 => n177, A2 => B(34), ZN => n182);
   U272 : NOR2_X1 port map( A1 => n34, A2 => B(33), ZN => n178);
   U273 : OAI21_X1 port map( B1 => n178, B2 => n179, A => n180, ZN => n292);
   U274 : OAI21_X1 port map( B1 => n1, B2 => n163, A => n165, ZN => n162);
   U275 : NAND2_X1 port map( A1 => n162, A2 => B(30), ZN => n169);
   U276 : XNOR2_X1 port map( A => n311, B => B(30), ZN => n286);
   U277 : NOR2_X1 port map( A1 => n162, A2 => B(30), ZN => n167);
   U278 : NOR2_X1 port map( A1 => n161, A2 => B(29), ZN => n163);
   U279 : NOR2_X1 port map( A1 => B(51), A2 => n237, ZN => n242);
   U280 : OAI21_X1 port map( B1 => n242, B2 => n243, A => n244, ZN => n241);
   U281 : OAI21_X1 port map( B1 => n242, B2 => n243, A => n244, ZN => n293);
   U282 : OAI21_X1 port map( B1 => n7, B2 => n227, A => n228, ZN => n225);
   U283 : NOR2_X1 port map( A1 => n221, A2 => B(46), ZN => n226);
   U284 : OAI21_X1 port map( B1 => n227, B2 => n226, A => n228, ZN => n294);
   U285 : OAI21_X1 port map( B1 => n211, B2 => n212, A => n213, ZN => n210);
   U286 : NAND2_X1 port map( A1 => n210, A2 => B(43), ZN => n215);
   U287 : OAI21_X1 port map( B1 => n160, B2 => B(43), A => A(43), ZN => n216);
   U288 : XNOR2_X1 port map( A => n210, B => B(43), ZN => n273);
   U289 : OAI21_X1 port map( B1 => n42, B2 => n198, A => n199, ZN => n196);
   U290 : NAND2_X1 port map( A1 => n295, A2 => B(39), ZN => n200);
   U291 : OAI21_X1 port map( B1 => n196, B2 => B(39), A => A(39), ZN => n201);
   U292 : XNOR2_X1 port map( A => n295, B => B(39), ZN => n277);
   U293 : OAI21_X1 port map( B1 => n197, B2 => n198, A => n199, ZN => n295);
   U294 : OAI21_X1 port map( B1 => n182, B2 => n183, A => n184, ZN => n181);
   U295 : NAND2_X1 port map( A1 => n296, A2 => B(35), ZN => n186);
   U296 : OAI21_X1 port map( B1 => n181, B2 => B(35), A => A(35), ZN => n187);
   U297 : XNOR2_X1 port map( A => n296, B => B(35), ZN => n281);
   U298 : OAI21_X1 port map( B1 => n58, B2 => n183, A => n184, ZN => n296);
   U299 : OAI21_X1 port map( B1 => n59, B2 => n168, A => n169, ZN => n166);
   U300 : NAND2_X1 port map( A1 => n297, A2 => B(31), ZN => n171);
   U301 : OAI21_X1 port map( B1 => n166, B2 => B(31), A => A(31), ZN => n172);
   U302 : XNOR2_X1 port map( A => n16, B => B(31), ZN => n285);
   U303 : OAI21_X1 port map( B1 => n167, B2 => n168, A => n169, ZN => n297);
   U304 : OAI21_X1 port map( B1 => n233, B2 => n52, A => n234, ZN => n232);
   U305 : XNOR2_X1 port map( A => n157, B => n261, ZN => n267);
   U306 : NAND2_X1 port map( A1 => n157, A2 => B(49), ZN => n236);
   U307 : NOR2_X1 port map( A1 => B(48), A2 => n229, ZN => n233);
   U308 : XNOR2_X1 port map( A => n298, B => n257, ZN => n275);
   U309 : NAND2_X1 port map( A1 => n202, A2 => B(41), ZN => n209);
   U310 : NOR2_X1 port map( A1 => n202, A2 => B(41), ZN => n207);
   U311 : NOR2_X1 port map( A1 => n62, A2 => B(50), ZN => n299);
   U312 : NAND2_X1 port map( A1 => n300, A2 => B(50), ZN => n240);
   U313 : XNOR2_X1 port map( A => n62, B => B(50), ZN => n266);
   U314 : OAI21_X1 port map( B1 => n307, B2 => n235, A => n236, ZN => n300);
   U315 : NOR2_X1 port map( A1 => n217, A2 => B(45), ZN => n301);
   U316 : OAI21_X1 port map( B1 => n60, B2 => n219, A => n220, ZN => n217);
   U317 : XNOR2_X1 port map( A => n302, B => n259, ZN => n271);
   U318 : NAND2_X1 port map( A1 => n217, A2 => B(45), ZN => n224);
   U319 : NOR2_X1 port map( A1 => n214, A2 => B(44), ZN => n218);
   U320 : OAI21_X1 port map( B1 => n218, B2 => n219, A => n220, ZN => n302);
   U321 : XNOR2_X1 port map( A => n266, B => n55, ZN => SUM(50));
   U322 : OAI21_X1 port map( B1 => n249, B2 => n248, A => n250, ZN => n247);
   U323 : NAND2_X1 port map( A1 => n308, A2 => B(54), ZN => net37303);
   U324 : XNOR2_X1 port map( A => n247, B => B(54), ZN => net37305);
   U325 : OAI21_X1 port map( B1 => n13, B2 => n190, A => n191, ZN => n188);
   U326 : XNOR2_X1 port map( A => n188, B => n255, ZN => n279);
   U327 : NAND2_X1 port map( A1 => n303, A2 => B(37), ZN => n195);
   U328 : NOR2_X1 port map( A1 => B(36), A2 => n185, ZN => n189);
   U329 : OAI21_X1 port map( B1 => n189, B2 => n190, A => n191, ZN => n303);
   U330 : OAI21_X1 port map( B1 => n6, B2 => n175, A => n176, ZN => n173);
   U331 : XNOR2_X1 port map( A => n12, B => n253, ZN => n283);
   U332 : NAND2_X1 port map( A1 => n304, A2 => B(33), ZN => n180);
   U333 : OAI21_X1 port map( B1 => net75169, B2 => net37062, A => net37064, ZN 
                           => n161);
   U334 : XNOR2_X1 port map( A => net37361, B => n251, ZN => n287);
   U335 : NAND2_X1 port map( A1 => n29, A2 => B(29), ZN => n165);
   U336 : XNOR2_X1 port map( A => n241, B => B(52), ZN => n264);
   U337 : NAND2_X1 port map( A1 => B(52), A2 => n293, ZN => n245);
   U338 : XNOR2_X1 port map( A => n273, B => A(43), ZN => SUM(43));
   U339 : NAND2_X1 port map( A1 => n41, A2 => B(44), ZN => n220);
   U340 : XNOR2_X1 port map( A => n158, B => n256, ZN => n276);
   U341 : NAND2_X1 port map( A1 => B(40), A2 => n158, ZN => n205);
   U342 : XNOR2_X1 port map( A => n309, B => n274, ZN => SUM(42));
   U343 : INV_X1 port map( A => A(42), ZN => n212);
   U344 : XNOR2_X1 port map( A => n294, B => B(47), ZN => n269);
   U345 : NAND2_X1 port map( A1 => n294, A2 => B(47), ZN => n230);
   U346 : NOR2_X1 port map( A1 => n56, A2 => B(53), ZN => n248);
   U347 : OAI21_X1 port map( B1 => n207, B2 => n208, A => n209, ZN => n206);
   U348 : OAI21_X1 port map( B1 => n43, B2 => n208, A => n209, ZN => n305);
   U349 : NOR2_X1 port map( A1 => B(48), A2 => n310, ZN => n306);
   U350 : NOR2_X1 port map( A1 => B(49), A2 => n232, ZN => n307);
   U351 : NAND2_X1 port map( A1 => B(48), A2 => n310, ZN => n234);
   U352 : NAND2_X1 port map( A1 => B(53), A2 => n56, ZN => n250);
   U353 : INV_X1 port map( A => A(49), ZN => n235);
   U354 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n308);
   U355 : XNOR2_X1 port map( A => n285, B => n51, ZN => SUM(31));
   U356 : INV_X1 port map( A => A(50), ZN => n239);
   U357 : XNOR2_X1 port map( A => n264, B => n57, ZN => SUM(52));
   U358 : XNOR2_X1 port map( A => n4, B => n277, ZN => SUM(39));
   U359 : INV_X1 port map( A => A(41), ZN => n208);
   U360 : NAND2_X1 port map( A1 => net37051, A2 => net37050, ZN => net37049);
   U361 : OAI21_X1 port map( B1 => n225, B2 => B(47), A => A(47), ZN => n231);
   U362 : XNOR2_X1 port map( A => n53, B => n269, ZN => SUM(47));
   U363 : XNOR2_X1 port map( A => n286, B => n159, ZN => SUM(30));
   U364 : XNOR2_X1 port map( A => n30, B => net37249, ZN => n288);
   U365 : XNOR2_X1 port map( A => A(38), B => n278, ZN => SUM(38));
   U366 : XNOR2_X1 port map( A => n290, B => B(46), ZN => n270);
   U367 : XNOR2_X1 port map( A => n289, B => B(51), ZN => n265);
   U368 : XNOR2_X1 port map( A => n281, B => A(35), ZN => SUM(35));
   U369 : OAI21_X1 port map( B1 => B(52), B2 => n293, A => A(52), ZN => n246);
   U370 : INV_X1 port map( A => A(32), ZN => n175);
   U371 : INV_X1 port map( A => A(40), ZN => n204);
   U372 : NAND2_X1 port map( A1 => n230, A2 => n231, ZN => n229);
   U373 : XNOR2_X1 port map( A => n5, B => n282, ZN => SUM(34));
   U374 : INV_X1 port map( A => A(30), ZN => n168);
   U375 : INV_X1 port map( A => A(46), ZN => n227);
   U376 : INV_X1 port map( A => A(51), ZN => n243);
   U377 : XNOR2_X1 port map( A => n267, B => n235, ZN => SUM(49));
   U378 : INV_X1 port map( A => n212, ZN => n309);
   U379 : NAND2_X1 port map( A1 => n33, A2 => n230, ZN => n310);
   U380 : INV_X1 port map( A => A(29), ZN => n164);
   U381 : OAI21_X1 port map( B1 => n15, B2 => n164, A => n165, ZN => n311);
   U382 : INV_X1 port map( A => A(38), ZN => n198);
   U383 : INV_X1 port map( A => A(37), ZN => n194);
   U384 : INV_X1 port map( A => A(44), ZN => n219);
   U385 : INV_X1 port map( A => A(36), ZN => n190);
   U386 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => n170);
   U387 : XNOR2_X1 port map( A => n170, B => n252, ZN => n284);
   U388 : XNOR2_X1 port map( A => n288, B => net37057, ZN => SUM(27));
   U389 : INV_X1 port map( A => A(34), ZN => n183);
   U390 : XNOR2_X1 port map( A => n265, B => n54, ZN => SUM(51));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_10_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_10_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_10_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_29_port, carry_1_port, net63046, net63041, 
      net62943, net63048, net62948, net68252, carry_62_port, net63042, 
      carry_61_port, carry_60_port, carry_59_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_12_port, carry_11_port, carry_10_port, net105170, 
      net105143, net105141, net84782, net93362, net84598, net84590, net84589, 
      net84134, net84133, carry_28_port, carry_27_port, carry_26_port, 
      carry_25_port, carry_24_port, carry_23_port, carry_22_port, carry_21_port
      , carry_20_port, carry_19_port, carry_18_port, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_59 : FA_X1 port map( A => carry_59_port, B => B(59), CI => A(59), CO => 
                           carry_60_port, S => SUM(59));
   U1_61 : FA_X1 port map( A => carry_61_port, B => B(61), CI => A(61), CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1 : OAI21_X1 port map( B1 => n133, B2 => n134, A => n135, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n75, A2 => B(31), ZN => n2);
   U3 : NAND2_X1 port map( A1 => carry_12_port, A2 => B(12), ZN => n12);
   U4 : INV_X1 port map( A => B(44), ZN => n179);
   U5 : INV_X1 port map( A => B(52), ZN => n183);
   U6 : INV_X1 port map( A => B(14), ZN => n23);
   U7 : INV_X1 port map( A => B(15), ZN => n24);
   U8 : INV_X1 port map( A => B(36), ZN => n175);
   U9 : INV_X1 port map( A => B(40), ZN => n177);
   U10 : INV_X1 port map( A => B(48), ZN => n181);
   U11 : NAND2_X1 port map( A1 => net84782, A2 => B(17), ZN => net84134);
   U12 : INV_X1 port map( A => B(32), ZN => n173);
   U13 : INV_X1 port map( A => B(51), ZN => n182);
   U14 : INV_X1 port map( A => B(56), ZN => n69);
   U15 : XNOR2_X1 port map( A => carry_12_port, B => B(12), ZN => n27);
   U16 : XNOR2_X1 port map( A => n26, B => n16, ZN => SUM(13));
   U17 : INV_X1 port map( A => B(13), ZN => n22);
   U18 : INV_X1 port map( A => B(31), ZN => n172);
   U19 : INV_X1 port map( A => B(30), ZN => n171);
   U20 : INV_X1 port map( A => B(39), ZN => n176);
   U21 : INV_X1 port map( A => B(43), ZN => n178);
   U22 : INV_X1 port map( A => B(47), ZN => n180);
   U23 : INV_X1 port map( A => B(35), ZN => n174);
   U24 : OAI21_X1 port map( B1 => n6, B2 => net105141, A => net105143, ZN => n5
                           );
   U25 : INV_X1 port map( A => A(15), ZN => n6);
   U26 : AND3_X1 port map( A1 => n122, A2 => n123, A3 => n178, ZN => n125);
   U27 : NAND3_X1 port map( A1 => net84589, A2 => net84590, A3 => n4, ZN => 
                           carry_22_port);
   U28 : NAND2_X1 port map( A1 => A(21), A2 => B(21), ZN => n4);
   U29 : NAND2_X1 port map( A1 => carry_21_port, A2 => A(21), ZN => net84589);
   U30 : NAND2_X1 port map( A1 => carry_21_port, A2 => B(21), ZN => net84590);
   U31 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => net93362);
   U32 : XNOR2_X1 port map( A => carry_21_port, B => net93362, ZN => SUM(21));
   U33 : NAND3_X1 port map( A1 => net84133, A2 => net84134, A3 => n3, ZN => 
                           carry_18_port);
   U34 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n3);
   U35 : NAND2_X1 port map( A1 => net84782, A2 => A(17), ZN => net84133);
   U36 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => net84598);
   U37 : XNOR2_X1 port map( A => net84782, B => net84598, ZN => SUM(17));
   U38 : NAND2_X2 port map( A1 => n7, A2 => n8, ZN => net84782);
   U39 : OAI21_X1 port map( B1 => n10, B2 => B(16), A => A(16), ZN => n8);
   U40 : OAI21_X1 port map( B1 => net105141, B2 => n6, A => net105143, ZN => 
                           n10);
   U41 : XNOR2_X1 port map( A => net105170, B => n6, ZN => SUM(15));
   U42 : NAND2_X1 port map( A1 => B(16), A2 => n5, ZN => n7);
   U43 : XNOR2_X1 port map( A => n5, B => B(16), ZN => n9);
   U44 : XNOR2_X1 port map( A => A(16), B => n9, ZN => SUM(16));
   U45 : OAI21_X1 port map( B1 => B(12), B2 => carry_12_port, A => A(12), ZN =>
                           n13);
   U46 : XNOR2_X1 port map( A => A(12), B => n27, ZN => SUM(12));
   U47 : NOR2_X1 port map( A1 => n18, A2 => B(15), ZN => net105141);
   U48 : XNOR2_X1 port map( A => n29, B => n23, ZN => n25);
   U49 : NAND2_X1 port map( A1 => n29, A2 => B(14), ZN => n21);
   U50 : NOR2_X1 port map( A1 => n14, A2 => B(14), ZN => n19);
   U51 : OAI21_X1 port map( B1 => n20, B2 => n19, A => n21, ZN => n18);
   U52 : XNOR2_X1 port map( A => n28, B => n24, ZN => net105170);
   U53 : NAND2_X1 port map( A1 => n28, A2 => B(15), ZN => net105143);
   U54 : OAI21_X1 port map( B1 => n19, B2 => n20, A => n21, ZN => n28);
   U55 : NAND2_X1 port map( A1 => n13, A2 => n12, ZN => n11);
   U56 : XNOR2_X1 port map( A => n11, B => n22, ZN => n26);
   U57 : NAND2_X1 port map( A1 => B(13), A2 => n11, ZN => n17);
   U58 : NOR2_X1 port map( A1 => B(13), A2 => n11, ZN => n15);
   U59 : INV_X1 port map( A => A(13), ZN => n16);
   U60 : OAI21_X1 port map( B1 => n15, B2 => n16, A => n17, ZN => n14);
   U61 : OAI21_X1 port map( B1 => n15, B2 => n30, A => n17, ZN => n29);
   U62 : XNOR2_X1 port map( A => n25, B => n20, ZN => SUM(14));
   U63 : INV_X1 port map( A => A(13), ZN => n30);
   U64 : INV_X1 port map( A => A(14), ZN => n20);
   U65 : OAI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n31);
   U66 : CLKBUF_X1 port map( A => A(29), Z => n32);
   U67 : AND2_X1 port map( A1 => n74, A2 => n33, ZN => n76);
   U68 : AND2_X1 port map( A1 => n73, A2 => n171, ZN => n33);
   U69 : AND2_X1 port map( A1 => n137, A2 => n34, ZN => n139);
   U70 : AND2_X1 port map( A1 => n136, A2 => n180, ZN => n34);
   U71 : NOR2_X1 port map( A1 => B(52), A2 => n223, ZN => n35);
   U72 : NOR2_X1 port map( A1 => n94, A2 => B(36), ZN => n36);
   U73 : NOR2_X1 port map( A1 => B(35), A2 => n91, ZN => n37);
   U74 : INV_X1 port map( A => n104, ZN => n38);
   U75 : OAI21_X1 port map( B1 => B(34), B2 => n87, A => A(34), ZN => n39);
   U76 : NAND2_X1 port map( A1 => n92, A2 => n39, ZN => n40);
   U77 : NOR2_X1 port map( A1 => n217, A2 => B(37), ZN => n41);
   U78 : XNOR2_X1 port map( A => n209, B => n77, ZN => SUM(30));
   U79 : INV_X1 port map( A => A(44), ZN => n42);
   U80 : CLKBUF_X1 port map( A => A(50), Z => n58);
   U81 : AND2_X1 port map( A1 => n108, A2 => n43, ZN => n110);
   U82 : AND2_X1 port map( A1 => n107, A2 => n176, ZN => n43);
   U83 : CLKBUF_X1 port map( A => A(45), Z => n44);
   U84 : NAND2_X1 port map( A1 => B(35), A2 => n40, ZN => n97);
   U85 : NOR2_X1 port map( A1 => B(45), A2 => n128, ZN => n45);
   U86 : NOR2_X1 port map( A1 => n83, A2 => B(33), ZN => n46);
   U87 : NOR2_X1 port map( A1 => n79, A2 => B(32), ZN => n47);
   U88 : NOR2_X1 port map( A1 => n216, A2 => B(41), ZN => n48);
   U89 : NOR2_X1 port map( A1 => n230, A2 => B(40), ZN => n49);
   U90 : OAI21_X1 port map( B1 => n50, B2 => n51, A => n52, ZN => carry_59_port
                           );
   U91 : NAND2_X1 port map( A1 => B(58), A2 => n53, ZN => n52);
   U92 : NOR2_X1 port map( A1 => B(58), A2 => n53, ZN => n51);
   U93 : INV_X1 port map( A => A(58), ZN => n50);
   U94 : XNOR2_X1 port map( A => n55, B => B(58), ZN => n54);
   U95 : OAI21_X1 port map( B1 => net63042, B2 => net63041, A => net63046, ZN 
                           => n53);
   U96 : INV_X1 port map( A => A(57), ZN => net63042);
   U97 : OAI21_X1 port map( B1 => net63041, B2 => net63042, A => net63046, ZN 
                           => n55);
   U98 : XNOR2_X1 port map( A => n54, B => A(58), ZN => SUM(58));
   U99 : CLKBUF_X1 port map( A => A(57), Z => net68252);
   U100 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => n56);
   U101 : CLKBUF_X1 port map( A => A(46), Z => n57);
   U102 : CLKBUF_X1 port map( A => A(54), Z => n59);
   U103 : BUF_X1 port map( A => A(49), Z => n60);
   U104 : INV_X1 port map( A => A(47), ZN => n61);
   U105 : NAND2_X1 port map( A1 => B(39), A2 => n106, ZN => n112);
   U106 : XNOR2_X1 port map( A => n106, B => n176, ZN => n200);
   U107 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => n91);
   U108 : CLKBUF_X1 port map( A => A(53), Z => n62);
   U109 : OAI21_X1 port map( B1 => n140, B2 => n139, A => n141, ZN => n63);
   U110 : OAI21_X1 port map( B1 => n61, B2 => n139, A => n141, ZN => n138);
   U111 : XNOR2_X1 port map( A => n203, B => n100, ZN => SUM(36));
   U112 : XNOR2_X1 port map( A => n56, B => n180, ZN => n192);
   U113 : XNOR2_X1 port map( A => n187, B => n159, ZN => SUM(52));
   U114 : INV_X1 port map( A => A(51), ZN => n155);
   U115 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => n106);
   U116 : NAND2_X1 port map( A1 => n151, A2 => n152, ZN => n150);
   U117 : XNOR2_X1 port map( A => n121, B => n178, ZN => n196);
   U118 : NAND2_X1 port map( A1 => n121, A2 => B(43), ZN => n127);
   U119 : XNOR2_X1 port map( A => n40, B => n174, ZN => n204);
   U120 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => n64);
   U121 : XNOR2_X1 port map( A => n191, B => n144, ZN => SUM(48));
   U122 : CLKBUF_X1 port map( A => A(55), Z => n65);
   U123 : INV_X1 port map( A => A(36), ZN => n100);
   U124 : INV_X1 port map( A => A(48), ZN => n144);
   U125 : XNOR2_X1 port map( A => n70, B => n67, ZN => SUM(56));
   U126 : INV_X1 port map( A => A(44), ZN => n130);
   U127 : XNOR2_X1 port map( A => n200, B => n111, ZN => SUM(39));
   U128 : OAI21_X1 port map( B1 => n67, B2 => n66, A => n68, ZN => n71);
   U129 : XNOR2_X1 port map( A => n71, B => B(57), ZN => net63048);
   U130 : INV_X1 port map( A => A(56), ZN => n67);
   U131 : OAI21_X1 port map( B1 => n67, B2 => n66, A => n68, ZN => net62948);
   U132 : NOR2_X1 port map( A1 => B(56), A2 => net62943, ZN => n66);
   U133 : NAND2_X1 port map( A1 => B(56), A2 => n64, ZN => n68);
   U134 : XNOR2_X1 port map( A => n64, B => n69, ZN => n70);
   U135 : XNOR2_X1 port map( A => net63048, B => net68252, ZN => SUM(57));
   U136 : NAND2_X1 port map( A1 => net62948, A2 => B(57), ZN => net63046);
   U137 : NOR2_X1 port map( A1 => net62948, A2 => B(57), ZN => net63041);
   U138 : OAI21_X1 port map( B1 => B(50), B2 => n219, A => A(50), ZN => n152);
   U139 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => n121);
   U140 : INV_X1 port map( A => A(30), ZN => n77);
   U141 : XNOR2_X1 port map( A => n199, B => n115, ZN => SUM(40));
   U142 : XNOR2_X1 port map( A => n204, B => n96, ZN => SUM(35));
   U143 : XNOR2_X1 port map( A => n196, B => n126, ZN => SUM(43));
   U144 : XNOR2_X1 port map( A => n195, B => n42, ZN => SUM(44));
   U145 : XNOR2_X1 port map( A => n192, B => n61, ZN => SUM(47));
   U146 : NOR2_X1 port map( A1 => B(53), A2 => n225, ZN => n162);
   U147 : OAI21_X1 port map( B1 => n162, B2 => n163, A => n164, ZN => n161);
   U148 : OAI21_X1 port map( B1 => n224, B2 => n163, A => n164, ZN => n211);
   U149 : OAI21_X1 port map( B1 => n224, B2 => n163, A => n164, ZN => n212);
   U150 : NOR2_X1 port map( A1 => B(48), A2 => n227, ZN => n143);
   U151 : OAI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n142);
   U152 : OAI21_X1 port map( B1 => n226, B2 => n144, A => n145, ZN => n213);
   U153 : OAI21_X1 port map( B1 => n144, B2 => n226, A => n145, ZN => n214);
   U154 : NOR2_X1 port map( A1 => B(44), A2 => n229, ZN => n129);
   U155 : OAI21_X1 port map( B1 => n129, B2 => n130, A => n131, ZN => n128);
   U156 : OAI21_X1 port map( B1 => n228, B2 => n42, A => n131, ZN => n215);
   U157 : OAI21_X1 port map( B1 => n114, B2 => n115, A => n116, ZN => n113);
   U158 : NAND2_X1 port map( A1 => n113, A2 => B(41), ZN => n120);
   U159 : XNOR2_X1 port map( A => n113, B => B(41), ZN => n198);
   U160 : NOR2_X1 port map( A1 => B(41), A2 => n216, ZN => n118);
   U161 : NOR2_X1 port map( A1 => n109, A2 => B(40), ZN => n114);
   U162 : OAI21_X1 port map( B1 => n49, B2 => n115, A => n116, ZN => n216);
   U163 : OAI21_X1 port map( B1 => n99, B2 => n100, A => n101, ZN => n98);
   U164 : NAND2_X1 port map( A1 => n98, A2 => B(37), ZN => n105);
   U165 : XNOR2_X1 port map( A => n217, B => B(37), ZN => n202);
   U166 : NOR2_X1 port map( A1 => n98, A2 => B(37), ZN => n103);
   U167 : NOR2_X1 port map( A1 => n94, A2 => B(36), ZN => n99);
   U168 : OAI21_X1 port map( B1 => n36, B2 => n100, A => n101, ZN => n217);
   U169 : OAI21_X1 port map( B1 => n47, B2 => n85, A => n86, ZN => n83);
   U170 : NAND2_X1 port map( A1 => n233, A2 => B(33), ZN => n90);
   U171 : XNOR2_X1 port map( A => n233, B => B(33), ZN => n206);
   U172 : NOR2_X1 port map( A1 => B(33), A2 => n83, ZN => n88);
   U173 : NOR2_X1 port map( A1 => n232, A2 => B(32), ZN => n84);
   U174 : NOR2_X1 port map( A1 => B(54), A2 => n161, ZN => n166);
   U175 : OAI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => n165);
   U176 : OAI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => n218);
   U177 : NOR2_X1 port map( A1 => B(49), A2 => n142, ZN => n147);
   U178 : OAI21_X1 port map( B1 => n147, B2 => n148, A => n149, ZN => n146);
   U179 : OAI21_X1 port map( B1 => n147, B2 => n148, A => n149, ZN => n219);
   U180 : OAI21_X1 port map( B1 => n134, B2 => n45, A => n135, ZN => n132);
   U181 : NOR2_X1 port map( A1 => n128, A2 => B(45), ZN => n133);
   U182 : OAI21_X1 port map( B1 => n48, B2 => n119, A => n120, ZN => n117);
   U183 : NAND2_X1 port map( A1 => B(42), A2 => n220, ZN => n122);
   U184 : OAI21_X1 port map( B1 => B(42), B2 => n117, A => A(42), ZN => n123);
   U185 : XNOR2_X1 port map( A => B(42), B => n220, ZN => n197);
   U186 : OAI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n220);
   U187 : OAI21_X1 port map( B1 => n103, B2 => n104, A => n105, ZN => n102);
   U188 : NAND2_X1 port map( A1 => n102, A2 => B(38), ZN => n107);
   U189 : OAI21_X1 port map( B1 => B(38), B2 => n102, A => A(38), ZN => n108);
   U190 : XNOR2_X1 port map( A => n221, B => B(38), ZN => n201);
   U191 : OAI21_X1 port map( B1 => n41, B2 => n104, A => n105, ZN => n221);
   U192 : OAI21_X1 port map( B1 => n46, B2 => n89, A => n90, ZN => n87);
   U193 : NAND2_X1 port map( A1 => n222, A2 => B(34), ZN => n92);
   U194 : OAI21_X1 port map( B1 => B(34), B2 => n87, A => A(34), ZN => n93);
   U195 : XNOR2_X1 port map( A => n222, B => B(34), ZN => n205);
   U196 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n222);
   U197 : OAI21_X1 port map( B1 => n154, B2 => n155, A => n156, ZN => n153);
   U198 : XNOR2_X1 port map( A => n153, B => n183, ZN => n187);
   U199 : NAND2_X1 port map( A1 => n153, A2 => B(52), ZN => n160);
   U200 : NOR2_X1 port map( A1 => B(52), A2 => n223, ZN => n158);
   U201 : NOR2_X1 port map( A1 => B(51), A2 => n150, ZN => n154);
   U202 : OAI21_X1 port map( B1 => n154, B2 => n155, A => n156, ZN => n223);
   U203 : OAI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n75);
   U204 : XNOR2_X1 port map( A => n75, B => n172, ZN => n208);
   U205 : NAND2_X1 port map( A1 => n31, A2 => B(31), ZN => n82);
   U206 : NOR2_X1 port map( A1 => n31, A2 => B(31), ZN => n80);
   U207 : NOR2_X1 port map( A1 => B(53), A2 => n157, ZN => n224);
   U208 : OAI21_X1 port map( B1 => n159, B2 => n158, A => n160, ZN => n157);
   U209 : NAND2_X1 port map( A1 => n225, A2 => B(53), ZN => n164);
   U210 : XNOR2_X1 port map( A => n157, B => B(53), ZN => n186);
   U211 : OAI21_X1 port map( B1 => n35, B2 => n159, A => n160, ZN => n225);
   U212 : NOR2_X1 port map( A1 => n227, A2 => B(48), ZN => n226);
   U213 : XNOR2_X1 port map( A => n63, B => n181, ZN => n191);
   U214 : NAND2_X1 port map( A1 => n138, A2 => B(48), ZN => n145);
   U215 : OAI21_X1 port map( B1 => n139, B2 => n140, A => n141, ZN => n227);
   U216 : NOR2_X1 port map( A1 => n124, A2 => B(44), ZN => n228);
   U217 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n124);
   U218 : XNOR2_X1 port map( A => n124, B => n179, ZN => n195);
   U219 : NAND2_X1 port map( A1 => n229, A2 => B(44), ZN => n131);
   U220 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n229);
   U221 : XNOR2_X1 port map( A => n186, B => n62, ZN => SUM(53));
   U222 : OAI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n109);
   U223 : XNOR2_X1 port map( A => n109, B => n177, ZN => n199);
   U224 : NAND2_X1 port map( A1 => n230, A2 => B(40), ZN => n116);
   U225 : OAI21_X1 port map( B1 => n111, B2 => n110, A => n112, ZN => n230);
   U226 : OAI21_X1 port map( B1 => n37, B2 => n96, A => n97, ZN => n94);
   U227 : XNOR2_X1 port map( A => n231, B => n175, ZN => n203);
   U228 : NAND2_X1 port map( A1 => n231, A2 => B(36), ZN => n101);
   U229 : NOR2_X1 port map( A1 => B(35), A2 => n91, ZN => n95);
   U230 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n231);
   U231 : OAI21_X1 port map( B1 => n2, B2 => n81, A => n82, ZN => n79);
   U232 : XNOR2_X1 port map( A => n79, B => n173, ZN => n207);
   U233 : NAND2_X1 port map( A1 => n232, A2 => B(32), ZN => n86);
   U234 : XNOR2_X1 port map( A => n146, B => B(50), ZN => n189);
   U235 : NAND2_X1 port map( A1 => B(50), A2 => n219, ZN => n151);
   U236 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => n232);
   U237 : XNOR2_X1 port map( A => B(55), B => n165, ZN => n184);
   U238 : NAND2_X1 port map( A1 => B(55), A2 => n218, ZN => n169);
   U239 : NAND2_X1 port map( A1 => A(29), A2 => B(29), ZN => n73);
   U240 : OAI21_X1 port map( B1 => B(29), B2 => A(29), A => carry_29_port, ZN 
                           => n74);
   U241 : XNOR2_X1 port map( A => n210, B => n32, ZN => SUM(29));
   U242 : NAND2_X1 port map( A1 => n215, A2 => B(45), ZN => n135);
   U243 : INV_X1 port map( A => A(45), ZN => n134);
   U244 : XNOR2_X1 port map( A => n132, B => B(46), ZN => n193);
   U245 : NAND2_X1 port map( A1 => n1, A2 => B(46), ZN => n136);
   U246 : NAND2_X1 port map( A1 => n56, A2 => B(47), ZN => n141);
   U247 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => n72);
   U248 : INV_X1 port map( A => A(53), ZN => n163);
   U249 : NAND2_X1 port map( A1 => n150, A2 => B(51), ZN => n156);
   U250 : XNOR2_X1 port map( A => n189, B => n58, ZN => SUM(50));
   U251 : INV_X1 port map( A => A(52), ZN => n159);
   U252 : XNOR2_X1 port map( A => n213, B => B(49), ZN => n190);
   U253 : XNOR2_X1 port map( A => n215, B => B(45), ZN => n194);
   U254 : OAI21_X1 port map( B1 => n218, B2 => B(55), A => A(55), ZN => n170);
   U255 : XNOR2_X1 port map( A => n65, B => n184, ZN => SUM(55));
   U256 : XNOR2_X1 port map( A => A(34), B => n205, ZN => SUM(34));
   U257 : XNOR2_X1 port map( A => n197, B => A(42), ZN => SUM(42));
   U258 : XNOR2_X1 port map( A => n201, B => A(38), ZN => SUM(38));
   U259 : XNOR2_X1 port map( A => n206, B => A(33), ZN => SUM(33));
   U260 : XNOR2_X1 port map( A => n198, B => A(41), ZN => SUM(41));
   U261 : XNOR2_X1 port map( A => n211, B => B(54), ZN => n185);
   U262 : NAND2_X1 port map( A1 => B(49), A2 => n214, ZN => n149);
   U263 : INV_X1 port map( A => A(49), ZN => n148);
   U264 : NAND2_X1 port map( A1 => B(54), A2 => n212, ZN => n168);
   U265 : INV_X1 port map( A => A(54), ZN => n167);
   U266 : OAI21_X1 port map( B1 => n1, B2 => B(46), A => A(46), ZN => n137);
   U267 : XNOR2_X1 port map( A => n193, B => n57, ZN => SUM(46));
   U268 : XNOR2_X1 port map( A => n208, B => n81, ZN => SUM(31));
   U269 : INV_X1 port map( A => A(37), ZN => n104);
   U270 : XNOR2_X1 port map( A => n150, B => n182, ZN => n188);
   U271 : XNOR2_X1 port map( A => n188, B => n155, ZN => SUM(51));
   U272 : XNOR2_X1 port map( A => n72, B => n171, ZN => n209);
   U273 : NAND2_X1 port map( A1 => B(30), A2 => n72, ZN => n78);
   U274 : XNOR2_X1 port map( A => n202, B => n38, ZN => SUM(37));
   U275 : XNOR2_X1 port map( A => carry_29_port, B => B(29), ZN => n210);
   U276 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => net62943);
   U277 : INV_X1 port map( A => A(47), ZN => n140);
   U278 : XNOR2_X1 port map( A => n44, B => n194, ZN => SUM(45));
   U279 : XNOR2_X1 port map( A => n190, B => n60, ZN => SUM(49));
   U280 : INV_X1 port map( A => A(33), ZN => n89);
   U281 : INV_X1 port map( A => A(31), ZN => n81);
   U282 : INV_X1 port map( A => A(43), ZN => n126);
   U283 : INV_X1 port map( A => A(32), ZN => n85);
   U284 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n233);
   U285 : INV_X1 port map( A => A(35), ZN => n96);
   U286 : INV_X1 port map( A => A(39), ZN => n111);
   U287 : INV_X1 port map( A => A(40), ZN => n115);
   U288 : INV_X1 port map( A => A(41), ZN => n119);
   U289 : XNOR2_X1 port map( A => n185, B => n59, ZN => SUM(54));
   U290 : XNOR2_X1 port map( A => n207, B => n85, ZN => SUM(32));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_11_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_11_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_11_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_28_port, 
      carry_27_port, carry_31_port, carry_30_port, carry_29_port, net65157, 
      net65109, net65108, net65107, net65097, net65016, net65015, net65014, 
      net64999, net64997, net64984, net65137, net65110, net64990, net70144, 
      net70164, net70301, net70408, net70411, net65146, net64998, net64996, 
      net65106, net65104, net70422, net65136, net65101, net65100, net65009, 
      net65007, net70443, net70247, net65162, net65010, net65008, net65004, 
      net65003, net65002, carry_26_port, net83984, net83981, net83841, net83840
      , net83839, net83830, net83828, net83824, net83822, net83818, net83817, 
      net83816, net83807, net83805, net84535, net83810, net90417, net84026, 
      net83821, net83980, net83833, net83829, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1 : CLKBUF_X1 port map( A => A(20), Z => n1);
   U2 : OAI21_X1 port map( B1 => n224, B2 => n225, A => n226, ZN => n2);
   U3 : BUF_X1 port map( A => n34, Z => n3);
   U4 : CLKBUF_X1 port map( A => A(22), Z => n4);
   U5 : BUF_X1 port map( A => net83810, Z => n12);
   U6 : AND2_X1 port map( A1 => n60, A2 => n5, ZN => n63);
   U7 : AND2_X1 port map( A1 => n61, A2 => n6, ZN => n5);
   U8 : INV_X1 port map( A => B(22), ZN => n6);
   U9 : NOR2_X1 port map( A1 => B(14), A2 => net83810, ZN => n7);
   U10 : NOR2_X1 port map( A1 => B(15), A2 => n49, ZN => n8);
   U11 : CLKBUF_X1 port map( A => A(31), Z => n9);
   U12 : NAND2_X1 port map( A1 => n308, A2 => B(35), ZN => n10);
   U13 : NAND3_X1 port map( A1 => n24, A2 => n25, A3 => n26, ZN => n11);
   U14 : NOR2_X1 port map( A1 => B(16), A2 => net83821, ZN => n13);
   U15 : CLKBUF_X1 port map( A => n144, Z => n14);
   U16 : CLKBUF_X1 port map( A => A(18), Z => net90417);
   U17 : INV_X1 port map( A => B(50), ZN => n277);
   U18 : INV_X1 port map( A => B(10), ZN => n43);
   U19 : INV_X1 port map( A => B(54), ZN => n278);
   U20 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n127);
   U21 : INV_X1 port map( A => n103, ZN => n128);
   U22 : INV_X1 port map( A => n101, ZN => n130);
   U23 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n133);
   U24 : NAND2_X1 port map( A1 => A(8), A2 => n94, ZN => n121);
   U25 : INV_X1 port map( A => B(33), ZN => n268);
   U26 : INV_X1 port map( A => B(37), ZN => n270);
   U27 : INV_X1 port map( A => B(46), ZN => n275);
   U28 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n125);
   U29 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n102);
   U30 : OAI221_X1 port map( B1 => n126, B2 => n74, C1 => n126, C2 => n73, A =>
                           n127, ZN => n103);
   U31 : INV_X1 port map( A => B(2), ZN => n73);
   U32 : INV_X1 port map( A => A(2), ZN => n74);
   U33 : INV_X1 port map( A => n105, ZN => n126);
   U34 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n100);
   U35 : OAI221_X1 port map( B1 => n128, B2 => n76, C1 => n128, C2 => n75, A =>
                           n129, ZN => n101);
   U36 : INV_X1 port map( A => B(3), ZN => n75);
   U37 : INV_X1 port map( A => A(3), ZN => n76);
   U38 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n129);
   U39 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n98);
   U40 : OAI221_X1 port map( B1 => n130, B2 => n78, C1 => n130, C2 => n77, A =>
                           n131, ZN => n99);
   U41 : INV_X1 port map( A => B(4), ZN => n77);
   U42 : INV_X1 port map( A => A(4), ZN => n78);
   U43 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n131);
   U44 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n96);
   U45 : OAI211_X1 port map( C1 => n132, C2 => n79, A => n120, B => n133, ZN =>
                           n97);
   U46 : INV_X1 port map( A => B(5), ZN => n79);
   U47 : INV_X1 port map( A => n99, ZN => n132);
   U48 : NAND2_X1 port map( A1 => A(5), A2 => n99, ZN => n120);
   U49 : INV_X1 port map( A => A(6), ZN => n81);
   U50 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n91);
   U51 : OAI211_X1 port map( C1 => n137, C2 => n84, A => n121, B => n138, ZN =>
                           n92);
   U52 : INV_X1 port map( A => B(8), ZN => n84);
   U53 : INV_X1 port map( A => n94, ZN => n137);
   U54 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n138);
   U55 : OAI222_X1 port map( A1 => n139, A2 => n85, B1 => n139, B2 => n86, C1 
                           => n86, C2 => n85, ZN => n117);
   U56 : INV_X1 port map( A => B(9), ZN => n85);
   U57 : INV_X1 port map( A => n92, ZN => n139);
   U58 : INV_X1 port map( A => A(9), ZN => n86);
   U59 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n115);
   U60 : INV_X1 port map( A => B(34), ZN => n269);
   U61 : INV_X1 port map( A => B(38), ZN => n271);
   U62 : INV_X1 port map( A => B(41), ZN => n272);
   U63 : INV_X1 port map( A => B(42), ZN => n273);
   U64 : INV_X1 port map( A => B(45), ZN => n274);
   U65 : XNOR2_X1 port map( A => B(0), B => CI, ZN => n118);
   U66 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n104);
   U67 : OAI211_X1 port map( C1 => n124, C2 => n72, A => n119, B => n125, ZN =>
                           n105);
   U68 : INV_X1 port map( A => n113, ZN => n124);
   U69 : INV_X1 port map( A => B(1), ZN => n72);
   U70 : NAND2_X1 port map( A1 => A(1), A2 => n113, ZN => n119);
   U71 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n112);
   U72 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => n113);
   U73 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n123);
   U74 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => CI, ZN => n122);
   U75 : XNOR2_X1 port map( A => n102, B => n103, ZN => SUM(3));
   U76 : XNOR2_X1 port map( A => n100, B => n101, ZN => SUM(4));
   U77 : XNOR2_X1 port map( A => n98, B => n99, ZN => SUM(5));
   U78 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n93);
   U79 : OAI221_X1 port map( B1 => n95, B2 => n83, C1 => n95, C2 => n82, A => 
                           n136, ZN => n94);
   U80 : INV_X1 port map( A => B(7), ZN => n82);
   U81 : INV_X1 port map( A => A(7), ZN => n83);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n136);
   U83 : XNOR2_X1 port map( A => n96, B => n97, ZN => SUM(6));
   U84 : INV_X1 port map( A => n135, ZN => n95);
   U85 : OAI222_X1 port map( A1 => n134, A2 => n80, B1 => n134, B2 => n81, C1 
                           => n81, C2 => n80, ZN => n135);
   U86 : INV_X1 port map( A => B(6), ZN => n80);
   U87 : INV_X1 port map( A => n97, ZN => n134);
   U88 : XNOR2_X1 port map( A => n91, B => n92, ZN => SUM(9));
   U89 : XNOR2_X1 port map( A => n116, B => n117, ZN => SUM(10));
   U90 : INV_X1 port map( A => B(49), ZN => n276);
   U91 : INV_X1 port map( A => B(58), ZN => net65097);
   U92 : XNOR2_X1 port map( A => A(0), B => n118, ZN => SUM(0));
   U93 : XNOR2_X1 port map( A => n104, B => n105, ZN => SUM(2));
   U94 : XNOR2_X1 port map( A => n112, B => n113, ZN => SUM(1));
   U95 : XNOR2_X1 port map( A => n93, B => n94, ZN => SUM(8));
   U96 : XNOR2_X1 port map( A => n95, B => n15, ZN => SUM(7));
   U97 : INV_X1 port map( A => B(53), ZN => n174);
   U98 : XOR2_X1 port map( A => B(7), B => A(7), Z => n15);
   U99 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n16);
   U100 : INV_X1 port map( A => n117, ZN => n41);
   U101 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n17);
   U102 : XNOR2_X1 port map( A => n17, B => n16, ZN => SUM(18));
   U103 : NOR2_X1 port map( A1 => B(18), A2 => net83833, ZN => net83839);
   U104 : NAND2_X1 port map( A1 => B(18), A2 => n16, ZN => net83841);
   U105 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => net83833);
   U106 : OAI21_X1 port map( B1 => B(17), B2 => n18, A => A(17), ZN => n20);
   U107 : OAI21_X1 port map( B1 => net83828, B2 => net83829, A => net83830, ZN 
                           => n18);
   U108 : INV_X1 port map( A => A(16), ZN => net83829);
   U109 : OAI21_X1 port map( B1 => n13, B2 => net83829, A => net83830, ZN => 
                           n22);
   U110 : NAND2_X1 port map( A1 => B(17), A2 => n22, ZN => n19);
   U111 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n21);
   U112 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => net83980);
   U113 : XNOR2_X1 port map( A => n21, B => n22, ZN => SUM(17));
   U114 : XOR2_X1 port map( A => A(30), B => B(30), Z => n23);
   U115 : XOR2_X1 port map( A => carry_30_port, B => n23, Z => SUM(30));
   U116 : NAND2_X1 port map( A1 => carry_30_port, A2 => A(30), ZN => n24);
   U117 : NAND2_X1 port map( A1 => carry_30_port, A2 => B(30), ZN => n25);
   U118 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n26);
   U119 : NAND3_X1 port map( A1 => n24, A2 => n25, A3 => n26, ZN => 
                           carry_31_port);
   U120 : XNOR2_X1 port map( A => net83980, B => net84026, ZN => SUM(16));
   U121 : NOR2_X1 port map( A1 => B(16), A2 => net83821, ZN => net83828);
   U122 : NAND2_X1 port map( A1 => B(16), A2 => net84026, ZN => net83830);
   U123 : OAI21_X1 port map( B1 => net83822, B2 => n27, A => net83824, ZN => 
                           net84026);
   U124 : INV_X1 port map( A => A(15), ZN => n27);
   U125 : OAI21_X1 port map( B1 => n8, B2 => n27, A => net83824, ZN => net83821
                           );
   U126 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => net83981);
   U127 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n33);
   U128 : OAI221_X1 port map( B1 => n41, B2 => n42, C1 => n41, C2 => n43, A => 
                           n44, ZN => n40);
   U129 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => n28);
   U130 : XNOR2_X1 port map( A => n28, B => n12, ZN => SUM(14));
   U131 : CLKBUF_X1 port map( A => A(14), Z => net84535);
   U132 : NOR2_X1 port map( A1 => B(14), A2 => net83810, ZN => net83816);
   U133 : NAND2_X1 port map( A1 => B(14), A2 => net83810, ZN => net83818);
   U134 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => net83810);
   U135 : OAI21_X1 port map( B1 => n29, B2 => B(13), A => A(13), ZN => n32);
   U136 : OAI21_X1 port map( B1 => net83805, B2 => n30, A => net83807, ZN => 
                           n29);
   U137 : INV_X1 port map( A => A(12), ZN => n30);
   U138 : OAI21_X1 port map( B1 => net83805, B2 => n30, A => net83807, ZN => 
                           n34);
   U139 : NAND2_X1 port map( A1 => B(13), A2 => n34, ZN => n31);
   U140 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => net83984);
   U141 : XNOR2_X1 port map( A => n33, B => n3, ZN => SUM(13));
   U142 : NOR2_X1 port map( A1 => B(24), A2 => n66, ZN => n35);
   U143 : NOR2_X1 port map( A1 => n313, A2 => B(54), ZN => n36);
   U144 : INV_X1 port map( A => A(33), ZN => n192);
   U145 : XNOR2_X1 port map( A => n115, B => n40, ZN => SUM(11));
   U146 : NAND2_X1 port map( A1 => B(11), A2 => n40, ZN => n48);
   U147 : INV_X1 port map( A => A(11), ZN => n47);
   U148 : NAND2_X1 port map( A1 => B(20), A2 => n141, ZN => n58);
   U149 : CLKBUF_X1 port map( A => A(21), Z => n37);
   U150 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n59);
   U151 : BUF_X1 port map( A => A(52), Z => n173);
   U152 : NOR2_X1 port map( A1 => B(53), A2 => n38, ZN => n262);
   U153 : NAND2_X1 port map( A1 => n259, A2 => n260, ZN => n38);
   U154 : CLKBUF_X1 port map( A => A(44), Z => n157);
   U155 : NAND2_X1 port map( A1 => B(24), A2 => n140, ZN => n90);
   U156 : XNOR2_X1 port map( A => n111, B => n141, ZN => SUM(20));
   U157 : CLKBUF_X1 port map( A => A(47), Z => n39);
   U158 : XNOR2_X1 port map( A => n114, B => n148, ZN => SUM(19));
   U159 : NOR2_X1 port map( A1 => B(23), A2 => n62, ZN => n67);
   U160 : OAI21_X1 port map( B1 => n145, B2 => n68, A => n69, ZN => n66);
   U161 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => n140);
   U162 : NOR2_X1 port map( A1 => B(19), A2 => n148, ZN => n52);
   U163 : OAI21_X1 port map( B1 => n52, B2 => n53, A => n54, ZN => n51);
   U164 : OAI21_X1 port map( B1 => n147, B2 => n53, A => n54, ZN => n141);
   U165 : NOR2_X1 port map( A1 => B(15), A2 => n49, ZN => net83822);
   U166 : OAI21_X1 port map( B1 => n46, B2 => n47, A => n48, ZN => n45);
   U167 : NAND2_X1 port map( A1 => B(12), A2 => n142, ZN => net83807);
   U168 : XNOR2_X1 port map( A => net83984, B => n142, ZN => SUM(12));
   U169 : NOR2_X1 port map( A1 => n45, A2 => B(12), ZN => net83805);
   U170 : NOR2_X1 port map( A1 => B(11), A2 => n40, ZN => n46);
   U171 : OAI21_X1 port map( B1 => n46, B2 => n47, A => n48, ZN => n142);
   U172 : NOR2_X1 port map( A1 => B(20), A2 => n51, ZN => n56);
   U173 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n55);
   U174 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n143);
   U175 : OAI21_X1 port map( B1 => n35, B2 => n88, A => n90, ZN => n89);
   U176 : OAI22_X1 port map( A1 => n144, A2 => B(25), B1 => n89, B2 => A(25), 
                           ZN => n71);
   U177 : XNOR2_X1 port map( A => n106, B => n14, ZN => SUM(25));
   U178 : NOR2_X1 port map( A1 => B(24), A2 => n66, ZN => n87);
   U179 : OAI21_X1 port map( B1 => n87, B2 => n88, A => n90, ZN => n144);
   U180 : NOR2_X1 port map( A1 => n71, A2 => n70, ZN => carry_26_port);
   U181 : NOR2_X1 port map( A1 => B(23), A2 => n146, ZN => n145);
   U182 : OAI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n62);
   U183 : OAI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n146);
   U184 : NAND2_X1 port map( A1 => n62, A2 => B(23), ZN => n69);
   U185 : NOR2_X1 port map( A1 => n50, A2 => B(19), ZN => n147);
   U186 : OAI21_X1 port map( B1 => net83839, B2 => net83840, A => net83841, ZN 
                           => n50);
   U187 : OAI21_X1 port map( B1 => net83839, B2 => net83840, A => net83841, ZN 
                           => n148);
   U188 : NAND2_X1 port map( A1 => B(19), A2 => n50, ZN => n54);
   U189 : OAI21_X1 port map( B1 => net83816, B2 => net83817, A => net83818, ZN 
                           => n49);
   U190 : NAND2_X1 port map( A1 => B(15), A2 => n149, ZN => net83824);
   U191 : XNOR2_X1 port map( A => net83981, B => n149, ZN => SUM(15));
   U192 : OAI21_X1 port map( B1 => n7, B2 => net83817, A => net83818, ZN => 
                           n149);
   U193 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n116);
   U194 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n44);
   U195 : INV_X1 port map( A => A(10), ZN => n42);
   U196 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n106);
   U197 : NOR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n70);
   U198 : INV_X1 port map( A => net84535, ZN => net83817);
   U199 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n108);
   U200 : INV_X1 port map( A => A(23), ZN => n68);
   U201 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n110);
   U202 : OAI21_X1 port map( B1 => B(21), B2 => n55, A => n37, ZN => n61);
   U203 : XNOR2_X1 port map( A => B(24), B => A(24), ZN => n107);
   U204 : INV_X1 port map( A => A(24), ZN => n88);
   U205 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n109);
   U206 : INV_X1 port map( A => n4, ZN => n64);
   U207 : XNOR2_X1 port map( A => n110, B => n143, ZN => SUM(21));
   U208 : NAND2_X1 port map( A1 => n143, A2 => B(21), ZN => n60);
   U209 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n114);
   U210 : INV_X1 port map( A => A(19), ZN => n53);
   U211 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n111);
   U212 : INV_X1 port map( A => n1, ZN => n57);
   U213 : INV_X1 port map( A => net90417, ZN => net83840);
   U214 : NAND2_X1 port map( A1 => B(22), A2 => n59, ZN => n65);
   U215 : XNOR2_X1 port map( A => n108, B => n146, ZN => SUM(23));
   U216 : XNOR2_X1 port map( A => n140, B => n107, ZN => SUM(24));
   U217 : XNOR2_X1 port map( A => n109, B => n59, ZN => SUM(22));
   U218 : NOR2_X1 port map( A1 => B(41), A2 => n216, ZN => n150);
   U219 : INV_X1 port map( A => n214, ZN => n151);
   U220 : OAI21_X1 port map( B1 => B(44), B2 => n310, A => A(44), ZN => n152);
   U221 : AND2_X1 port map( A1 => n185, A2 => n153, ZN => n187);
   U222 : AND2_X1 port map( A1 => n184, A2 => n160, ZN => n153);
   U223 : OAI21_X1 port map( B1 => n212, B2 => B(40), A => A(40), ZN => n154);
   U224 : NOR2_X1 port map( A1 => n208, A2 => B(39), ZN => n155);
   U225 : NOR2_X1 port map( A1 => n201, A2 => B(37), ZN => n156);
   U226 : NAND2_X1 port map( A1 => n217, A2 => n154, ZN => n158);
   U227 : NAND2_X1 port map( A1 => n152, A2 => n232, ZN => n159);
   U228 : INV_X1 port map( A => B(32), ZN => n160);
   U229 : NOR2_X1 port map( A1 => n2, A2 => B(43), ZN => n161);
   U230 : NOR2_X1 port map( A1 => n194, A2 => B(35), ZN => n162);
   U231 : NOR2_X1 port map( A1 => B(38), A2 => n204, ZN => n163);
   U232 : NOR2_X1 port map( A1 => B(42), A2 => n319, ZN => n164);
   U233 : NOR2_X1 port map( A1 => n190, A2 => B(34), ZN => n165);
   U234 : NOR2_X1 port map( A1 => n314, A2 => B(33), ZN => n166);
   U235 : NAND2_X1 port map( A1 => net65003, A2 => net65004, ZN => net65002);
   U236 : NAND2_X1 port map( A1 => B(58), A2 => net65002, ZN => net65010);
   U237 : NOR2_X1 port map( A1 => B(58), A2 => net65002, ZN => net70443);
   U238 : NOR2_X1 port map( A1 => B(58), A2 => net65002, ZN => net65008);
   U239 : NAND2_X1 port map( A1 => net65146, A2 => B(57), ZN => net65003);
   U240 : NAND2_X1 port map( A1 => net65004, A2 => net65003, ZN => net70411);
   U241 : OAI21_X1 port map( B1 => net65146, B2 => B(57), A => A(57), ZN => 
                           net65004);
   U242 : XNOR2_X1 port map( A => net64996, B => B(57), ZN => net65109);
   U243 : CLKBUF_X1 port map( A => A(57), Z => net70301);
   U244 : OAI21_X1 port map( B1 => net70247, B2 => net65008, A => net65010, ZN 
                           => net65162);
   U245 : NOR2_X1 port map( A1 => net65162, A2 => B(59), ZN => net65100);
   U246 : INV_X1 port map( A => A(58), ZN => net70247);
   U247 : OAI21_X1 port map( B1 => net70408, B2 => net70247, A => net65010, ZN 
                           => net65007);
   U248 : OAI21_X1 port map( B1 => net65009, B2 => net70443, A => net65010, ZN 
                           => net70422);
   U249 : INV_X1 port map( A => A(58), ZN => net65009);
   U250 : OAI21_X1 port map( B1 => net65100, B2 => net65101, A => n167, ZN => 
                           net65136);
   U251 : XNOR2_X1 port map( A => net65136, B => B(60), ZN => net65106);
   U252 : INV_X1 port map( A => A(59), ZN => net65101);
   U253 : OAI21_X1 port map( B1 => net65101, B2 => net65100, A => n167, ZN => 
                           net65104);
   U254 : NAND2_X1 port map( A1 => net70422, A2 => B(59), ZN => n167);
   U255 : XNOR2_X1 port map( A => net65009, B => net65108, ZN => SUM(58));
   U256 : CLKBUF_X1 port map( A => A(59), Z => net70164);
   U257 : XNOR2_X1 port map( A => net65007, B => B(59), ZN => net65107);
   U258 : XNOR2_X1 port map( A => net65106, B => A(60), ZN => SUM(60));
   U259 : NAND2_X1 port map( A1 => B(60), A2 => net65104, ZN => net65016);
   U260 : NOR2_X1 port map( A1 => B(60), A2 => net65104, ZN => net65015);
   U261 : OAI21_X1 port map( B1 => net64997, B2 => net64998, A => net64999, ZN 
                           => net65146);
   U262 : INV_X1 port map( A => A(56), ZN => net64998);
   U263 : OAI21_X1 port map( B1 => net64997, B2 => net64998, A => net64999, ZN 
                           => net64996);
   U264 : CLKBUF_X1 port map( A => A(56), Z => net70144);
   U265 : INV_X1 port map( A => A(60), ZN => net65014);
   U266 : INV_X1 port map( A => A(50), ZN => n168);
   U267 : NAND2_X1 port map( A1 => n303, A2 => B(51), ZN => n258);
   U268 : CLKBUF_X1 port map( A => A(51), Z => n169);
   U269 : INV_X1 port map( A => A(54), ZN => n170);
   U270 : NOR2_X1 port map( A1 => B(58), A2 => net70411, ZN => net70408);
   U271 : NOR2_X1 port map( A1 => B(51), A2 => n252, ZN => n171);
   U272 : NOR2_X1 port map( A1 => B(51), A2 => n252, ZN => n256);
   U273 : INV_X1 port map( A => A(45), ZN => n172);
   U274 : OAI21_X1 port map( B1 => n265, B2 => n266, A => n267, ZN => n175);
   U275 : NAND2_X1 port map( A1 => n259, A2 => n260, ZN => n176);
   U276 : XNOR2_X1 port map( A => n158, B => n272, ZN => n292);
   U277 : NAND2_X1 port map( A1 => B(41), A2 => n158, ZN => n222);
   U278 : INV_X1 port map( A => A(42), ZN => n225);
   U279 : INV_X1 port map( A => A(38), ZN => n210);
   U280 : XNOR2_X1 port map( A => n295, B => n210, ZN => SUM(38));
   U281 : NAND2_X1 port map( A1 => n217, A2 => n218, ZN => n216);
   U282 : INV_X1 port map( A => A(41), ZN => n221);
   U283 : XNOR2_X1 port map( A => n288, B => n235, ZN => SUM(45));
   U284 : XNOR2_X1 port map( A => n283, B => n168, ZN => SUM(50));
   U285 : XNOR2_X1 port map( A => n296, B => n206, ZN => SUM(37));
   U286 : INV_X1 port map( A => A(46), ZN => n239);
   U287 : XNOR2_X1 port map( A => n284, B => n250, ZN => SUM(49));
   U288 : OAI21_X1 port map( B1 => B(52), B2 => n255, A => A(52), ZN => n260);
   U289 : OAI21_X1 port map( B1 => net65014, B2 => net65015, A => net65016, ZN 
                           => carry_61_port);
   U290 : XNOR2_X1 port map( A => n300, B => n192, ZN => SUM(33));
   U291 : XNOR2_X1 port map( A => n301, B => n188, ZN => SUM(32));
   U292 : XNOR2_X1 port map( A => net65110, B => net70144, ZN => SUM(56));
   U293 : XNOR2_X1 port map( A => n245, B => n276, ZN => n284);
   U294 : INV_X1 port map( A => A(34), ZN => n196);
   U295 : XNOR2_X1 port map( A => n287, B => n239, ZN => SUM(46));
   U296 : OAI21_X1 port map( B1 => n178, B2 => n182, A => n179, ZN => n181);
   U297 : XNOR2_X1 port map( A => n181, B => B(56), ZN => net65110);
   U298 : INV_X1 port map( A => A(55), ZN => n178);
   U299 : OAI21_X1 port map( B1 => n182, B2 => n178, A => n179, ZN => net65137)
                           ;
   U300 : OAI21_X1 port map( B1 => n177, B2 => n178, A => n179, ZN => net64990)
                           ;
   U301 : NOR2_X1 port map( A1 => net65157, A2 => B(55), ZN => n182);
   U302 : NAND2_X1 port map( A1 => n175, A2 => B(55), ZN => n179);
   U303 : XNOR2_X1 port map( A => n180, B => A(55), ZN => SUM(55));
   U304 : XNOR2_X1 port map( A => net64984, B => B(55), ZN => n180);
   U305 : NOR2_X1 port map( A1 => B(55), A2 => n175, ZN => n177);
   U306 : NOR2_X1 port map( A1 => B(56), A2 => net64990, ZN => net64997);
   U307 : NAND2_X1 port map( A1 => B(56), A2 => net65137, ZN => net64999);
   U308 : XNOR2_X1 port map( A => n291, B => n225, ZN => SUM(42));
   U309 : XNOR2_X1 port map( A => n292, B => n221, ZN => SUM(41));
   U310 : NOR2_X1 port map( A1 => n316, A2 => B(50), ZN => n253);
   U311 : OAI21_X1 port map( B1 => n253, B2 => n168, A => n254, ZN => n252);
   U312 : OAI21_X1 port map( B1 => n315, B2 => n168, A => n254, ZN => n303);
   U313 : NOR2_X1 port map( A1 => B(46), A2 => n233, ZN => n238);
   U314 : OAI21_X1 port map( B1 => n238, B2 => n239, A => n240, ZN => n237);
   U315 : OAI21_X1 port map( B1 => n317, B2 => n239, A => n240, ZN => n304);
   U316 : OAI21_X1 port map( B1 => n239, B2 => n317, A => n240, ZN => n305);
   U317 : OAI21_X1 port map( B1 => n164, B2 => n225, A => n226, ZN => n223);
   U318 : NAND2_X1 port map( A1 => n306, A2 => B(43), ZN => n230);
   U319 : XNOR2_X1 port map( A => n223, B => B(43), ZN => n290);
   U320 : NOR2_X1 port map( A1 => B(43), A2 => n2, ZN => n228);
   U321 : NOR2_X1 port map( A1 => n219, A2 => B(42), ZN => n224);
   U322 : OAI21_X1 port map( B1 => n224, B2 => n225, A => n226, ZN => n306);
   U323 : OAI21_X1 port map( B1 => n163, B2 => n210, A => n211, ZN => n208);
   U324 : NAND2_X1 port map( A1 => n307, A2 => B(39), ZN => n215);
   U325 : XNOR2_X1 port map( A => n307, B => B(39), ZN => n294);
   U326 : NOR2_X1 port map( A1 => B(39), A2 => n208, ZN => n213);
   U327 : NOR2_X1 port map( A1 => n320, A2 => B(38), ZN => n209);
   U328 : OAI21_X1 port map( B1 => n209, B2 => n210, A => n211, ZN => n307);
   U329 : OAI21_X1 port map( B1 => n165, B2 => n196, A => n197, ZN => n194);
   U330 : XNOR2_X1 port map( A => n308, B => B(35), ZN => n298);
   U331 : NOR2_X1 port map( A1 => B(35), A2 => n194, ZN => n199);
   U332 : NOR2_X1 port map( A1 => n190, A2 => B(34), ZN => n195);
   U333 : OAI21_X1 port map( B1 => n195, B2 => n196, A => n197, ZN => n308);
   U334 : OAI21_X1 port map( B1 => n171, B2 => n257, A => n258, ZN => n255);
   U335 : NOR2_X1 port map( A1 => B(47), A2 => n237, ZN => n242);
   U336 : OAI21_X1 port map( B1 => n242, B2 => n243, A => n244, ZN => n241);
   U337 : OAI21_X1 port map( B1 => n242, B2 => n243, A => n244, ZN => n309);
   U338 : OAI21_X1 port map( B1 => n228, B2 => n229, A => n230, ZN => n227);
   U339 : NAND2_X1 port map( A1 => B(44), A2 => n310, ZN => n232);
   U340 : XNOR2_X1 port map( A => n227, B => B(44), ZN => n289);
   U341 : OAI21_X1 port map( B1 => n161, B2 => n229, A => n230, ZN => n310);
   U342 : OAI21_X1 port map( B1 => n155, B2 => n214, A => n215, ZN => n212);
   U343 : NAND2_X1 port map( A1 => n212, A2 => B(40), ZN => n217);
   U344 : OAI21_X1 port map( B1 => n212, B2 => B(40), A => A(40), ZN => n218);
   U345 : XNOR2_X1 port map( A => B(40), B => n311, ZN => n293);
   U346 : OAI21_X1 port map( B1 => n214, B2 => n213, A => n215, ZN => n311);
   U347 : OAI21_X1 port map( B1 => n162, B2 => n200, A => n10, ZN => n198);
   U348 : NAND2_X1 port map( A1 => B(36), A2 => n198, ZN => n202);
   U349 : OAI21_X1 port map( B1 => n198, B2 => B(36), A => A(36), ZN => n203);
   U350 : XNOR2_X1 port map( A => B(36), B => n312, ZN => n297);
   U351 : OAI21_X1 port map( B1 => n199, B2 => n200, A => n10, ZN => n312);
   U352 : OAI21_X1 port map( B1 => n262, B2 => n263, A => n264, ZN => n261);
   U353 : XNOR2_X1 port map( A => n261, B => n278, ZN => n279);
   U354 : NAND2_X1 port map( A1 => n261, A2 => B(54), ZN => n267);
   U355 : NOR2_X1 port map( A1 => n313, A2 => B(54), ZN => n265);
   U356 : OAI21_X1 port map( B1 => n262, B2 => n263, A => n264, ZN => n313);
   U357 : OAI21_X1 port map( B1 => n187, B2 => n188, A => n189, ZN => n186);
   U358 : XNOR2_X1 port map( A => n314, B => n268, ZN => n300);
   U359 : NAND2_X1 port map( A1 => n186, A2 => B(33), ZN => n193);
   U360 : NOR2_X1 port map( A1 => n186, A2 => B(33), ZN => n191);
   U361 : OAI21_X1 port map( B1 => n187, B2 => n188, A => n189, ZN => n314);
   U362 : OAI21_X1 port map( B1 => n36, B2 => n266, A => n267, ZN => net64984);
   U363 : OAI21_X1 port map( B1 => n170, B2 => n36, A => n267, ZN => net65157);
   U364 : NOR2_X1 port map( A1 => n316, A2 => B(50), ZN => n315);
   U365 : OAI21_X1 port map( B1 => n249, B2 => n250, A => n251, ZN => n248);
   U366 : XNOR2_X1 port map( A => n248, B => n277, ZN => n283);
   U367 : NAND2_X1 port map( A1 => n248, A2 => B(50), ZN => n254);
   U368 : NOR2_X1 port map( A1 => B(49), A2 => n245, ZN => n249);
   U369 : OAI21_X1 port map( B1 => n250, B2 => n249, A => n251, ZN => n316);
   U370 : NOR2_X1 port map( A1 => n233, A2 => B(46), ZN => n317);
   U371 : OAI21_X1 port map( B1 => n234, B2 => n235, A => n236, ZN => n233);
   U372 : XNOR2_X1 port map( A => n318, B => n275, ZN => n287);
   U373 : NAND2_X1 port map( A1 => n318, A2 => B(46), ZN => n240);
   U374 : NOR2_X1 port map( A1 => B(45), A2 => n231, ZN => n234);
   U375 : OAI21_X1 port map( B1 => n234, B2 => n172, A => n236, ZN => n318);
   U376 : OAI21_X1 port map( B1 => n220, B2 => n221, A => n222, ZN => n219);
   U377 : XNOR2_X1 port map( A => n319, B => n273, ZN => n291);
   U378 : NAND2_X1 port map( A1 => n219, A2 => B(42), ZN => n226);
   U379 : NOR2_X1 port map( A1 => B(41), A2 => n216, ZN => n220);
   U380 : OAI21_X1 port map( B1 => n150, B2 => n221, A => n222, ZN => n319);
   U381 : OAI21_X1 port map( B1 => n156, B2 => n206, A => n207, ZN => n204);
   U382 : XNOR2_X1 port map( A => n320, B => n271, ZN => n295);
   U383 : NAND2_X1 port map( A1 => n204, A2 => B(38), ZN => n211);
   U384 : NOR2_X1 port map( A1 => B(37), A2 => n201, ZN => n205);
   U385 : OAI21_X1 port map( B1 => n205, B2 => n206, A => n207, ZN => n320);
   U386 : OAI21_X1 port map( B1 => n166, B2 => n192, A => n193, ZN => n190);
   U387 : XNOR2_X1 port map( A => n321, B => n269, ZN => n299);
   U388 : NAND2_X1 port map( A1 => n321, A2 => B(34), ZN => n197);
   U389 : OAI21_X1 port map( B1 => n191, B2 => n192, A => n193, ZN => n321);
   U390 : XNOR2_X1 port map( A => n322, B => B(52), ZN => n281);
   U391 : NAND2_X1 port map( A1 => B(52), A2 => n255, ZN => n259);
   U392 : NAND2_X1 port map( A1 => B(49), A2 => n245, ZN => n251);
   U393 : NAND2_X1 port map( A1 => B(47), A2 => n305, ZN => n244);
   U394 : INV_X1 port map( A => A(47), ZN => n243);
   U395 : NAND2_X1 port map( A1 => n152, A2 => n232, ZN => n231);
   U396 : XNOR2_X1 port map( A => n309, B => B(48), ZN => n285);
   U397 : NAND2_X1 port map( A1 => B(48), A2 => n241, ZN => n246);
   U398 : XNOR2_X1 port map( A => n159, B => n274, ZN => n288);
   U399 : NAND2_X1 port map( A1 => n159, A2 => B(45), ZN => n236);
   U400 : NAND2_X1 port map( A1 => n176, A2 => B(53), ZN => n264);
   U401 : INV_X1 port map( A => A(54), ZN => n266);
   U402 : XNOR2_X1 port map( A => net65107, B => net70164, ZN => SUM(59));
   U403 : XNOR2_X1 port map( A => A(40), B => n293, ZN => SUM(40));
   U404 : XNOR2_X1 port map( A => n304, B => B(47), ZN => n286);
   U405 : XNOR2_X1 port map( A => A(36), B => n297, ZN => SUM(36));
   U406 : XNOR2_X1 port map( A => net65109, B => net70301, ZN => SUM(57));
   U407 : XNOR2_X1 port map( A => n281, B => n173, ZN => SUM(52));
   U408 : XNOR2_X1 port map( A => n299, B => n196, ZN => SUM(34));
   U409 : XNOR2_X1 port map( A => n11, B => B(31), ZN => n302);
   U410 : OAI21_X1 port map( B1 => A(31), B2 => B(31), A => carry_31_port, ZN 
                           => n185);
   U411 : XNOR2_X1 port map( A => n289, B => n157, ZN => SUM(44));
   U412 : XNOR2_X1 port map( A => n303, B => B(51), ZN => n282);
   U413 : NAND2_X1 port map( A1 => B(31), A2 => A(31), ZN => n184);
   U414 : XNOR2_X1 port map( A => n302, B => n9, ZN => SUM(31));
   U415 : OAI21_X1 port map( B1 => n241, B2 => B(48), A => A(48), ZN => n247);
   U416 : XNOR2_X1 port map( A => n285, B => A(48), ZN => SUM(48));
   U417 : XNOR2_X1 port map( A => n294, B => n151, ZN => SUM(39));
   U418 : XNOR2_X1 port map( A => n298, B => A(35), ZN => SUM(35));
   U419 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => n183);
   U420 : INV_X1 port map( A => A(43), ZN => n229);
   U421 : INV_X1 port map( A => A(51), ZN => n257);
   U422 : OAI21_X1 port map( B1 => n257, B2 => n256, A => n258, ZN => n322);
   U423 : XNOR2_X1 port map( A => n286, B => n39, ZN => SUM(47));
   U424 : XNOR2_X1 port map( A => n176, B => n174, ZN => n280);
   U425 : XNOR2_X1 port map( A => n280, B => n263, ZN => SUM(53));
   U426 : INV_X1 port map( A => A(35), ZN => n200);
   U427 : XNOR2_X1 port map( A => n183, B => n160, ZN => n301);
   U428 : NAND2_X1 port map( A1 => n183, A2 => B(32), ZN => n189);
   U429 : INV_X1 port map( A => A(37), ZN => n206);
   U430 : XNOR2_X1 port map( A => A(43), B => n290, ZN => SUM(43));
   U431 : INV_X1 port map( A => A(39), ZN => n214);
   U432 : INV_X1 port map( A => A(45), ZN => n235);
   U433 : INV_X1 port map( A => A(49), ZN => n250);
   U434 : XNOR2_X1 port map( A => net70411, B => net65097, ZN => net65108);
   U435 : INV_X1 port map( A => A(53), ZN => n263);
   U436 : XNOR2_X1 port map( A => n282, B => n169, ZN => SUM(51));
   U437 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => n201);
   U438 : XNOR2_X1 port map( A => n201, B => n270, ZN => n296);
   U439 : NAND2_X1 port map( A1 => n201, A2 => B(37), ZN => n207);
   U440 : INV_X1 port map( A => A(32), ZN => n188);
   U441 : XNOR2_X1 port map( A => n279, B => n170, ZN => SUM(54));
   U442 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => n245);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_12_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_12_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_12_DW01_add_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_27_port, carry_26_port, carry_25_port, carry_24_port
      , carry_23_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_28_port, net70461, carry_58_port, net84116, net84513, net84661, 
      net84660, net84796, net90269, net90287, net90373, carry_9_port, 
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, carry_1_port, carry_11_port, carry_10_port, 
      net84515, net84514, net84113, net84112, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_15_port, carry_14_port, carry_13_port
      , carry_12_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => carry_61_port, B => B(61), CI => A(61), CO => 
                           carry_62_port, S => SUM(61));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1 : XNOR2_X1 port map( A => n6, B => n1, ZN => SUM(13));
   U2 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n1);
   U3 : XNOR2_X1 port map( A => n3, B => n2, ZN => SUM(16));
   U4 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n2);
   U5 : CLKBUF_X1 port map( A => carry_16_port, Z => n3);
   U6 : BUF_X1 port map( A => A(16), Z => n4);
   U7 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => n12, ZN => n5);
   U8 : CLKBUF_X1 port map( A => carry_13_port, Z => n6);
   U9 : NAND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => n7);
   U10 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n8);
   U11 : NAND2_X1 port map( A1 => A(13), A2 => B(13), ZN => n9);
   U12 : NAND3_X1 port map( A1 => n7, A2 => n8, A3 => n9, ZN => carry_14_port);
   U13 : NAND2_X1 port map( A1 => carry_16_port, A2 => n4, ZN => n10);
   U14 : NAND2_X1 port map( A1 => carry_16_port, A2 => B(16), ZN => n11);
   U15 : NAND2_X1 port map( A1 => n4, A2 => B(16), ZN => n12);
   U16 : NAND3_X1 port map( A1 => n11, A2 => n10, A3 => n12, ZN => 
                           carry_17_port);
   U17 : CLKBUF_X1 port map( A => carry_21_port, Z => n13);
   U18 : AND2_X1 port map( A1 => n102, A2 => n14, ZN => n104);
   U19 : AND2_X1 port map( A1 => n101, A2 => n15, ZN => n14);
   U20 : INV_X1 port map( A => B(38), ZN => n15);
   U21 : NOR2_X1 port map( A1 => n78, A2 => B(32), ZN => n16);
   U22 : OAI21_X1 port map( B1 => n117, B2 => n116, A => n118, ZN => n17);
   U23 : AND2_X2 port map( A1 => n113, A2 => n50, ZN => n116);
   U24 : NAND2_X1 port map( A1 => B(50), A2 => n141, ZN => n147);
   U25 : INV_X1 port map( A => B(55), ZN => n181);
   U26 : INV_X1 port map( A => B(39), ZN => n174);
   U27 : INV_X1 port map( A => B(46), ZN => n177);
   U28 : INV_X1 port map( A => B(31), ZN => n171);
   U29 : INV_X1 port map( A => B(34), ZN => n172);
   U30 : INV_X1 port map( A => B(50), ZN => n179);
   U31 : INV_X1 port map( A => B(47), ZN => n178);
   U32 : INV_X1 port map( A => B(51), ZN => n180);
   U33 : INV_X1 port map( A => A(55), ZN => n164);
   U34 : INV_X1 port map( A => A(56), ZN => n183);
   U35 : INV_X1 port map( A => B(35), ZN => n173);
   U36 : INV_X1 port map( A => B(43), ZN => n176);
   U37 : INV_X1 port map( A => B(30), ZN => n170);
   U38 : XNOR2_X1 port map( A => n244, B => n66, ZN => SUM(60));
   U39 : XNOR2_X1 port map( A => n188, B => n164, ZN => SUM(55));
   U40 : INV_X1 port map( A => B(29), ZN => n169);
   U41 : INV_X1 port map( A => B(42), ZN => n175);
   U42 : INV_X1 port map( A => B(20), ZN => n29);
   U43 : XNOR2_X1 port map( A => carry_19_port, B => net90373, ZN => SUM(19));
   U44 : NAND2_X1 port map( A1 => carry_19_port, A2 => B(19), ZN => net84661);
   U45 : NAND2_X1 port map( A1 => carry_19_port, A2 => net90269, ZN => net84660
                           );
   U46 : NAND3_X1 port map( A1 => net84112, A2 => net84113, A3 => n18, ZN => 
                           carry_18_port);
   U47 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n18);
   U48 : NAND2_X1 port map( A1 => n5, A2 => B(17), ZN => net84113);
   U49 : NAND2_X1 port map( A1 => carry_17_port, A2 => A(17), ZN => net84112);
   U50 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => net84116);
   U51 : CLKBUF_X1 port map( A => carry_17_port, Z => net84796);
   U52 : NAND3_X1 port map( A1 => net84515, A2 => net84514, A3 => n19, ZN => 
                           carry_12_port);
   U53 : NAND2_X1 port map( A1 => A(11), A2 => B(11), ZN => n19);
   U54 : NAND2_X1 port map( A1 => carry_11_port, A2 => A(11), ZN => net84514);
   U55 : NAND2_X1 port map( A1 => carry_11_port, A2 => B(11), ZN => net84515);
   U56 : XOR2_X1 port map( A => A(11), B => B(11), Z => net84513);
   U57 : CLKBUF_X1 port map( A => carry_11_port, Z => net90287);
   U58 : NAND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => carry_9_port
                           );
   U59 : NAND2_X1 port map( A1 => A(8), A2 => B(8), ZN => n23);
   U60 : NAND2_X1 port map( A1 => carry_8_port, A2 => B(8), ZN => n22);
   U61 : NAND2_X1 port map( A1 => carry_8_port, A2 => n24, ZN => n21);
   U62 : CLKBUF_X1 port map( A => A(8), Z => n24);
   U63 : XOR2_X1 port map( A => n24, B => B(8), Z => n20);
   U64 : XOR2_X1 port map( A => carry_8_port, B => n20, Z => SUM(8));
   U65 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => net90373);
   U66 : CLKBUF_X1 port map( A => A(19), Z => net90269);
   U67 : NAND3_X1 port map( A1 => n42, A2 => n43, A3 => n44, ZN => n25);
   U68 : NOR2_X1 port map( A1 => B(51), A2 => n231, ZN => n26);
   U69 : OAI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n27);
   U70 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n30);
   U71 : CLKBUF_X1 port map( A => n25, Z => n28);
   U72 : XNOR2_X1 port map( A => A(20), B => n29, ZN => n35);
   U73 : XNOR2_X1 port map( A => n30, B => n28, ZN => SUM(22));
   U74 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n31);
   U75 : NAND3_X1 port map( A1 => net84660, A2 => net84661, A3 => n31, ZN => 
                           carry_20_port);
   U76 : CLKBUF_X1 port map( A => A(20), Z => n32);
   U77 : AND2_X1 port map( A1 => n69, A2 => n33, ZN => n71);
   U78 : AND2_X1 port map( A1 => n68, A2 => n169, ZN => n33);
   U79 : XOR2_X1 port map( A => net90287, B => net84513, Z => SUM(11));
   U80 : XNOR2_X1 port map( A => n13, B => n34, ZN => SUM(21));
   U81 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n34);
   U82 : XOR2_X1 port map( A => carry_20_port, B => n35, Z => SUM(20));
   U83 : NAND2_X1 port map( A1 => carry_20_port, A2 => n32, ZN => n36);
   U84 : NAND2_X1 port map( A1 => carry_20_port, A2 => B(20), ZN => n37);
   U85 : NAND2_X1 port map( A1 => A(20), A2 => B(20), ZN => n38);
   U86 : NAND3_X1 port map( A1 => n36, A2 => n37, A3 => n38, ZN => 
                           carry_21_port);
   U87 : CLKBUF_X1 port map( A => A(21), Z => n39);
   U88 : INV_X1 port map( A => n154, ZN => n40);
   U89 : CLKBUF_X1 port map( A => A(37), Z => n41);
   U90 : NAND2_X1 port map( A1 => carry_21_port, A2 => n39, ZN => n42);
   U91 : NAND2_X1 port map( A1 => carry_21_port, A2 => B(21), ZN => n43);
   U92 : NAND2_X1 port map( A1 => A(21), A2 => B(21), ZN => n44);
   U93 : NAND3_X1 port map( A1 => n43, A2 => n42, A3 => n44, ZN => 
                           carry_22_port);
   U94 : NAND2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => n45);
   U95 : NAND2_X1 port map( A1 => n25, A2 => B(22), ZN => n46);
   U96 : NAND2_X1 port map( A1 => A(22), A2 => B(22), ZN => n47);
   U97 : NAND3_X1 port map( A1 => n46, A2 => n45, A3 => n47, ZN => 
                           carry_23_port);
   U98 : INV_X1 port map( A => n158, ZN => n48);
   U99 : NAND2_X1 port map( A1 => B(55), A2 => n160, ZN => n165);
   U100 : XNOR2_X1 port map( A => n160, B => n181, ZN => n188);
   U101 : NAND2_X1 port map( A1 => n161, A2 => n162, ZN => n160);
   U102 : XNOR2_X1 port map( A => net84116, B => net84796, ZN => SUM(17));
   U103 : INV_X1 port map( A => A(46), ZN => n49);
   U104 : AND2_X1 port map( A1 => n114, A2 => n175, ZN => n50);
   U105 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => n51);
   U106 : XNOR2_X1 port map( A => n192, B => n150, ZN => SUM(51));
   U107 : XOR2_X1 port map( A => A(26), B => B(26), Z => n52);
   U108 : XOR2_X1 port map( A => carry_26_port, B => n52, Z => SUM(26));
   U109 : NAND2_X1 port map( A1 => carry_26_port, A2 => A(26), ZN => n53);
   U110 : NAND2_X1 port map( A1 => carry_26_port, A2 => B(26), ZN => n54);
   U111 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n55);
   U112 : NAND3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => 
                           carry_27_port);
   U113 : NOR2_X1 port map( A1 => B(34), A2 => n51, ZN => n56);
   U114 : XNOR2_X1 port map( A => n57, B => n175, ZN => n201);
   U115 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => n57);
   U116 : INV_X1 port map( A => A(57), ZN => n166);
   U117 : XNOR2_X1 port map( A => n212, B => n80, ZN => SUM(31));
   U118 : NOR2_X1 port map( A1 => n74, A2 => B(31), ZN => n58);
   U119 : NOR2_X1 port map( A1 => B(30), A2 => n70, ZN => n59);
   U120 : XNOR2_X1 port map( A => n213, B => n76, ZN => SUM(30));
   U121 : OAI21_X1 port map( B1 => n61, B2 => n63, A => n112, ZN => n60);
   U122 : XNOR2_X1 port map( A => n214, B => n72, ZN => SUM(29));
   U123 : XNOR2_X1 port map( A => n208, B => n94, ZN => SUM(35));
   U124 : XNOR2_X1 port map( A => n196, B => n135, ZN => SUM(47));
   U125 : INV_X1 port map( A => A(47), ZN => n135);
   U126 : XNOR2_X1 port map( A => n200, B => n121, ZN => SUM(43));
   U127 : INV_X1 port map( A => A(40), ZN => n61);
   U128 : NAND2_X1 port map( A1 => B(38), A2 => n100, ZN => n106);
   U129 : INV_X1 port map( A => n125, ZN => n62);
   U130 : INV_X1 port map( A => A(52), ZN => n154);
   U131 : INV_X1 port map( A => A(39), ZN => n109);
   U132 : INV_X1 port map( A => A(53), ZN => n158);
   U133 : XNOR2_X1 port map( A => n193, B => n146, ZN => SUM(50));
   U134 : NOR2_X1 port map( A1 => B(40), A2 => n107, ZN => n63);
   U135 : NOR2_X1 port map( A1 => n240, A2 => B(35), ZN => n64);
   U136 : INV_X1 port map( A => A(51), ZN => n150);
   U137 : XNOR2_X1 port map( A => n127, B => n177, ZN => n197);
   U138 : NAND2_X1 port map( A1 => B(46), A2 => n127, ZN => n132);
   U139 : XNOR2_X1 port map( A => n197, B => n49, ZN => SUM(46));
   U140 : INV_X1 port map( A => A(50), ZN => n146);
   U141 : INV_X1 port map( A => A(44), ZN => n125);
   U142 : INV_X1 port map( A => A(48), ZN => n139);
   U143 : INV_X1 port map( A => n61, ZN => n65);
   U144 : OAI21_X1 port map( B1 => B(54), B2 => n156, A => A(54), ZN => n162);
   U145 : OAI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => 
                           carry_58_port);
   U146 : XNOR2_X1 port map( A => A(60), B => B(60), ZN => n66);
   U147 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => n100);
   U148 : INV_X1 port map( A => A(43), ZN => n121);
   U149 : XNOR2_X1 port map( A => n201, B => n117, ZN => SUM(42));
   U150 : OAI21_X1 port map( B1 => B(49), B2 => n228, A => A(49), ZN => n143);
   U151 : NAND2_X1 port map( A1 => B(53), A2 => n217, ZN => n159);
   U152 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => n127);
   U153 : XNOR2_X1 port map( A => n204, B => n109, ZN => SUM(39));
   U154 : INV_X1 port map( A => A(35), ZN => n94);
   U155 : NOR2_X1 port map( A1 => B(52), A2 => n27, ZN => n153);
   U156 : OAI21_X1 port map( B1 => n153, B2 => n154, A => n155, ZN => n152);
   U157 : OAI21_X1 port map( B1 => n233, B2 => n154, A => n155, ZN => n216);
   U158 : OAI21_X1 port map( B1 => n233, B2 => n154, A => n155, ZN => n217);
   U159 : NOR2_X1 port map( A1 => B(55), A2 => n160, ZN => n163);
   U160 : OAI21_X1 port map( B1 => n163, B2 => n164, A => n165, ZN => n218);
   U161 : OAI21_X1 port map( B1 => n163, B2 => n164, A => n165, ZN => n219);
   U162 : NOR2_X1 port map( A1 => B(47), A2 => n236, ZN => n134);
   U163 : OAI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n133);
   U164 : OAI21_X1 port map( B1 => n235, B2 => n135, A => n136, ZN => n220);
   U165 : OAI21_X1 port map( B1 => n235, B2 => n135, A => n136, ZN => n221);
   U166 : NOR2_X1 port map( A1 => B(39), A2 => n103, ZN => n108);
   U167 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n107);
   U168 : OAI21_X1 port map( B1 => n237, B2 => n109, A => n110, ZN => n222);
   U169 : OAI21_X1 port map( B1 => n58, B2 => n80, A => n81, ZN => n78);
   U170 : NAND2_X1 port map( A1 => B(32), A2 => n223, ZN => n84);
   U171 : XNOR2_X1 port map( A => n223, B => B(32), ZN => n211);
   U172 : NOR2_X1 port map( A1 => n74, A2 => B(31), ZN => n79);
   U173 : OAI21_X1 port map( B1 => n80, B2 => n79, A => n81, ZN => n223);
   U174 : OAI21_X1 port map( B1 => n182, B2 => n183, A => n185, ZN => n184);
   U175 : NAND2_X1 port map( A1 => B(57), A2 => n224, ZN => n168);
   U176 : XNOR2_X1 port map( A => B(57), B => n184, ZN => n186);
   U177 : NOR2_X1 port map( A1 => B(57), A2 => n224, ZN => n167);
   U178 : NOR2_X1 port map( A1 => B(56), A2 => n219, ZN => n182);
   U179 : OAI21_X1 port map( B1 => n182, B2 => n183, A => n185, ZN => n224);
   U180 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => n119);
   U181 : NAND2_X1 port map( A1 => B(44), A2 => n119, ZN => n126);
   U182 : XNOR2_X1 port map( A => B(44), B => n225, ZN => n199);
   U183 : NOR2_X1 port map( A1 => n119, A2 => B(44), ZN => n124);
   U184 : NOR2_X1 port map( A1 => B(43), A2 => n115, ZN => n120);
   U185 : OAI21_X1 port map( B1 => n121, B2 => n120, A => n122, ZN => n225);
   U186 : OAI21_X1 port map( B1 => n64, B2 => n94, A => n95, ZN => n92);
   U187 : NAND2_X1 port map( A1 => B(36), A2 => n226, ZN => n99);
   U188 : XNOR2_X1 port map( A => n226, B => B(36), ZN => n207);
   U189 : NOR2_X1 port map( A1 => B(36), A2 => n92, ZN => n97);
   U190 : NOR2_X1 port map( A1 => B(35), A2 => n88, ZN => n93);
   U191 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n226);
   U192 : NOR2_X1 port map( A1 => B(53), A2 => n152, ZN => n157);
   U193 : OAI21_X1 port map( B1 => n157, B2 => n158, A => n159, ZN => n156);
   U194 : OAI21_X1 port map( B1 => n157, B2 => n158, A => n159, ZN => n227);
   U195 : NOR2_X1 port map( A1 => B(48), A2 => n133, ZN => n138);
   U196 : OAI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n137);
   U197 : OAI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n228);
   U198 : OAI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n123);
   U199 : NAND2_X1 port map( A1 => n229, A2 => B(45), ZN => n128);
   U200 : OAI21_X1 port map( B1 => B(45), B2 => n123, A => A(45), ZN => n129);
   U201 : XNOR2_X1 port map( A => n229, B => B(45), ZN => n198);
   U202 : OAI21_X1 port map( B1 => n125, B2 => n124, A => n126, ZN => n229);
   U203 : OAI21_X1 port map( B1 => n63, B2 => n61, A => n112, ZN => n111);
   U204 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n96);
   U205 : NAND2_X1 port map( A1 => n242, A2 => B(37), ZN => n101);
   U206 : OAI21_X1 port map( B1 => B(37), B2 => n96, A => A(37), ZN => n102);
   U207 : XNOR2_X1 port map( A => n242, B => B(37), ZN => n206);
   U208 : OAI21_X1 port map( B1 => n16, B2 => n83, A => n84, ZN => n82);
   U209 : NAND2_X1 port map( A1 => B(33), A2 => n230, ZN => n86);
   U210 : OAI21_X1 port map( B1 => B(33), B2 => n230, A => A(33), ZN => n87);
   U211 : XNOR2_X1 port map( A => B(33), B => n82, ZN => n210);
   U212 : OAI21_X1 port map( B1 => n16, B2 => n83, A => n84, ZN => n230);
   U213 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n144);
   U214 : XNOR2_X1 port map( A => n231, B => n180, ZN => n192);
   U215 : NAND2_X1 port map( A1 => B(51), A2 => n144, ZN => n151);
   U216 : NOR2_X1 port map( A1 => B(51), A2 => n144, ZN => n149);
   U217 : NOR2_X1 port map( A1 => B(50), A2 => n141, ZN => n145);
   U218 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n231);
   U219 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n70);
   U220 : XNOR2_X1 port map( A => n70, B => n170, ZN => n213);
   U221 : NAND2_X1 port map( A1 => B(30), A2 => n232, ZN => n77);
   U222 : NOR2_X1 port map( A1 => B(30), A2 => n232, ZN => n75);
   U223 : OAI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n232);
   U224 : NOR2_X1 port map( A1 => n27, A2 => B(52), ZN => n233);
   U225 : OAI21_X1 port map( B1 => n26, B2 => n150, A => n151, ZN => n148);
   U226 : NAND2_X1 port map( A1 => n148, A2 => B(52), ZN => n155);
   U227 : XNOR2_X1 port map( A => n234, B => B(52), ZN => n191);
   U228 : OAI21_X1 port map( B1 => n26, B2 => n150, A => n151, ZN => n234);
   U229 : NOR2_X1 port map( A1 => n130, A2 => B(47), ZN => n235);
   U230 : OAI21_X1 port map( B1 => n131, B2 => n49, A => n132, ZN => n130);
   U231 : XNOR2_X1 port map( A => n236, B => n178, ZN => n196);
   U232 : NAND2_X1 port map( A1 => n130, A2 => B(47), ZN => n136);
   U233 : NOR2_X1 port map( A1 => B(46), A2 => n127, ZN => n131);
   U234 : OAI21_X1 port map( B1 => n131, B2 => n49, A => n132, ZN => n236);
   U235 : NOR2_X1 port map( A1 => n238, A2 => B(39), ZN => n237);
   U236 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n103);
   U237 : XNOR2_X1 port map( A => n103, B => n174, ZN => n204);
   U238 : NAND2_X1 port map( A1 => n238, A2 => B(39), ZN => n110);
   U239 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n238);
   U240 : NAND2_X1 port map( A1 => B(56), A2 => n219, ZN => n185);
   U241 : XNOR2_X1 port map( A => B(56), B => n218, ZN => n187);
   U242 : XNOR2_X1 port map( A => B(53), B => n216, ZN => n190);
   U243 : XNOR2_X1 port map( A => A(57), B => n186, ZN => SUM(57));
   U244 : XNOR2_X1 port map( A => n191, B => n40, ZN => SUM(52));
   U245 : XNOR2_X1 port map( A => B(48), B => n220, ZN => n195);
   U246 : XNOR2_X1 port map( A => B(54), B => n227, ZN => n189);
   U247 : NAND2_X1 port map( A1 => B(54), A2 => n227, ZN => n161);
   U248 : XNOR2_X1 port map( A => n190, B => n48, ZN => SUM(53));
   U249 : NAND2_X1 port map( A1 => B(48), A2 => n221, ZN => n140);
   U250 : XNOR2_X1 port map( A => B(49), B => n137, ZN => n194);
   U251 : NAND2_X1 port map( A1 => B(49), A2 => n228, ZN => n142);
   U252 : XNOR2_X1 port map( A => A(56), B => n187, ZN => SUM(56));
   U253 : OAI21_X1 port map( B1 => n117, B2 => n116, A => n118, ZN => n115);
   U254 : XNOR2_X1 port map( A => n239, B => n176, ZN => n200);
   U255 : NAND2_X1 port map( A1 => B(43), A2 => n17, ZN => n122);
   U256 : OAI21_X1 port map( B1 => n117, B2 => n116, A => n118, ZN => n239);
   U257 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n88);
   U258 : XNOR2_X1 port map( A => n240, B => n173, ZN => n208);
   U259 : NAND2_X1 port map( A1 => B(35), A2 => n88, ZN => n95);
   U260 : NOR2_X1 port map( A1 => B(34), A2 => n85, ZN => n89);
   U261 : OAI21_X1 port map( B1 => n56, B2 => n90, A => n91, ZN => n240);
   U262 : OAI21_X1 port map( B1 => n59, B2 => n76, A => n77, ZN => n74);
   U263 : XNOR2_X1 port map( A => n241, B => n171, ZN => n212);
   U264 : NAND2_X1 port map( A1 => n241, A2 => B(31), ZN => n81);
   U265 : NAND2_X1 port map( A1 => B(40), A2 => n222, ZN => n112);
   U266 : XNOR2_X1 port map( A => n60, B => B(41), ZN => n202);
   U267 : NAND2_X1 port map( A1 => B(41), A2 => n60, ZN => n113);
   U268 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => n241);
   U269 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n68);
   U270 : OAI21_X1 port map( B1 => A(28), B2 => B(28), A => carry_28_port, ZN 
                           => n69);
   U271 : XNOR2_X1 port map( A => n215, B => A(28), ZN => SUM(28));
   U272 : XNOR2_X1 port map( A => A(33), B => n210, ZN => SUM(33));
   U273 : XNOR2_X1 port map( A => A(48), B => n195, ZN => SUM(48));
   U274 : XNOR2_X1 port map( A => B(40), B => n222, ZN => n203);
   U275 : XNOR2_X1 port map( A => A(32), B => n211, ZN => SUM(32));
   U276 : XNOR2_X1 port map( A => n206, B => n41, ZN => SUM(37));
   U277 : NAND2_X1 port map( A1 => n69, A2 => n68, ZN => n67);
   U278 : XNOR2_X1 port map( A => n67, B => n169, ZN => n214);
   U279 : NAND2_X1 port map( A1 => B(29), A2 => n67, ZN => n73);
   U280 : XNOR2_X1 port map( A => carry_28_port, B => B(28), ZN => n215);
   U281 : OAI21_X1 port map( B1 => n111, B2 => B(41), A => A(41), ZN => n114);
   U282 : XNOR2_X1 port map( A => n202, B => A(41), ZN => SUM(41));
   U283 : INV_X1 port map( A => A(32), ZN => n83);
   U284 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => n85);
   U285 : XNOR2_X1 port map( A => n51, B => n172, ZN => n209);
   U286 : NAND2_X1 port map( A1 => B(34), A2 => n85, ZN => n91);
   U287 : XNOR2_X1 port map( A => A(36), B => n207, ZN => SUM(36));
   U288 : INV_X1 port map( A => A(34), ZN => n90);
   U289 : INV_X1 port map( A => A(31), ZN => n80);
   U290 : XNOR2_X1 port map( A => n198, B => A(45), ZN => SUM(45));
   U291 : XNOR2_X1 port map( A => A(49), B => n194, ZN => SUM(49));
   U292 : XNOR2_X1 port map( A => n199, B => n62, ZN => SUM(44));
   U293 : XNOR2_X1 port map( A => n189, B => A(54), ZN => SUM(54));
   U294 : INV_X1 port map( A => A(42), ZN => n117);
   U295 : INV_X1 port map( A => A(36), ZN => n98);
   U296 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n242);
   U297 : INV_X1 port map( A => A(38), ZN => n105);
   U298 : INV_X1 port map( A => A(30), ZN => n76);
   U299 : NAND2_X1 port map( A1 => B(42), A2 => n57, ZN => n118);
   U300 : INV_X1 port map( A => A(29), ZN => n72);
   U301 : XNOR2_X1 port map( A => n203, B => n65, ZN => SUM(40));
   U302 : XNOR2_X1 port map( A => n209, B => n90, ZN => SUM(34));
   U303 : XNOR2_X1 port map( A => n100, B => n15, ZN => n205);
   U304 : XNOR2_X1 port map( A => n205, B => n105, ZN => SUM(38));
   U305 : NAND2_X1 port map( A1 => n142, A2 => n143, ZN => n141);
   U306 : XNOR2_X1 port map( A => n141, B => n179, ZN => n193);
   U307 : CLKBUF_X1 port map( A => carry_59_port, Z => net70461);
   U308 : XNOR2_X1 port map( A => net70461, B => n243, ZN => SUM(59));
   U309 : XNOR2_X1 port map( A => A(59), B => B(59), ZN => n243);
   U310 : NAND3_X1 port map( A1 => n245, A2 => n246, A3 => n247, ZN => n244);
   U311 : NAND2_X1 port map( A1 => carry_59_port, A2 => A(59), ZN => n245);
   U312 : NAND2_X1 port map( A1 => carry_59_port, A2 => B(59), ZN => n246);
   U313 : NAND2_X1 port map( A1 => A(59), A2 => B(59), ZN => n247);
   U314 : NAND3_X1 port map( A1 => n246, A2 => n245, A3 => n247, ZN => 
                           carry_60_port);
   U315 : NAND2_X1 port map( A1 => n244, A2 => A(60), ZN => n248);
   U316 : NAND2_X1 port map( A1 => carry_60_port, A2 => B(60), ZN => n249);
   U317 : NAND2_X1 port map( A1 => A(60), A2 => B(60), ZN => n250);
   U318 : NAND3_X1 port map( A1 => n248, A2 => n249, A3 => n250, ZN => 
                           carry_61_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_13_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_13_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_13_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , net18124, carry_45_port, carry_44_port, net29754, net29753, net29752, 
      carry_43_port, carry_42_port, carry_41_port, carry_40_port, carry_39_port
      , carry_38_port, carry_37_port, carry_36_port, carry_35_port, 
      carry_34_port, carry_33_port, carry_32_port, carry_31_port, carry_30_port
      , carry_29_port, carry_28_port, carry_27_port, carry_26_port, 
      carry_25_port, carry_24_port, carry_23_port, carry_22_port, carry_21_port
      , carry_20_port, carry_19_port, carry_18_port, carry_17_port, 
      carry_16_port, carry_15_port, carry_14_port, carry_13_port, net84281, 
      net84280, net89911, net89905, net89896, net89886, net89863, net89850, 
      net89849, net89825, net89823, net90207, net90206, net93331, net89932, 
      net89927, net89922, net93330, net90245, net90234, net90233, net90229, 
      net90223, net90221, net90202, net89919, net89908, net89865, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => B(13), B => A(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1 : BUF_X1 port map( A => A(23), Z => n2);
   U2 : BUF_X1 port map( A => A(34), Z => n1);
   U3 : BUF_X1 port map( A => A(43), Z => n3);
   U4 : BUF_X1 port map( A => A(32), Z => n4);
   U5 : XNOR2_X1 port map( A => n5, B => net29752, ZN => SUM(43));
   U6 : AND3_X1 port map( A1 => n165, A2 => n164, A3 => n166, ZN => n5);
   U7 : AND2_X1 port map( A1 => net90202, A2 => n26, ZN => n6);
   U8 : CLKBUF_X1 port map( A => net89905, Z => n33);
   U9 : BUF_X1 port map( A => A(7), Z => n25);
   U10 : NAND3_X1 port map( A1 => n131, A2 => n130, A3 => n132, ZN => n7);
   U11 : CLKBUF_X1 port map( A => carry_15_port, Z => n8);
   U12 : NAND3_X1 port map( A1 => n155, A2 => n154, A3 => n153, ZN => n9);
   U13 : NAND3_X1 port map( A1 => n199, A2 => n200, A3 => n201, ZN => n10);
   U14 : NAND3_X1 port map( A1 => n184, A2 => n185, A3 => n186, ZN => n11);
   U15 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => n12);
   U16 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => n13);
   U17 : XOR2_X1 port map( A => A(31), B => B(31), Z => n14);
   U18 : XOR2_X1 port map( A => carry_31_port, B => n14, Z => SUM(31));
   U19 : NAND2_X1 port map( A1 => carry_31_port, A2 => A(31), ZN => n15);
   U20 : NAND2_X1 port map( A1 => carry_31_port, A2 => B(31), ZN => n16);
   U21 : NAND2_X1 port map( A1 => A(31), A2 => B(31), ZN => n17);
   U22 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => n17, ZN => 
                           carry_32_port);
   U23 : XOR2_X1 port map( A => A(32), B => B(32), Z => n18);
   U24 : XOR2_X1 port map( A => carry_32_port, B => n18, Z => SUM(32));
   U25 : NAND2_X1 port map( A1 => carry_32_port, A2 => n4, ZN => n19);
   U26 : NAND2_X1 port map( A1 => carry_32_port, A2 => B(32), ZN => n20);
   U27 : NAND2_X1 port map( A1 => n4, A2 => B(32), ZN => n21);
   U28 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => 
                           carry_33_port);
   U29 : INV_X1 port map( A => B(38), ZN => n100);
   U30 : INV_X1 port map( A => B(7), ZN => net89823);
   U31 : INV_X1 port map( A => B(35), ZN => n193);
   U32 : INV_X1 port map( A => B(42), ZN => n133);
   U33 : INV_X1 port map( A => B(11), ZN => n43);
   U34 : INV_X1 port map( A => A(4), ZN => n49);
   U35 : INV_X1 port map( A => B(4), ZN => n48);
   U36 : INV_X1 port map( A => B(9), ZN => net90223);
   U37 : INV_X1 port map( A => B(43), ZN => n91);
   U38 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n64);
   U39 : OAI21_X1 port map( B1 => n76, B2 => n55, A => n77, ZN => n65);
   U40 : INV_X1 port map( A => n67, ZN => n76);
   U41 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n77);
   U42 : NOR2_X1 port map( A1 => A(2), A2 => B(2), ZN => n55);
   U43 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n62);
   U44 : OAI21_X1 port map( B1 => n78, B2 => n56, A => n79, ZN => n63);
   U45 : INV_X1 port map( A => n65, ZN => n78);
   U46 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n79);
   U47 : NOR2_X1 port map( A1 => A(3), A2 => B(3), ZN => n56);
   U48 : INV_X1 port map( A => A(6), ZN => n51);
   U49 : INV_X1 port map( A => B(6), ZN => n50);
   U50 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n60);
   U51 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n61);
   U52 : NAND2_X1 port map( A1 => n85, A2 => n63, ZN => n80);
   U53 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n81);
   U54 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => n85);
   U55 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n58);
   U56 : OAI21_X1 port map( B1 => n82, B2 => n57, A => n83, ZN => n59);
   U57 : INV_X1 port map( A => n61, ZN => n82);
   U58 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n83);
   U59 : NOR2_X1 port map( A1 => A(5), A2 => B(5), ZN => n57);
   U60 : INV_X1 port map( A => B(15), ZN => n124);
   U61 : INV_X1 port map( A => B(39), ZN => n128);
   U62 : INV_X1 port map( A => B(56), ZN => n192);
   U63 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n66);
   U64 : OAI21_X1 port map( B1 => n74, B2 => n54, A => n75, ZN => n67);
   U65 : INV_X1 port map( A => n69, ZN => n74);
   U66 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n75);
   U67 : NOR2_X1 port map( A1 => A(1), A2 => B(1), ZN => n54);
   U68 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n68);
   U69 : NAND2_X1 port map( A1 => B(0), A2 => CI, ZN => n73);
   U70 : NAND2_X1 port map( A1 => A(0), A2 => CI, ZN => n72);
   U71 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n71);
   U72 : XNOR2_X1 port map( A => n64, B => n65, ZN => SUM(3));
   U73 : XNOR2_X1 port map( A => n62, B => n63, ZN => SUM(4));
   U74 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => net18124);
   U75 : NAND2_X1 port map( A1 => n86, A2 => n59, ZN => n52);
   U76 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n53);
   U77 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => n86);
   U78 : XNOR2_X1 port map( A => n60, B => n61, ZN => SUM(5));
   U79 : XNOR2_X1 port map( A => n58, B => n59, ZN => SUM(6));
   U80 : INV_X1 port map( A => B(48), ZN => n167);
   U81 : XNOR2_X1 port map( A => B(0), B => CI, ZN => n70);
   U82 : XNOR2_X1 port map( A => n66, B => n67, ZN => SUM(2));
   U83 : XNOR2_X1 port map( A => n68, B => n69, ZN => SUM(1));
   U84 : XNOR2_X1 port map( A => A(0), B => n70, ZN => SUM(0));
   U85 : XOR2_X1 port map( A => B(7), B => n25, Z => n22);
   U86 : NAND2_X1 port map( A1 => net90202, A2 => n26, ZN => net89908);
   U87 : XNOR2_X1 port map( A => carry_28_port, B => n23, ZN => SUM(28));
   U88 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n23);
   U89 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => net89865);
   U90 : XNOR2_X1 port map( A => net89865, B => net89908, ZN => SUM(10));
   U91 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => net90206);
   U92 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => net90207);
   U93 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => n26);
   U94 : NAND3_X1 port map( A1 => net90234, A2 => net90229, A3 => net90233, ZN 
                           => n27);
   U95 : NAND2_X1 port map( A1 => net89927, A2 => B(8), ZN => net90233);
   U96 : INV_X1 port map( A => net89919, ZN => net90229);
   U97 : NAND2_X1 port map( A1 => n30, A2 => net89850, ZN => net90234);
   U98 : NAND2_X1 port map( A1 => B(7), A2 => n25, ZN => n24);
   U99 : NAND2_X1 port map( A1 => B(7), A2 => n25, ZN => net89932);
   U100 : CLKBUF_X1 port map( A => A(8), Z => n30);
   U101 : NAND2_X1 port map( A1 => net90221, A2 => net90223, ZN => n28);
   U102 : INV_X1 port map( A => A(9), ZN => net90221);
   U103 : INV_X1 port map( A => net90221, ZN => net90245);
   U104 : NAND2_X1 port map( A1 => B(9), A2 => net90245, ZN => net90202);
   U105 : AOI21_X1 port map( B1 => net89927, B2 => n29, A => net89919, ZN => 
                           net89922);
   U106 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => net89849);
   U107 : AND2_X1 port map( A1 => A(8), A2 => B(8), ZN => net89919);
   U108 : OR2_X1 port map( A1 => A(8), A2 => B(8), ZN => n29);
   U109 : NAND2_X1 port map( A1 => net89896, A2 => n24, ZN => net89850);
   U110 : INV_X1 port map( A => A(7), ZN => net89825);
   U111 : XNOR2_X1 port map( A => A(9), B => B(9), ZN => net93330);
   U112 : NAND2_X1 port map( A1 => n84, A2 => net18124, ZN => net89896);
   U113 : XNOR2_X1 port map( A => net93330, B => net93331, ZN => SUM(9));
   U114 : INV_X1 port map( A => net89922, ZN => net93331);
   U115 : NAND2_X1 port map( A1 => net89886, A2 => net89932, ZN => net89927);
   U116 : CLKBUF_X1 port map( A => A(41), Z => n31);
   U117 : CLKBUF_X1 port map( A => n45, Z => n32);
   U118 : BUF_X1 port map( A => A(25), Z => n34);
   U119 : NAND2_X1 port map( A1 => carry_28_port, A2 => A(28), ZN => n35);
   U120 : NAND2_X1 port map( A1 => carry_28_port, A2 => B(28), ZN => n36);
   U121 : NAND2_X1 port map( A1 => A(28), A2 => B(28), ZN => n37);
   U122 : NAND3_X1 port map( A1 => n35, A2 => n36, A3 => n37, ZN => 
                           carry_29_port);
   U123 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => n38);
   U124 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => n39);
   U125 : NAND3_X1 port map( A1 => n149, A2 => n150, A3 => n151, ZN => n40);
   U126 : NAND2_X1 port map( A1 => n41, A2 => B(12), ZN => net84281);
   U127 : OAI21_X1 port map( B1 => n6, B2 => net90206, A => net90207, ZN => 
                           net89911);
   U128 : OAI21_X1 port map( B1 => n6, B2 => net90206, A => net90207, ZN => n45
                           );
   U129 : OAI21_X1 port map( B1 => n46, B2 => n43, A => n44, ZN => n41);
   U130 : NOR2_X1 port map( A1 => net89911, A2 => A(11), ZN => n42);
   U131 : OAI21_X1 port map( B1 => n42, B2 => n43, A => n44, ZN => net89905);
   U132 : NOR2_X1 port map( A1 => net89911, A2 => A(11), ZN => n46);
   U133 : NAND2_X1 port map( A1 => A(11), A2 => n45, ZN => n44);
   U134 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => net89863);
   U135 : XNOR2_X1 port map( A => n47, B => n90, ZN => SUM(18));
   U136 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n47);
   U137 : NAND3_X1 port map( A1 => n72, A2 => n71, A3 => n73, ZN => n69);
   U138 : NAND2_X1 port map( A1 => A(12), A2 => net89905, ZN => net84280);
   U139 : NAND2_X1 port map( A1 => n84, A2 => net18124, ZN => net89886);
   U140 : NAND2_X1 port map( A1 => net89825, A2 => net89823, ZN => n84);
   U141 : XNOR2_X1 port map( A => net89849, B => net89850, ZN => SUM(8));
   U142 : XNOR2_X1 port map( A => net89863, B => n32, ZN => SUM(11));
   U143 : CLKBUF_X1 port map( A => A(35), Z => n87);
   U144 : XNOR2_X1 port map( A => n94, B => n88, ZN => SUM(19));
   U145 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n88);
   U146 : NAND3_X1 port map( A1 => n180, A2 => n181, A3 => n182, ZN => n89);
   U147 : CLKBUF_X1 port map( A => carry_18_port, Z => n90);
   U148 : XNOR2_X1 port map( A => A(43), B => n91, ZN => net29752);
   U149 : CLKBUF_X1 port map( A => carry_29_port, Z => n92);
   U150 : NAND3_X1 port map( A1 => n106, A2 => n107, A3 => n108, ZN => n93);
   U151 : CLKBUF_X1 port map( A => n89, Z => n94);
   U152 : NAND3_X1 port map( A1 => n104, A2 => n103, A3 => n102, ZN => n95);
   U153 : NAND3_X1 port map( A1 => n102, A2 => n103, A3 => n104, ZN => n96);
   U154 : NAND3_X1 port map( A1 => n157, A2 => n158, A3 => n159, ZN => n97);
   U155 : XNOR2_X1 port map( A => n98, B => n33, ZN => SUM(12));
   U156 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n98);
   U157 : XNOR2_X1 port map( A => n99, B => n97, ZN => SUM(26));
   U158 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n99);
   U159 : XNOR2_X1 port map( A => A(38), B => n100, ZN => n152);
   U160 : XOR2_X1 port map( A => A(33), B => B(33), Z => n101);
   U161 : XOR2_X1 port map( A => n101, B => n13, Z => SUM(33));
   U162 : NAND2_X1 port map( A1 => A(33), A2 => B(33), ZN => n102);
   U163 : NAND2_X1 port map( A1 => A(33), A2 => carry_33_port, ZN => n103);
   U164 : NAND2_X1 port map( A1 => B(33), A2 => n12, ZN => n104);
   U165 : NAND3_X1 port map( A1 => n102, A2 => n103, A3 => n104, ZN => 
                           carry_34_port);
   U166 : XOR2_X1 port map( A => A(34), B => B(34), Z => n105);
   U167 : XOR2_X1 port map( A => n105, B => n96, Z => SUM(34));
   U168 : NAND2_X1 port map( A1 => n1, A2 => B(34), ZN => n106);
   U169 : NAND2_X1 port map( A1 => n1, A2 => n95, ZN => n107);
   U170 : NAND2_X1 port map( A1 => B(34), A2 => carry_34_port, ZN => n108);
   U171 : NAND3_X1 port map( A1 => n106, A2 => n107, A3 => n108, ZN => 
                           carry_35_port);
   U172 : XOR2_X1 port map( A => A(23), B => B(23), Z => n109);
   U173 : XOR2_X1 port map( A => carry_23_port, B => n109, Z => SUM(23));
   U174 : NAND2_X1 port map( A1 => carry_23_port, A2 => n2, ZN => n110);
   U175 : NAND2_X1 port map( A1 => carry_23_port, A2 => B(23), ZN => n111);
   U176 : NAND2_X1 port map( A1 => n2, A2 => B(23), ZN => n112);
   U177 : NAND3_X1 port map( A1 => n110, A2 => n111, A3 => n112, ZN => 
                           carry_24_port);
   U178 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n113);
   U179 : NAND3_X1 port map( A1 => net84280, A2 => net84281, A3 => n113, ZN => 
                           carry_13_port);
   U180 : XOR2_X1 port map( A => A(36), B => B(36), Z => n114);
   U181 : XOR2_X1 port map( A => carry_36_port, B => n114, Z => SUM(36));
   U182 : NAND2_X1 port map( A1 => n10, A2 => A(36), ZN => n115);
   U183 : NAND2_X1 port map( A1 => carry_36_port, A2 => B(36), ZN => n116);
   U184 : NAND2_X1 port map( A1 => A(36), A2 => B(36), ZN => n117);
   U185 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => 
                           carry_37_port);
   U186 : CLKBUF_X1 port map( A => A(26), Z => n123);
   U187 : XOR2_X1 port map( A => A(55), B => B(55), Z => n118);
   U188 : XOR2_X1 port map( A => carry_55_port, B => n118, Z => SUM(55));
   U189 : NAND2_X1 port map( A1 => carry_55_port, A2 => A(55), ZN => n119);
   U190 : NAND2_X1 port map( A1 => carry_55_port, A2 => B(55), ZN => n120);
   U191 : NAND2_X1 port map( A1 => A(55), A2 => B(55), ZN => n121);
   U192 : NAND3_X1 port map( A1 => n119, A2 => n120, A3 => n121, ZN => 
                           carry_56_port);
   U193 : NAND3_X1 port map( A1 => n196, A2 => n195, A3 => n197, ZN => n122);
   U194 : XNOR2_X1 port map( A => A(15), B => n124, ZN => n129);
   U195 : XNOR2_X1 port map( A => n127, B => n125, ZN => SUM(16));
   U196 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n125);
   U197 : NAND3_X1 port map( A1 => n146, A2 => n145, A3 => n147, ZN => n126);
   U198 : CLKBUF_X1 port map( A => n7, Z => n127);
   U199 : XNOR2_X1 port map( A => A(39), B => n128, ZN => n134);
   U200 : XOR2_X1 port map( A => n129, B => n8, Z => SUM(15));
   U201 : NAND2_X1 port map( A1 => carry_15_port, A2 => A(15), ZN => n130);
   U202 : NAND2_X1 port map( A1 => carry_15_port, A2 => B(15), ZN => n131);
   U203 : NAND2_X1 port map( A1 => A(15), A2 => B(15), ZN => n132);
   U204 : NAND3_X1 port map( A1 => n131, A2 => n130, A3 => n132, ZN => 
                           carry_16_port);
   U205 : XNOR2_X1 port map( A => A(42), B => n133, ZN => n163);
   U206 : XOR2_X1 port map( A => carry_39_port, B => n134, Z => SUM(39));
   U207 : NAND2_X1 port map( A1 => carry_39_port, A2 => A(39), ZN => n135);
   U208 : NAND2_X1 port map( A1 => n9, A2 => B(39), ZN => n136);
   U209 : NAND2_X1 port map( A1 => A(39), A2 => B(39), ZN => n137);
   U210 : NAND3_X1 port map( A1 => n136, A2 => n135, A3 => n137, ZN => 
                           carry_40_port);
   U211 : NAND2_X1 port map( A1 => n7, A2 => A(16), ZN => n138);
   U212 : NAND2_X1 port map( A1 => carry_16_port, A2 => B(16), ZN => n139);
   U213 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => n140);
   U214 : NAND3_X1 port map( A1 => n138, A2 => n139, A3 => n140, ZN => 
                           carry_17_port);
   U215 : NAND2_X1 port map( A1 => n89, A2 => A(19), ZN => n141);
   U216 : NAND2_X1 port map( A1 => carry_19_port, A2 => B(19), ZN => n142);
   U217 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n143);
   U218 : NAND3_X1 port map( A1 => n141, A2 => n142, A3 => n143, ZN => 
                           carry_20_port);
   U219 : XOR2_X1 port map( A => A(41), B => B(41), Z => n144);
   U220 : XOR2_X1 port map( A => carry_41_port, B => n144, Z => SUM(41));
   U221 : NAND2_X1 port map( A1 => carry_41_port, A2 => n31, ZN => n145);
   U222 : NAND2_X1 port map( A1 => carry_41_port, A2 => B(41), ZN => n146);
   U223 : NAND2_X1 port map( A1 => n31, A2 => B(41), ZN => n147);
   U224 : NAND3_X1 port map( A1 => n145, A2 => n146, A3 => n147, ZN => 
                           carry_42_port);
   U225 : XOR2_X1 port map( A => A(37), B => B(37), Z => n148);
   U226 : XOR2_X1 port map( A => n148, B => n39, Z => SUM(37));
   U227 : NAND2_X1 port map( A1 => A(37), A2 => B(37), ZN => n149);
   U228 : NAND2_X1 port map( A1 => A(37), A2 => n38, ZN => n150);
   U229 : NAND2_X1 port map( A1 => B(37), A2 => carry_37_port, ZN => n151);
   U230 : NAND3_X1 port map( A1 => n149, A2 => n150, A3 => n151, ZN => 
                           carry_38_port);
   U231 : XOR2_X1 port map( A => n152, B => carry_38_port, Z => SUM(38));
   U232 : NAND2_X1 port map( A1 => A(38), A2 => B(38), ZN => n153);
   U233 : NAND2_X1 port map( A1 => A(38), A2 => n40, ZN => n154);
   U234 : NAND2_X1 port map( A1 => B(38), A2 => carry_38_port, ZN => n155);
   U235 : NAND3_X1 port map( A1 => n155, A2 => n154, A3 => n153, ZN => 
                           carry_39_port);
   U236 : XOR2_X1 port map( A => A(25), B => B(25), Z => n156);
   U237 : XOR2_X1 port map( A => n156, B => carry_25_port, Z => SUM(25));
   U238 : NAND2_X1 port map( A1 => n34, A2 => B(25), ZN => n157);
   U239 : NAND2_X1 port map( A1 => n34, A2 => carry_25_port, ZN => n158);
   U240 : NAND2_X1 port map( A1 => B(25), A2 => carry_25_port, ZN => n159);
   U241 : NAND3_X1 port map( A1 => n159, A2 => n158, A3 => n157, ZN => 
                           carry_26_port);
   U242 : NAND2_X1 port map( A1 => n123, A2 => B(26), ZN => n160);
   U243 : NAND2_X1 port map( A1 => n123, A2 => n97, ZN => n161);
   U244 : NAND2_X1 port map( A1 => B(26), A2 => carry_26_port, ZN => n162);
   U245 : NAND3_X1 port map( A1 => n160, A2 => n161, A3 => n162, ZN => 
                           carry_27_port);
   U246 : XOR2_X1 port map( A => carry_42_port, B => n163, Z => SUM(42));
   U247 : NAND2_X1 port map( A1 => A(42), A2 => n126, ZN => n164);
   U248 : NAND2_X1 port map( A1 => carry_42_port, A2 => B(42), ZN => n165);
   U249 : NAND2_X1 port map( A1 => A(42), A2 => B(42), ZN => n166);
   U250 : NAND3_X1 port map( A1 => n165, A2 => n164, A3 => n166, ZN => 
                           carry_43_port);
   U251 : XNOR2_X1 port map( A => A(48), B => n167, ZN => n168);
   U252 : XOR2_X1 port map( A => carry_48_port, B => n168, Z => SUM(48));
   U253 : NAND2_X1 port map( A1 => carry_48_port, A2 => A(48), ZN => n169);
   U254 : NAND2_X1 port map( A1 => carry_48_port, A2 => B(48), ZN => n170);
   U255 : NAND2_X1 port map( A1 => A(48), A2 => B(48), ZN => n171);
   U256 : NAND3_X1 port map( A1 => n169, A2 => n170, A3 => n171, ZN => 
                           carry_49_port);
   U257 : XOR2_X1 port map( A => A(57), B => B(57), Z => n172);
   U258 : XOR2_X1 port map( A => carry_57_port, B => n172, Z => SUM(57));
   U259 : NAND2_X1 port map( A1 => n122, A2 => A(57), ZN => n173);
   U260 : NAND2_X1 port map( A1 => carry_57_port, A2 => B(57), ZN => n174);
   U261 : NAND2_X1 port map( A1 => A(57), A2 => B(57), ZN => n175);
   U262 : NAND3_X1 port map( A1 => n173, A2 => n174, A3 => n175, ZN => 
                           carry_58_port);
   U263 : XOR2_X1 port map( A => A(52), B => B(52), Z => n176);
   U264 : XOR2_X1 port map( A => carry_52_port, B => n176, Z => SUM(52));
   U265 : NAND2_X1 port map( A1 => carry_52_port, A2 => A(52), ZN => n177);
   U266 : NAND2_X1 port map( A1 => carry_52_port, A2 => B(52), ZN => n178);
   U267 : NAND2_X1 port map( A1 => A(52), A2 => B(52), ZN => n179);
   U268 : NAND3_X1 port map( A1 => n177, A2 => n178, A3 => n179, ZN => 
                           carry_53_port);
   U269 : NAND2_X1 port map( A1 => carry_18_port, A2 => A(18), ZN => n180);
   U270 : NAND2_X1 port map( A1 => carry_18_port, A2 => B(18), ZN => n181);
   U271 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n182);
   U272 : NAND3_X1 port map( A1 => n181, A2 => n180, A3 => n182, ZN => 
                           carry_19_port);
   U273 : XOR2_X1 port map( A => A(29), B => B(29), Z => n183);
   U274 : XOR2_X1 port map( A => n92, B => n183, Z => SUM(29));
   U275 : NAND2_X1 port map( A1 => carry_29_port, A2 => A(29), ZN => n184);
   U276 : NAND2_X1 port map( A1 => carry_29_port, A2 => B(29), ZN => n185);
   U277 : NAND2_X1 port map( A1 => A(29), A2 => B(29), ZN => n186);
   U278 : NAND3_X1 port map( A1 => n184, A2 => n185, A3 => n186, ZN => 
                           carry_30_port);
   U279 : XOR2_X1 port map( A => A(30), B => B(30), Z => n187);
   U280 : XOR2_X1 port map( A => carry_30_port, B => n187, Z => SUM(30));
   U281 : NAND2_X1 port map( A1 => n11, A2 => A(30), ZN => n188);
   U282 : NAND2_X1 port map( A1 => carry_30_port, A2 => B(30), ZN => n189);
   U283 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n190);
   U284 : NAND3_X1 port map( A1 => n188, A2 => n189, A3 => n190, ZN => 
                           carry_31_port);
   U285 : CLKBUF_X1 port map( A => carry_56_port, Z => n191);
   U286 : XNOR2_X1 port map( A => A(56), B => n192, ZN => n194);
   U287 : XNOR2_X1 port map( A => A(35), B => n193, ZN => n198);
   U288 : XOR2_X1 port map( A => n191, B => n194, Z => SUM(56));
   U289 : NAND2_X1 port map( A1 => carry_56_port, A2 => A(56), ZN => n195);
   U290 : NAND2_X1 port map( A1 => carry_56_port, A2 => B(56), ZN => n196);
   U291 : NAND2_X1 port map( A1 => A(56), A2 => B(56), ZN => n197);
   U292 : NAND3_X1 port map( A1 => n196, A2 => n195, A3 => n197, ZN => 
                           carry_57_port);
   U293 : XOR2_X1 port map( A => carry_35_port, B => n198, Z => SUM(35));
   U294 : NAND2_X1 port map( A1 => n93, A2 => n87, ZN => n199);
   U295 : NAND2_X1 port map( A1 => carry_35_port, A2 => B(35), ZN => n200);
   U296 : NAND2_X1 port map( A1 => n87, A2 => B(35), ZN => n201);
   U297 : NAND3_X1 port map( A1 => n199, A2 => n200, A3 => n201, ZN => 
                           carry_36_port);
   U298 : NAND2_X1 port map( A1 => carry_43_port, A2 => B(43), ZN => net29754);
   U299 : NAND2_X1 port map( A1 => n3, A2 => carry_43_port, ZN => net29753);
   U300 : NAND2_X1 port map( A1 => n3, A2 => B(43), ZN => n202);
   U301 : NAND3_X1 port map( A1 => net29754, A2 => net29753, A3 => n202, ZN => 
                           carry_44_port);
   U302 : XOR2_X1 port map( A => net18124, B => n22, Z => SUM(7));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_14_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_14_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_14_DW01_add_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_4_port,
      carry_3_port, carry_2_port, carry_1_port, net17921, net17991, net18132, 
      net69934, net69933, net69932, net98250, net98278, net93358, net69924, 
      net69923, net90419, net90405, net69954, net69949, net69945, net69944, 
      net69930, net69928, net69927, net17910, net25732, net18111, net17868, 
      net17867, net17866, carry_6_port, carry_5_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_20 : FA_X1 port map( A => B(20), B => A(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_14 : FA_X1 port map( A => B(14), B => A(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           net18111, S => SUM(6));
   U1 : BUF_X1 port map( A => A(25), Z => n4);
   U2 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => n12, ZN => n1);
   U3 : OAI21_X1 port map( B1 => A(7), B2 => B(7), A => net18111, ZN => n2);
   U4 : CLKBUF_X1 port map( A => A(22), Z => n3);
   U5 : CLKBUF_X1 port map( A => net18111, Z => net98278);
   U6 : BUF_X1 port map( A => A(15), Z => n50);
   U7 : CLKBUF_X1 port map( A => A(30), Z => n5);
   U8 : CLKBUF_X1 port map( A => A(34), Z => n6);
   U9 : CLKBUF_X1 port map( A => A(9), Z => n43);
   U10 : NAND2_X1 port map( A1 => net69954, A2 => B(9), ZN => n7);
   U11 : XNOR2_X1 port map( A => n8, B => carry_36_port, ZN => SUM(36));
   U12 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n8);
   U13 : XOR2_X1 port map( A => A(26), B => B(26), Z => n9);
   U14 : XOR2_X1 port map( A => carry_26_port, B => n9, Z => SUM(26));
   U15 : NAND2_X1 port map( A1 => carry_26_port, A2 => A(26), ZN => n10);
   U16 : NAND2_X1 port map( A1 => carry_26_port, A2 => B(26), ZN => n11);
   U17 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n12);
   U18 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => n12, ZN => 
                           carry_27_port);
   U19 : XOR2_X1 port map( A => A(31), B => B(31), Z => n13);
   U20 : XOR2_X1 port map( A => carry_31_port, B => n13, Z => SUM(31));
   U21 : NAND2_X1 port map( A1 => carry_31_port, A2 => A(31), ZN => n14);
   U22 : NAND2_X1 port map( A1 => carry_31_port, A2 => B(31), ZN => n15);
   U23 : NAND2_X1 port map( A1 => A(31), A2 => B(31), ZN => n16);
   U24 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => 
                           carry_32_port);
   U25 : XOR2_X1 port map( A => A(21), B => B(21), Z => n17);
   U26 : XOR2_X1 port map( A => carry_21_port, B => n17, Z => SUM(21));
   U27 : NAND2_X1 port map( A1 => carry_21_port, A2 => A(21), ZN => n18);
   U28 : NAND2_X1 port map( A1 => carry_21_port, A2 => B(21), ZN => n19);
   U29 : NAND2_X1 port map( A1 => A(21), A2 => B(21), ZN => n20);
   U30 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => 
                           carry_22_port);
   U31 : NAND3_X1 port map( A1 => n127, A2 => n128, A3 => n129, ZN => n21);
   U32 : NAND3_X1 port map( A1 => n152, A2 => n153, A3 => n154, ZN => n22);
   U33 : NAND3_X1 port map( A1 => n69, A2 => n68, A3 => n67, ZN => n23);
   U34 : NAND3_X1 port map( A1 => n69, A2 => n68, A3 => n67, ZN => n24);
   U35 : NAND3_X1 port map( A1 => n73, A2 => n72, A3 => n71, ZN => n25);
   U36 : NOR2_X1 port map( A1 => B(9), A2 => net69927, ZN => n26);
   U37 : XOR2_X1 port map( A => A(58), B => B(58), Z => n27);
   U38 : XOR2_X1 port map( A => carry_58_port, B => n27, Z => SUM(58));
   U39 : NAND2_X1 port map( A1 => carry_58_port, A2 => A(58), ZN => n28);
   U40 : NAND2_X1 port map( A1 => carry_58_port, A2 => B(58), ZN => n29);
   U41 : NAND2_X1 port map( A1 => A(58), A2 => B(58), ZN => n30);
   U42 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => 
                           carry_59_port);
   U43 : INV_X1 port map( A => B(48), ZN => n103);
   U44 : INV_X1 port map( A => B(23), ZN => n32);
   U45 : XNOR2_X1 port map( A => n31, B => carry_11_port, ZN => SUM(11));
   U46 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => n31);
   U47 : XNOR2_X1 port map( A => A(23), B => n32, ZN => n159);
   U48 : XNOR2_X1 port map( A => n97, B => n33, ZN => SUM(16));
   U49 : AND3_X1 port map( A1 => n96, A2 => n95, A3 => n94, ZN => n33);
   U50 : OAI21_X1 port map( B1 => net69945, B2 => n26, A => n7, ZN => net93358)
                           ;
   U51 : XOR2_X1 port map( A => n134, B => n21, Z => SUM(28));
   U52 : OAI21_X1 port map( B1 => A(7), B2 => B(7), A => net18111, ZN => 
                           net69924);
   U53 : NAND3_X1 port map( A1 => n37, A2 => n35, A3 => n36, ZN => carry_6_port
                           );
   U54 : NAND2_X1 port map( A1 => A(5), A2 => B(5), ZN => n36);
   U55 : NAND2_X1 port map( A1 => carry_5_port, A2 => B(5), ZN => n37);
   U56 : NAND3_X1 port map( A1 => net17866, A2 => net17867, A3 => net17868, ZN 
                           => carry_5_port);
   U57 : NAND2_X1 port map( A1 => n39, A2 => A(5), ZN => n35);
   U58 : NAND3_X1 port map( A1 => net17866, A2 => net17867, A3 => net17868, ZN 
                           => n39);
   U59 : CLKBUF_X1 port map( A => A(5), Z => net18132);
   U60 : XOR2_X1 port map( A => n40, B => B(5), Z => net17991);
   U61 : NAND2_X1 port map( A1 => carry_4_port, A2 => n38, ZN => net17866);
   U62 : NAND3_X1 port map( A1 => net17866, A2 => net17867, A3 => net17868, ZN 
                           => n40);
   U63 : CLKBUF_X1 port map( A => A(4), Z => n38);
   U64 : XOR2_X1 port map( A => n38, B => B(4), Z => n34);
   U65 : NAND2_X1 port map( A1 => carry_4_port, A2 => B(4), ZN => net17867);
   U66 : NAND2_X1 port map( A1 => A(4), A2 => B(4), ZN => net17868);
   U67 : XOR2_X1 port map( A => carry_4_port, B => n34, Z => SUM(4));
   U68 : NOR2_X1 port map( A1 => net25732, A2 => B(8), ZN => n41);
   U69 : OAI21_X1 port map( B1 => n41, B2 => net69928, A => net69930, ZN => 
                           net69954);
   U70 : NAND2_X1 port map( A1 => net25732, A2 => B(8), ZN => net69930);
   U71 : NOR2_X1 port map( A1 => net90405, A2 => B(8), ZN => net90419);
   U72 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => net17910);
   U73 : NAND2_X1 port map( A1 => net69924, A2 => net69923, ZN => net25732);
   U74 : NAND2_X1 port map( A1 => n2, A2 => net69923, ZN => net90405);
   U75 : OAI21_X1 port map( B1 => net69944, B2 => net69945, A => n7, ZN => n42)
                           ;
   U76 : INV_X1 port map( A => n42, ZN => net69933);
   U77 : INV_X1 port map( A => n43, ZN => net69945);
   U78 : NOR2_X1 port map( A1 => net69927, A2 => B(9), ZN => net69944);
   U79 : OAI21_X1 port map( B1 => net90419, B2 => net69928, A => net69930, ZN 
                           => net69927);
   U80 : INV_X1 port map( A => A(8), ZN => net69928);
   U81 : XNOR2_X1 port map( A => net69954, B => net69949, ZN => SUM(9));
   U82 : XNOR2_X1 port map( A => A(9), B => B(9), ZN => net69949);
   U83 : XNOR2_X1 port map( A => net17910, B => net90405, ZN => SUM(8));
   U84 : XNOR2_X1 port map( A => A(7), B => B(7), ZN => net17921);
   U85 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => net69923);
   U86 : XNOR2_X1 port map( A => n44, B => net93358, ZN => SUM(10));
   U87 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n44);
   U88 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => net69934);
   U89 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => net69932);
   U90 : CLKBUF_X1 port map( A => net69933, Z => net98250);
   U91 : BUF_X1 port map( A => carry_25_port, Z => n51);
   U92 : XNOR2_X1 port map( A => carry_13_port, B => n45, ZN => SUM(13));
   U93 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n45);
   U94 : XNOR2_X1 port map( A => n169, B => n46, ZN => SUM(17));
   U95 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n46);
   U96 : XNOR2_X1 port map( A => n52, B => n47, ZN => SUM(19));
   U97 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n47);
   U98 : AOI21_X1 port map( B1 => net69933, B2 => net69932, A => net69934, ZN 
                           => n48);
   U99 : NAND3_X1 port map( A1 => n100, A2 => n99, A3 => n98, ZN => n49);
   U100 : AOI21_X1 port map( B1 => net98250, B2 => net69932, A => net69934, ZN 
                           => carry_11_port);
   U101 : CLKBUF_X1 port map( A => carry_19_port, Z => n52);
   U102 : NAND3_X1 port map( A1 => n95, A2 => n96, A3 => n94, ZN => n53);
   U103 : XOR2_X1 port map( A => A(35), B => B(35), Z => n54);
   U104 : XOR2_X1 port map( A => n54, B => carry_35_port, Z => SUM(35));
   U105 : NAND2_X1 port map( A1 => A(35), A2 => B(35), ZN => n55);
   U106 : NAND2_X1 port map( A1 => A(35), A2 => n22, ZN => n56);
   U107 : NAND2_X1 port map( A1 => B(35), A2 => carry_35_port, ZN => n57);
   U108 : NAND3_X1 port map( A1 => n55, A2 => n56, A3 => n57, ZN => 
                           carry_36_port);
   U109 : NAND2_X1 port map( A1 => A(36), A2 => B(36), ZN => n58);
   U110 : NAND2_X1 port map( A1 => A(36), A2 => carry_36_port, ZN => n59);
   U111 : NAND2_X1 port map( A1 => B(36), A2 => carry_36_port, ZN => n60);
   U112 : NAND3_X1 port map( A1 => n60, A2 => n59, A3 => n58, ZN => 
                           carry_37_port);
   U113 : XOR2_X1 port map( A => A(25), B => B(25), Z => n61);
   U114 : XOR2_X1 port map( A => n51, B => n61, Z => SUM(25));
   U115 : NAND2_X1 port map( A1 => carry_25_port, A2 => n4, ZN => n62);
   U116 : NAND2_X1 port map( A1 => carry_25_port, A2 => B(25), ZN => n63);
   U117 : NAND2_X1 port map( A1 => n4, A2 => B(25), ZN => n64);
   U118 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => 
                           carry_26_port);
   U119 : XNOR2_X1 port map( A => n65, B => n77, ZN => SUM(33));
   U120 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n65);
   U121 : XOR2_X1 port map( A => A(38), B => B(38), Z => n66);
   U122 : XOR2_X1 port map( A => n66, B => carry_38_port, Z => SUM(38));
   U123 : NAND2_X1 port map( A1 => A(38), A2 => B(38), ZN => n67);
   U124 : NAND2_X1 port map( A1 => A(38), A2 => carry_38_port, ZN => n68);
   U125 : NAND2_X1 port map( A1 => B(38), A2 => carry_38_port, ZN => n69);
   U126 : NAND3_X1 port map( A1 => n69, A2 => n68, A3 => n67, ZN => 
                           carry_39_port);
   U127 : XOR2_X1 port map( A => A(39), B => B(39), Z => n70);
   U128 : XOR2_X1 port map( A => n70, B => n24, Z => SUM(39));
   U129 : NAND2_X1 port map( A1 => A(39), A2 => B(39), ZN => n71);
   U130 : NAND2_X1 port map( A1 => A(39), A2 => carry_39_port, ZN => n72);
   U131 : NAND2_X1 port map( A1 => B(39), A2 => n23, ZN => n73);
   U132 : NAND3_X1 port map( A1 => n73, A2 => n72, A3 => n71, ZN => 
                           carry_40_port);
   U133 : NAND3_X1 port map( A1 => n86, A2 => n85, A3 => n84, ZN => n74);
   U134 : CLKBUF_X1 port map( A => carry_51_port, Z => n75);
   U135 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n76);
   U136 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n77);
   U137 : NAND3_X1 port map( A1 => n157, A2 => n156, A3 => n158, ZN => n78);
   U138 : NAND3_X1 port map( A1 => n156, A2 => n157, A3 => n158, ZN => n79);
   U139 : XOR2_X1 port map( A => A(32), B => B(32), Z => n80);
   U140 : XOR2_X1 port map( A => n80, B => carry_32_port, Z => SUM(32));
   U141 : NAND2_X1 port map( A1 => A(32), A2 => B(32), ZN => n81);
   U142 : NAND2_X1 port map( A1 => A(32), A2 => carry_32_port, ZN => n82);
   U143 : NAND2_X1 port map( A1 => B(32), A2 => carry_32_port, ZN => n83);
   U144 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => 
                           carry_33_port);
   U145 : NAND2_X1 port map( A1 => A(33), A2 => B(33), ZN => n84);
   U146 : NAND2_X1 port map( A1 => A(33), A2 => carry_33_port, ZN => n85);
   U147 : NAND2_X1 port map( A1 => B(33), A2 => n76, ZN => n86);
   U148 : NAND3_X1 port map( A1 => n86, A2 => n85, A3 => n84, ZN => 
                           carry_34_port);
   U149 : NAND2_X1 port map( A1 => n48, A2 => A(11), ZN => n87);
   U150 : NAND2_X1 port map( A1 => n48, A2 => B(11), ZN => n88);
   U151 : NAND2_X1 port map( A1 => A(11), A2 => B(11), ZN => n89);
   U152 : NAND3_X1 port map( A1 => n88, A2 => n87, A3 => n89, ZN => 
                           carry_12_port);
   U153 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => n90);
   U154 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => n91);
   U155 : XNOR2_X1 port map( A => n92, B => carry_48_port, ZN => SUM(48));
   U156 : XOR2_X1 port map( A => A(48), B => n103, Z => n92);
   U157 : XOR2_X1 port map( A => A(15), B => B(15), Z => n93);
   U158 : XOR2_X1 port map( A => carry_15_port, B => n93, Z => SUM(15));
   U159 : NAND2_X1 port map( A1 => n50, A2 => B(15), ZN => n94);
   U160 : NAND2_X1 port map( A1 => carry_15_port, A2 => n50, ZN => n95);
   U161 : NAND2_X1 port map( A1 => carry_15_port, A2 => B(15), ZN => n96);
   U162 : NAND3_X1 port map( A1 => n96, A2 => n95, A3 => n94, ZN => 
                           carry_16_port);
   U163 : XOR2_X1 port map( A => A(16), B => B(16), Z => n97);
   U164 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => n98);
   U165 : NAND2_X1 port map( A1 => carry_16_port, A2 => A(16), ZN => n99);
   U166 : NAND2_X1 port map( A1 => B(16), A2 => n53, ZN => n100);
   U167 : NAND3_X1 port map( A1 => n100, A2 => n99, A3 => n98, ZN => 
                           carry_17_port);
   U168 : XNOR2_X1 port map( A => A(60), B => B(60), ZN => n104);
   U169 : XNOR2_X1 port map( A => net17921, B => net98278, ZN => SUM(7));
   U170 : XNOR2_X1 port map( A => n101, B => carry_59_port, ZN => SUM(59));
   U171 : XNOR2_X1 port map( A => A(59), B => B(59), ZN => n101);
   U172 : CLKBUF_X1 port map( A => n74, Z => n102);
   U173 : XNOR2_X1 port map( A => n104, B => carry_60_port, ZN => SUM(60));
   U174 : XNOR2_X1 port map( A => carry_43_port, B => n105, ZN => SUM(43));
   U175 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n105);
   U176 : XOR2_X1 port map( A => A(50), B => B(50), Z => n106);
   U177 : XOR2_X1 port map( A => carry_50_port, B => n106, Z => SUM(50));
   U178 : NAND2_X1 port map( A1 => carry_50_port, A2 => A(50), ZN => n107);
   U179 : NAND2_X1 port map( A1 => carry_50_port, A2 => B(50), ZN => n108);
   U180 : NAND2_X1 port map( A1 => A(50), A2 => B(50), ZN => n109);
   U181 : NAND3_X1 port map( A1 => n107, A2 => n108, A3 => n109, ZN => 
                           carry_51_port);
   U182 : XOR2_X1 port map( A => A(51), B => B(51), Z => n110);
   U183 : XOR2_X1 port map( A => n75, B => n110, Z => SUM(51));
   U184 : NAND2_X1 port map( A1 => carry_51_port, A2 => A(51), ZN => n111);
   U185 : NAND2_X1 port map( A1 => carry_51_port, A2 => B(51), ZN => n112);
   U186 : NAND2_X1 port map( A1 => A(51), A2 => B(51), ZN => n113);
   U187 : NAND3_X1 port map( A1 => n111, A2 => n112, A3 => n113, ZN => 
                           carry_52_port);
   U188 : XOR2_X1 port map( A => A(40), B => B(40), Z => n114);
   U189 : XOR2_X1 port map( A => n114, B => carry_40_port, Z => SUM(40));
   U190 : NAND2_X1 port map( A1 => A(40), A2 => B(40), ZN => n115);
   U191 : NAND2_X1 port map( A1 => A(40), A2 => n25, ZN => n116);
   U192 : NAND2_X1 port map( A1 => B(40), A2 => carry_40_port, ZN => n117);
   U193 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => 
                           carry_41_port);
   U194 : XOR2_X1 port map( A => A(41), B => B(41), Z => n118);
   U195 : XOR2_X1 port map( A => n118, B => n91, Z => SUM(41));
   U196 : NAND2_X1 port map( A1 => A(41), A2 => B(41), ZN => n119);
   U197 : NAND2_X1 port map( A1 => n90, A2 => A(41), ZN => n120);
   U198 : NAND2_X1 port map( A1 => B(41), A2 => carry_41_port, ZN => n121);
   U199 : NAND3_X1 port map( A1 => n121, A2 => n120, A3 => n119, ZN => 
                           carry_42_port);
   U200 : XOR2_X1 port map( A => A(30), B => B(30), Z => n122);
   U201 : XOR2_X1 port map( A => carry_30_port, B => n122, Z => SUM(30));
   U202 : NAND2_X1 port map( A1 => carry_30_port, A2 => n5, ZN => n123);
   U203 : NAND2_X1 port map( A1 => carry_30_port, A2 => B(30), ZN => n124);
   U204 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n125);
   U205 : NAND3_X1 port map( A1 => n123, A2 => n124, A3 => n125, ZN => 
                           carry_31_port);
   U206 : XOR2_X1 port map( A => A(27), B => B(27), Z => n126);
   U207 : XOR2_X1 port map( A => n1, B => n126, Z => SUM(27));
   U208 : NAND2_X1 port map( A1 => n1, A2 => A(27), ZN => n127);
   U209 : NAND2_X1 port map( A1 => carry_27_port, A2 => B(27), ZN => n128);
   U210 : NAND2_X1 port map( A1 => A(27), A2 => B(27), ZN => n129);
   U211 : NAND3_X1 port map( A1 => n127, A2 => n128, A3 => n129, ZN => 
                           carry_28_port);
   U212 : XOR2_X1 port map( A => A(46), B => B(46), Z => n130);
   U213 : XOR2_X1 port map( A => carry_46_port, B => n130, Z => SUM(46));
   U214 : NAND2_X1 port map( A1 => carry_46_port, A2 => A(46), ZN => n131);
   U215 : NAND2_X1 port map( A1 => carry_46_port, A2 => B(46), ZN => n132);
   U216 : NAND2_X1 port map( A1 => A(46), A2 => B(46), ZN => n133);
   U217 : NAND3_X1 port map( A1 => n131, A2 => n132, A3 => n133, ZN => 
                           carry_47_port);
   U218 : XOR2_X1 port map( A => A(28), B => B(28), Z => n134);
   U219 : NAND2_X1 port map( A1 => n21, A2 => A(28), ZN => n135);
   U220 : NAND2_X1 port map( A1 => carry_28_port, A2 => B(28), ZN => n136);
   U221 : NAND2_X1 port map( A1 => A(28), A2 => B(28), ZN => n137);
   U222 : NAND3_X1 port map( A1 => n135, A2 => n136, A3 => n137, ZN => 
                           carry_29_port);
   U223 : NAND2_X1 port map( A1 => A(59), A2 => B(59), ZN => n138);
   U224 : NAND2_X1 port map( A1 => A(59), A2 => carry_59_port, ZN => n139);
   U225 : NAND2_X1 port map( A1 => B(59), A2 => carry_59_port, ZN => n140);
   U226 : NAND3_X1 port map( A1 => n138, A2 => n139, A3 => n140, ZN => 
                           carry_60_port);
   U227 : NAND2_X1 port map( A1 => A(60), A2 => B(60), ZN => n141);
   U228 : NAND2_X1 port map( A1 => A(60), A2 => carry_60_port, ZN => n142);
   U229 : NAND2_X1 port map( A1 => B(60), A2 => carry_60_port, ZN => n143);
   U230 : NAND3_X1 port map( A1 => n141, A2 => n142, A3 => n143, ZN => 
                           carry_61_port);
   U231 : XOR2_X1 port map( A => A(47), B => B(47), Z => n144);
   U232 : XOR2_X1 port map( A => n144, B => carry_47_port, Z => SUM(47));
   U233 : NAND2_X1 port map( A1 => A(47), A2 => B(47), ZN => n145);
   U234 : NAND2_X1 port map( A1 => A(47), A2 => carry_47_port, ZN => n146);
   U235 : NAND2_X1 port map( A1 => B(47), A2 => carry_47_port, ZN => n147);
   U236 : NAND3_X1 port map( A1 => n145, A2 => n146, A3 => n147, ZN => 
                           carry_48_port);
   U237 : NAND2_X1 port map( A1 => A(48), A2 => B(48), ZN => n148);
   U238 : NAND2_X1 port map( A1 => A(48), A2 => carry_48_port, ZN => n149);
   U239 : NAND2_X1 port map( A1 => B(48), A2 => carry_48_port, ZN => n150);
   U240 : NAND3_X1 port map( A1 => n150, A2 => n149, A3 => n148, ZN => 
                           carry_49_port);
   U241 : XOR2_X1 port map( A => A(34), B => B(34), Z => n151);
   U242 : XOR2_X1 port map( A => n102, B => n151, Z => SUM(34));
   U243 : NAND2_X1 port map( A1 => n74, A2 => n6, ZN => n152);
   U244 : NAND2_X1 port map( A1 => carry_34_port, A2 => B(34), ZN => n153);
   U245 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => n154);
   U246 : NAND3_X1 port map( A1 => n152, A2 => n153, A3 => n154, ZN => 
                           carry_35_port);
   U247 : XOR2_X1 port map( A => A(22), B => B(22), Z => n155);
   U248 : XOR2_X1 port map( A => n155, B => carry_22_port, Z => SUM(22));
   U249 : NAND2_X1 port map( A1 => n3, A2 => B(22), ZN => n156);
   U250 : NAND2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => n157);
   U251 : NAND2_X1 port map( A1 => B(22), A2 => carry_22_port, ZN => n158);
   U252 : NAND3_X1 port map( A1 => n158, A2 => n157, A3 => n156, ZN => 
                           carry_23_port);
   U253 : XOR2_X1 port map( A => n159, B => n79, Z => SUM(23));
   U254 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n160);
   U255 : NAND2_X1 port map( A1 => A(23), A2 => n78, ZN => n161);
   U256 : NAND2_X1 port map( A1 => carry_23_port, A2 => B(23), ZN => n162);
   U257 : NAND3_X1 port map( A1 => n160, A2 => n161, A3 => n162, ZN => 
                           carry_24_port);
   U258 : NAND2_X1 port map( A1 => carry_19_port, A2 => A(19), ZN => n163);
   U259 : NAND2_X1 port map( A1 => carry_19_port, A2 => B(19), ZN => n164);
   U260 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n165);
   U261 : NAND3_X1 port map( A1 => n164, A2 => n163, A3 => n165, ZN => 
                           carry_20_port);
   U262 : NAND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => n166);
   U263 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n167);
   U264 : NAND2_X1 port map( A1 => A(13), A2 => B(13), ZN => n168);
   U265 : NAND3_X1 port map( A1 => n167, A2 => n166, A3 => n168, ZN => 
                           carry_14_port);
   U266 : CLKBUF_X1 port map( A => n49, Z => n169);
   U267 : XOR2_X1 port map( A => net18132, B => net17991, Z => SUM(5));
   U268 : NAND2_X1 port map( A1 => n49, A2 => A(17), ZN => n170);
   U269 : NAND2_X1 port map( A1 => carry_17_port, A2 => B(17), ZN => n171);
   U270 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n172);
   U271 : NAND3_X1 port map( A1 => n170, A2 => n171, A3 => n172, ZN => 
                           carry_18_port);
   U272 : NAND2_X1 port map( A1 => carry_43_port, A2 => A(43), ZN => n173);
   U273 : NAND2_X1 port map( A1 => carry_43_port, A2 => B(43), ZN => n174);
   U274 : NAND2_X1 port map( A1 => A(43), A2 => B(43), ZN => n175);
   U275 : NAND3_X1 port map( A1 => n173, A2 => n174, A3 => n175, ZN => 
                           carry_44_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_0_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_0_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_0_DW01_add_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_33_port, carry_32_port, 
      carry_31_port, carry_30_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_13_port, carry_10_port, net17757, net17756, 
      net17755, net17893, net17909, net17908, net17907, net17916, net18110, 
      carry_2_port, carry_1_port, net17953, net25658, net25657, net25656, 
      net25665, net25729, net25739, net25741, net25651, carry_3_port, net17990,
      carry_9_port, net99960, net99950, net25731, net25663, net17872, net17871,
      net17870, carry_4_port, net25652, net25650, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235 : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => n86, ZN => n1);
   U2 : CLKBUF_X1 port map( A => A(4), Z => net25663);
   U3 : NAND3_X1 port map( A1 => n217, A2 => n218, A3 => n219, ZN => n2);
   U4 : NAND3_X1 port map( A1 => n175, A2 => n174, A3 => n176, ZN => n3);
   U5 : XOR2_X1 port map( A => B(44), B => A(44), Z => n4);
   U6 : XOR2_X1 port map( A => carry_44_port, B => n4, Z => SUM(44));
   U7 : NAND2_X1 port map( A1 => carry_44_port, A2 => B(44), ZN => n5);
   U8 : NAND2_X1 port map( A1 => carry_44_port, A2 => A(44), ZN => n6);
   U9 : NAND2_X1 port map( A1 => B(44), A2 => A(44), ZN => n7);
   U10 : NAND3_X1 port map( A1 => n5, A2 => n6, A3 => n7, ZN => carry_45_port);
   U11 : XNOR2_X1 port map( A => carry_21_port, B => n8, ZN => SUM(21));
   U12 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n8);
   U13 : OR2_X1 port map( A1 => A(5), A2 => B(5), ZN => n9);
   U14 : NAND2_X1 port map( A1 => n43, A2 => n9, ZN => n44);
   U15 : XOR2_X1 port map( A => B(51), B => A(51), Z => n10);
   U16 : XOR2_X1 port map( A => carry_51_port, B => n10, Z => SUM(51));
   U17 : NAND2_X1 port map( A1 => carry_51_port, A2 => B(51), ZN => n11);
   U18 : NAND2_X1 port map( A1 => carry_51_port, A2 => A(51), ZN => n12);
   U19 : NAND2_X1 port map( A1 => B(51), A2 => A(51), ZN => n13);
   U20 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => 
                           carry_52_port);
   U21 : XOR2_X1 port map( A => B(58), B => A(58), Z => n14);
   U22 : XOR2_X1 port map( A => carry_58_port, B => n14, Z => SUM(58));
   U23 : NAND2_X1 port map( A1 => carry_58_port, A2 => B(58), ZN => n15);
   U24 : NAND2_X1 port map( A1 => carry_58_port, A2 => A(58), ZN => n16);
   U25 : NAND2_X1 port map( A1 => B(58), A2 => A(58), ZN => n17);
   U26 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => n17, ZN => 
                           carry_59_port);
   U27 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => n18);
   U28 : XOR2_X1 port map( A => B(53), B => A(53), Z => n19);
   U29 : XOR2_X1 port map( A => carry_53_port, B => n19, Z => SUM(53));
   U30 : NAND2_X1 port map( A1 => carry_53_port, A2 => B(53), ZN => n20);
   U31 : NAND2_X1 port map( A1 => carry_53_port, A2 => A(53), ZN => n21);
   U32 : NAND2_X1 port map( A1 => B(53), A2 => A(53), ZN => n22);
   U33 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => 
                           carry_54_port);
   U34 : NAND3_X1 port map( A1 => n217, A2 => n218, A3 => n219, ZN => n23);
   U35 : NAND3_X1 port map( A1 => n204, A2 => n203, A3 => n202, ZN => n24);
   U36 : NAND3_X1 port map( A1 => n153, A2 => n152, A3 => n151, ZN => n25);
   U37 : NAND3_X1 port map( A1 => n175, A2 => n174, A3 => n176, ZN => n26);
   U38 : NAND3_X1 port map( A1 => n175, A2 => n174, A3 => n176, ZN => n27);
   U39 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => n28);
   U40 : NAND3_X1 port map( A1 => n114, A2 => n113, A3 => n112, ZN => n29);
   U41 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => n30);
   U42 : NAND3_X1 port map( A1 => n75, A2 => n76, A3 => n77, ZN => n31);
   U43 : NAND3_X1 port map( A1 => n76, A2 => n75, A3 => n77, ZN => n32);
   U44 : NAND3_X1 port map( A1 => n102, A2 => n101, A3 => n100, ZN => n33);
   U45 : NAND3_X1 port map( A1 => n138, A2 => n137, A3 => n136, ZN => n34);
   U46 : NAND3_X1 port map( A1 => n166, A2 => n165, A3 => n164, ZN => n35);
   U47 : NAND3_X1 port map( A1 => n166, A2 => n165, A3 => n164, ZN => n36);
   U48 : CLKBUF_X1 port map( A => B(2), Z => n37);
   U49 : NAND2_X1 port map( A1 => n59, A2 => A(9), ZN => n38);
   U50 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n39);
   U51 : NAND3_X1 port map( A1 => n138, A2 => n137, A3 => n136, ZN => 
                           carry_30_port);
   U52 : NAND3_X1 port map( A1 => n114, A2 => n113, A3 => n112, ZN => 
                           carry_40_port);
   U53 : NAND3_X1 port map( A1 => n102, A2 => n101, A3 => n100, ZN => 
                           carry_50_port);
   U54 : NAND2_X1 port map( A1 => n40, A2 => B(3), ZN => net25650);
   U55 : NAND3_X1 port map( A1 => net25650, A2 => net25652, A3 => net25651, ZN 
                           => net25731);
   U56 : NAND3_X1 port map( A1 => net25650, A2 => net25651, A3 => net25652, ZN 
                           => net25741);
   U57 : NAND3_X1 port map( A1 => net25650, A2 => net25652, A3 => net25651, ZN 
                           => carry_4_port);
   U58 : NAND3_X1 port map( A1 => net25658, A2 => net25657, A3 => net25656, ZN 
                           => n40);
   U59 : CLKBUF_X1 port map( A => n40, Z => net25665);
   U60 : CLKBUF_X1 port map( A => B(3), Z => net25739);
   U61 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => net25652);
   U62 : NAND3_X1 port map( A1 => net25658, A2 => net25657, A3 => net25656, ZN 
                           => carry_3_port);
   U63 : NAND2_X1 port map( A1 => n44, A2 => n42, ZN => net99950);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n42, ZN => net99960);
   U65 : NAND3_X1 port map( A1 => net17871, A2 => net17870, A3 => net17872, ZN 
                           => n43);
   U66 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n42);
   U67 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => net17916);
   U68 : NAND2_X1 port map( A1 => carry_4_port, A2 => net25663, ZN => net17871)
                           ;
   U69 : NAND3_X1 port map( A1 => net17870, A2 => net17872, A3 => net17871, ZN 
                           => net17893);
   U70 : NAND2_X1 port map( A1 => n41, A2 => net25663, ZN => net17872);
   U71 : NAND2_X1 port map( A1 => net25731, A2 => n41, ZN => net17870);
   U72 : BUF_X1 port map( A => B(4), Z => n41);
   U73 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => net17953);
   U74 : XNOR2_X1 port map( A => net99950, B => n45, ZN => SUM(6));
   U75 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n45);
   U76 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => net17755);
   U77 : NAND2_X1 port map( A1 => net99960, A2 => B(6), ZN => net17757);
   U78 : NAND2_X1 port map( A1 => net99960, A2 => A(6), ZN => net17756);
   U79 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => n54);
   U80 : XNOR2_X1 port map( A => n47, B => n46, ZN => SUM(7));
   U81 : XOR2_X1 port map( A => A(7), B => n52, Z => n46);
   U82 : NAND3_X1 port map( A1 => net17757, A2 => net17756, A3 => net17755, ZN 
                           => n47);
   U83 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n48);
   U84 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => net17990);
   U85 : NAND3_X1 port map( A1 => net17756, A2 => net17757, A3 => net17755, ZN 
                           => n53);
   U86 : NAND2_X1 port map( A1 => A(7), A2 => B(7), ZN => n50);
   U87 : INV_X1 port map( A => A(7), ZN => n51);
   U88 : INV_X1 port map( A => B(7), ZN => n52);
   U89 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n49);
   U90 : XNOR2_X1 port map( A => n60, B => n58, ZN => SUM(9));
   U91 : XNOR2_X1 port map( A => A(9), B => B(9), ZN => n58);
   U92 : NAND3_X1 port map( A1 => n56, A2 => n61, A3 => n57, ZN => n60);
   U93 : NAND2_X1 port map( A1 => n59, A2 => A(9), ZN => net17907);
   U94 : NAND2_X1 port map( A1 => A(9), A2 => B(9), ZN => net17909);
   U95 : NAND2_X1 port map( A1 => carry_9_port, A2 => B(9), ZN => net17908);
   U96 : NAND2_X1 port map( A1 => net17990, A2 => A(8), ZN => n61);
   U97 : NAND3_X1 port map( A1 => n56, A2 => n61, A3 => n57, ZN => n59);
   U98 : NAND2_X1 port map( A1 => net17990, A2 => B(8), ZN => n56);
   U99 : NAND3_X1 port map( A1 => n56, A2 => n55, A3 => n57, ZN => carry_9_port
                           );
   U100 : NAND2_X1 port map( A1 => A(8), A2 => B(8), ZN => n57);
   U101 : NAND2_X1 port map( A1 => n48, A2 => A(8), ZN => n55);
   U102 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => net18110);
   U103 : XOR2_X1 port map( A => A(14), B => B(14), Z => n62);
   U104 : XOR2_X1 port map( A => n3, B => n62, Z => SUM(14));
   U105 : NAND2_X1 port map( A1 => n27, A2 => A(14), ZN => n63);
   U106 : NAND2_X1 port map( A1 => n26, A2 => B(14), ZN => n64);
   U107 : NAND2_X1 port map( A1 => A(14), A2 => B(14), ZN => n65);
   U108 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => 
                           carry_15_port);
   U109 : XNOR2_X1 port map( A => carry_10_port, B => n66, ZN => SUM(10));
   U110 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n66);
   U111 : XNOR2_X1 port map( A => n67, B => n170, ZN => SUM(12));
   U112 : AND3_X1 port map( A1 => n185, A2 => n186, A3 => n187, ZN => n67);
   U113 : XNOR2_X1 port map( A => n68, B => n36, ZN => SUM(23));
   U114 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n68);
   U115 : XNOR2_X1 port map( A => n184, B => n69, ZN => SUM(11));
   U116 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => n69);
   U117 : XOR2_X1 port map( A => B(35), B => A(35), Z => n70);
   U118 : XOR2_X1 port map( A => n24, B => n70, Z => SUM(35));
   U119 : NAND2_X1 port map( A1 => n24, A2 => B(35), ZN => n71);
   U120 : NAND2_X1 port map( A1 => carry_35_port, A2 => A(35), ZN => n72);
   U121 : NAND2_X1 port map( A1 => B(35), A2 => A(35), ZN => n73);
   U122 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => 
                           carry_36_port);
   U123 : XOR2_X1 port map( A => A(28), B => B(28), Z => n74);
   U124 : XOR2_X1 port map( A => carry_28_port, B => n74, Z => SUM(28));
   U125 : NAND2_X1 port map( A1 => carry_28_port, A2 => A(28), ZN => n75);
   U126 : NAND2_X1 port map( A1 => carry_28_port, A2 => B(28), ZN => n76);
   U127 : NAND2_X1 port map( A1 => A(28), A2 => B(28), ZN => n77);
   U128 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n94, ZN => n78);
   U129 : NAND3_X1 port map( A1 => n167, A2 => n168, A3 => n169, ZN => n79);
   U130 : XNOR2_X1 port map( A => n87, B => n80, ZN => SUM(13));
   U131 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n80);
   U132 : NAND3_X1 port map( A1 => n85, A2 => n84, A3 => n86, ZN => n81);
   U133 : NAND2_X1 port map( A1 => carry_3_port, A2 => A(3), ZN => net25651);
   U134 : CLKBUF_X1 port map( A => A(3), Z => net25729);
   U135 : NAND3_X1 port map( A1 => n108, A2 => n109, A3 => n110, ZN => n82);
   U136 : XNOR2_X1 port map( A => n83, B => n89, ZN => SUM(19));
   U137 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n83);
   U138 : NAND2_X1 port map( A1 => n78, A2 => A(21), ZN => n84);
   U139 : NAND2_X1 port map( A1 => n78, A2 => B(21), ZN => n85);
   U140 : NAND2_X1 port map( A1 => A(21), A2 => B(21), ZN => n86);
   U141 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => n86, ZN => 
                           carry_22_port);
   U142 : NAND3_X1 port map( A1 => n171, A2 => n172, A3 => n173, ZN => n87);
   U143 : NAND3_X1 port map( A1 => n233, A2 => n234, A3 => n235, ZN => n88);
   U144 : NAND3_X1 port map( A1 => n150, A2 => n149, A3 => n148, ZN => n89);
   U145 : NAND3_X1 port map( A1 => n178, A2 => n179, A3 => n180, ZN => n90);
   U146 : XOR2_X1 port map( A => A(20), B => B(20), Z => n91);
   U147 : XOR2_X1 port map( A => n25, B => n91, Z => SUM(20));
   U148 : NAND2_X1 port map( A1 => n25, A2 => A(20), ZN => n92);
   U149 : NAND2_X1 port map( A1 => carry_20_port, A2 => B(20), ZN => n93);
   U150 : NAND2_X1 port map( A1 => A(20), A2 => B(20), ZN => n94);
   U151 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n94, ZN => 
                           carry_21_port);
   U152 : XOR2_X1 port map( A => B(48), B => A(48), Z => n95);
   U153 : XOR2_X1 port map( A => carry_48_port, B => n95, Z => SUM(48));
   U154 : NAND2_X1 port map( A1 => carry_48_port, A2 => B(48), ZN => n96);
   U155 : NAND2_X1 port map( A1 => carry_48_port, A2 => A(48), ZN => n97);
   U156 : NAND2_X1 port map( A1 => B(48), A2 => A(48), ZN => n98);
   U157 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => 
                           carry_49_port);
   U158 : XOR2_X1 port map( A => A(49), B => B(49), Z => n99);
   U159 : XOR2_X1 port map( A => n99, B => n30, Z => SUM(49));
   U160 : NAND2_X1 port map( A1 => A(49), A2 => B(49), ZN => n100);
   U161 : NAND2_X1 port map( A1 => A(49), A2 => carry_49_port, ZN => n101);
   U162 : NAND2_X1 port map( A1 => B(49), A2 => n30, ZN => n102);
   U163 : XOR2_X1 port map( A => A(50), B => B(50), Z => n103);
   U164 : XOR2_X1 port map( A => n103, B => n33, Z => SUM(50));
   U165 : NAND2_X1 port map( A1 => A(50), A2 => B(50), ZN => n104);
   U166 : NAND2_X1 port map( A1 => A(50), A2 => n33, ZN => n105);
   U167 : NAND2_X1 port map( A1 => B(50), A2 => carry_50_port, ZN => n106);
   U168 : NAND3_X1 port map( A1 => n104, A2 => n105, A3 => n106, ZN => 
                           carry_51_port);
   U169 : XOR2_X1 port map( A => B(38), B => A(38), Z => n107);
   U170 : XOR2_X1 port map( A => n23, B => n107, Z => SUM(38));
   U171 : NAND2_X1 port map( A1 => carry_38_port, A2 => B(38), ZN => n108);
   U172 : NAND2_X1 port map( A1 => n2, A2 => A(38), ZN => n109);
   U173 : NAND2_X1 port map( A1 => B(38), A2 => A(38), ZN => n110);
   U174 : NAND3_X1 port map( A1 => n108, A2 => n109, A3 => n110, ZN => 
                           carry_39_port);
   U175 : XOR2_X1 port map( A => A(39), B => B(39), Z => n111);
   U176 : XOR2_X1 port map( A => n111, B => n82, Z => SUM(39));
   U177 : NAND2_X1 port map( A1 => A(39), A2 => B(39), ZN => n112);
   U178 : NAND2_X1 port map( A1 => carry_39_port, A2 => A(39), ZN => n113);
   U179 : NAND2_X1 port map( A1 => B(39), A2 => carry_39_port, ZN => n114);
   U180 : XOR2_X1 port map( A => A(40), B => B(40), Z => n115);
   U181 : XOR2_X1 port map( A => n115, B => n29, Z => SUM(40));
   U182 : NAND2_X1 port map( A1 => A(40), A2 => B(40), ZN => n116);
   U183 : NAND2_X1 port map( A1 => A(40), A2 => carry_40_port, ZN => n117);
   U184 : NAND2_X1 port map( A1 => carry_40_port, A2 => B(40), ZN => n118);
   U185 : NAND3_X1 port map( A1 => n116, A2 => n117, A3 => n118, ZN => 
                           carry_41_port);
   U186 : XOR2_X1 port map( A => B(61), B => A(61), Z => n119);
   U187 : XOR2_X1 port map( A => carry_61_port, B => n119, Z => SUM(61));
   U188 : NAND2_X1 port map( A1 => carry_61_port, A2 => B(61), ZN => n120);
   U189 : NAND2_X1 port map( A1 => carry_61_port, A2 => A(61), ZN => n121);
   U190 : NAND2_X1 port map( A1 => B(61), A2 => A(61), ZN => n122);
   U191 : NAND3_X1 port map( A1 => n120, A2 => n121, A3 => n122, ZN => 
                           carry_62_port);
   U192 : XOR2_X1 port map( A => A(32), B => B(32), Z => n123);
   U193 : XOR2_X1 port map( A => carry_32_port, B => n123, Z => SUM(32));
   U194 : NAND2_X1 port map( A1 => carry_32_port, A2 => A(32), ZN => n124);
   U195 : NAND2_X1 port map( A1 => carry_32_port, A2 => B(32), ZN => n125);
   U196 : NAND2_X1 port map( A1 => A(32), A2 => B(32), ZN => n126);
   U197 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => 
                           carry_33_port);
   U198 : XOR2_X1 port map( A => A(24), B => B(24), Z => n127);
   U199 : XOR2_X1 port map( A => carry_24_port, B => n127, Z => SUM(24));
   U200 : NAND2_X1 port map( A1 => n79, A2 => A(24), ZN => n128);
   U201 : NAND2_X1 port map( A1 => carry_24_port, A2 => B(24), ZN => n129);
   U202 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n130);
   U203 : NAND3_X1 port map( A1 => n128, A2 => n129, A3 => n130, ZN => 
                           carry_25_port);
   U204 : XOR2_X1 port map( A => B(54), B => A(54), Z => n131);
   U205 : XOR2_X1 port map( A => carry_54_port, B => n131, Z => SUM(54));
   U206 : NAND2_X1 port map( A1 => carry_54_port, A2 => B(54), ZN => n132);
   U207 : NAND2_X1 port map( A1 => carry_54_port, A2 => A(54), ZN => n133);
   U208 : NAND2_X1 port map( A1 => B(54), A2 => A(54), ZN => n134);
   U209 : NAND3_X1 port map( A1 => n132, A2 => n133, A3 => n134, ZN => 
                           carry_55_port);
   U210 : XOR2_X1 port map( A => A(29), B => B(29), Z => n135);
   U211 : XOR2_X1 port map( A => n135, B => n32, Z => SUM(29));
   U212 : NAND2_X1 port map( A1 => A(29), A2 => B(29), ZN => n136);
   U213 : NAND2_X1 port map( A1 => A(29), A2 => n31, ZN => n137);
   U214 : NAND2_X1 port map( A1 => B(29), A2 => n31, ZN => n138);
   U215 : XOR2_X1 port map( A => A(30), B => B(30), Z => n139);
   U216 : XOR2_X1 port map( A => n139, B => carry_30_port, Z => SUM(30));
   U217 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n140);
   U218 : NAND2_X1 port map( A1 => A(30), A2 => carry_30_port, ZN => n141);
   U219 : NAND2_X1 port map( A1 => B(30), A2 => n34, ZN => n142);
   U220 : NAND3_X1 port map( A1 => n142, A2 => n141, A3 => n140, ZN => 
                           carry_31_port);
   U221 : NAND3_X1 port map( A1 => n206, A2 => n207, A3 => n208, ZN => n143);
   U222 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n144);
   U223 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n145);
   U224 : NAND3_X1 port map( A1 => n191, A2 => n190, A3 => n192, ZN => n146);
   U225 : XOR2_X1 port map( A => A(18), B => B(18), Z => n147);
   U226 : XOR2_X1 port map( A => n147, B => n88, Z => SUM(18));
   U227 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n148);
   U228 : NAND2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => n149);
   U229 : NAND2_X1 port map( A1 => B(18), A2 => carry_18_port, ZN => n150);
   U230 : NAND3_X1 port map( A1 => n148, A2 => n149, A3 => n150, ZN => 
                           carry_19_port);
   U231 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n151);
   U232 : NAND2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => n152);
   U233 : NAND2_X1 port map( A1 => B(19), A2 => carry_19_port, ZN => n153);
   U234 : NAND3_X1 port map( A1 => n151, A2 => n152, A3 => n153, ZN => 
                           carry_20_port);
   U235 : NAND3_X1 port map( A1 => n186, A2 => n185, A3 => n187, ZN => n154);
   U236 : XOR2_X1 port map( A => B(45), B => A(45), Z => n155);
   U237 : XOR2_X1 port map( A => carry_45_port, B => n155, Z => SUM(45));
   U238 : NAND2_X1 port map( A1 => carry_45_port, A2 => B(45), ZN => n156);
   U239 : NAND2_X1 port map( A1 => carry_45_port, A2 => A(45), ZN => n157);
   U240 : NAND2_X1 port map( A1 => B(45), A2 => A(45), ZN => n158);
   U241 : NAND3_X1 port map( A1 => n156, A2 => n157, A3 => n158, ZN => 
                           carry_46_port);
   U242 : XOR2_X1 port map( A => A(31), B => B(31), Z => n159);
   U243 : XOR2_X1 port map( A => carry_31_port, B => n159, Z => SUM(31));
   U244 : NAND2_X1 port map( A1 => carry_31_port, A2 => A(31), ZN => n160);
   U245 : NAND2_X1 port map( A1 => carry_31_port, A2 => B(31), ZN => n161);
   U246 : NAND2_X1 port map( A1 => A(31), A2 => B(31), ZN => n162);
   U247 : NAND3_X1 port map( A1 => n160, A2 => n161, A3 => n162, ZN => 
                           carry_32_port);
   U248 : XOR2_X1 port map( A => A(22), B => B(22), Z => n163);
   U249 : XOR2_X1 port map( A => n163, B => n1, Z => SUM(22));
   U250 : NAND2_X1 port map( A1 => A(22), A2 => B(22), ZN => n164);
   U251 : NAND2_X1 port map( A1 => A(22), A2 => n81, ZN => n165);
   U252 : NAND2_X1 port map( A1 => B(22), A2 => carry_22_port, ZN => n166);
   U253 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n167);
   U254 : NAND2_X1 port map( A1 => A(23), A2 => n35, ZN => n168);
   U255 : NAND2_X1 port map( A1 => B(23), A2 => n35, ZN => n169);
   U256 : NAND3_X1 port map( A1 => n169, A2 => n168, A3 => n167, ZN => 
                           carry_24_port);
   U257 : XOR2_X1 port map( A => A(12), B => B(12), Z => n170);
   U258 : NAND2_X1 port map( A1 => n154, A2 => A(12), ZN => n171);
   U259 : NAND2_X1 port map( A1 => n154, A2 => B(12), ZN => n172);
   U260 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n173);
   U261 : NAND3_X1 port map( A1 => n171, A2 => n172, A3 => n173, ZN => 
                           carry_13_port);
   U262 : NAND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => n174);
   U263 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n175);
   U264 : NAND2_X1 port map( A1 => A(13), A2 => B(13), ZN => n176);
   U265 : XOR2_X1 port map( A => A(15), B => B(15), Z => n177);
   U266 : XOR2_X1 port map( A => carry_15_port, B => n177, Z => SUM(15));
   U267 : NAND2_X1 port map( A1 => n28, A2 => A(15), ZN => n178);
   U268 : NAND2_X1 port map( A1 => n28, A2 => B(15), ZN => n179);
   U269 : NAND2_X1 port map( A1 => A(15), A2 => B(15), ZN => n180);
   U270 : NAND3_X1 port map( A1 => n179, A2 => n178, A3 => n180, ZN => 
                           carry_16_port);
   U271 : CLKBUF_X1 port map( A => A(2), Z => n181);
   U272 : XOR2_X1 port map( A => n37, B => n181, Z => n182);
   U273 : XOR2_X1 port map( A => carry_2_port, B => n182, Z => SUM(2));
   U274 : NAND2_X1 port map( A1 => carry_2_port, A2 => n181, ZN => net25656);
   U275 : NAND2_X1 port map( A1 => B(2), A2 => carry_2_port, ZN => net25657);
   U276 : NAND2_X1 port map( A1 => A(2), A2 => B(2), ZN => net25658);
   U277 : XOR2_X1 port map( A => net25739, B => net25729, Z => n183);
   U278 : XOR2_X1 port map( A => net25665, B => n183, Z => SUM(3));
   U279 : XNOR2_X1 port map( A => net17953, B => net25741, ZN => SUM(4));
   U280 : NAND3_X1 port map( A1 => n190, A2 => n191, A3 => n192, ZN => n184);
   U281 : XNOR2_X1 port map( A => net18110, B => n48, ZN => SUM(8));
   U282 : NAND2_X1 port map( A1 => n146, A2 => A(11), ZN => n185);
   U283 : NAND2_X1 port map( A1 => n146, A2 => B(11), ZN => n186);
   U284 : NAND2_X1 port map( A1 => A(11), A2 => B(11), ZN => n187);
   U285 : NAND3_X1 port map( A1 => n38, A2 => net17908, A3 => net17909, ZN => 
                           n188);
   U286 : NAND3_X1 port map( A1 => net17908, A2 => net17909, A3 => net17907, ZN
                           => n189);
   U287 : XNOR2_X1 port map( A => net17893, B => net17916, ZN => SUM(5));
   U288 : NAND2_X1 port map( A1 => n188, A2 => A(10), ZN => n190);
   U289 : NAND2_X1 port map( A1 => n189, A2 => B(10), ZN => n191);
   U290 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => n192);
   U291 : NAND3_X1 port map( A1 => n38, A2 => net17908, A3 => net17909, ZN => 
                           carry_10_port);
   U292 : XOR2_X1 port map( A => B(41), B => A(41), Z => n193);
   U293 : XOR2_X1 port map( A => carry_41_port, B => n193, Z => SUM(41));
   U294 : NAND2_X1 port map( A1 => carry_41_port, A2 => B(41), ZN => n194);
   U295 : NAND2_X1 port map( A1 => carry_41_port, A2 => A(41), ZN => n195);
   U296 : NAND2_X1 port map( A1 => B(41), A2 => A(41), ZN => n196);
   U297 : NAND3_X1 port map( A1 => n194, A2 => n195, A3 => n196, ZN => 
                           carry_42_port);
   U298 : XOR2_X1 port map( A => A(33), B => B(33), Z => n197);
   U299 : XOR2_X1 port map( A => n197, B => n18, Z => SUM(33));
   U300 : NAND2_X1 port map( A1 => A(33), A2 => B(33), ZN => n198);
   U301 : NAND2_X1 port map( A1 => A(33), A2 => carry_33_port, ZN => n199);
   U302 : NAND2_X1 port map( A1 => B(33), A2 => n18, ZN => n200);
   U303 : XOR2_X1 port map( A => A(34), B => B(34), Z => n201);
   U304 : XOR2_X1 port map( A => n201, B => n145, Z => SUM(34));
   U305 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => n202);
   U306 : NAND2_X1 port map( A1 => n144, A2 => A(34), ZN => n203);
   U307 : NAND2_X1 port map( A1 => B(34), A2 => n144, ZN => n204);
   U308 : NAND3_X1 port map( A1 => n204, A2 => n203, A3 => n202, ZN => 
                           carry_35_port);
   U309 : XOR2_X1 port map( A => A(25), B => B(25), Z => n205);
   U310 : XOR2_X1 port map( A => carry_25_port, B => n205, Z => SUM(25));
   U311 : NAND2_X1 port map( A1 => carry_25_port, A2 => A(25), ZN => n206);
   U312 : NAND2_X1 port map( A1 => carry_25_port, A2 => B(25), ZN => n207);
   U313 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n208);
   U314 : NAND3_X1 port map( A1 => n206, A2 => n207, A3 => n208, ZN => 
                           carry_26_port);
   U315 : NAND3_X1 port map( A1 => n213, A2 => n214, A3 => n215, ZN => n209);
   U316 : NAND3_X1 port map( A1 => n222, A2 => n221, A3 => n223, ZN => n210);
   U317 : NAND3_X1 port map( A1 => n231, A2 => n230, A3 => n229, ZN => n211);
   U318 : XOR2_X1 port map( A => A(36), B => B(36), Z => n212);
   U319 : XOR2_X1 port map( A => n212, B => n39, Z => SUM(36));
   U320 : NAND2_X1 port map( A1 => A(36), A2 => B(36), ZN => n213);
   U321 : NAND2_X1 port map( A1 => A(36), A2 => carry_36_port, ZN => n214);
   U322 : NAND2_X1 port map( A1 => B(36), A2 => carry_36_port, ZN => n215);
   U323 : NAND3_X1 port map( A1 => n213, A2 => n214, A3 => n215, ZN => 
                           carry_37_port);
   U324 : XOR2_X1 port map( A => A(37), B => B(37), Z => n216);
   U325 : XOR2_X1 port map( A => n216, B => n209, Z => SUM(37));
   U326 : NAND2_X1 port map( A1 => A(37), A2 => B(37), ZN => n217);
   U327 : NAND2_X1 port map( A1 => carry_37_port, A2 => A(37), ZN => n218);
   U328 : NAND2_X1 port map( A1 => B(37), A2 => n209, ZN => n219);
   U329 : NAND3_X1 port map( A1 => n217, A2 => n218, A3 => n219, ZN => 
                           carry_38_port);
   U330 : XOR2_X1 port map( A => A(26), B => B(26), Z => n220);
   U331 : XOR2_X1 port map( A => n220, B => n143, Z => SUM(26));
   U332 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n221);
   U333 : NAND2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => n222);
   U334 : NAND2_X1 port map( A1 => B(26), A2 => carry_26_port, ZN => n223);
   U335 : NAND3_X1 port map( A1 => n223, A2 => n222, A3 => n221, ZN => 
                           carry_27_port);
   U336 : XOR2_X1 port map( A => A(27), B => B(27), Z => n224);
   U337 : XOR2_X1 port map( A => n224, B => n210, Z => SUM(27));
   U338 : NAND2_X1 port map( A1 => A(27), A2 => B(27), ZN => n225);
   U339 : NAND2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => n226);
   U340 : NAND2_X1 port map( A1 => B(27), A2 => carry_27_port, ZN => n227);
   U341 : NAND3_X1 port map( A1 => n225, A2 => n226, A3 => n227, ZN => 
                           carry_28_port);
   U342 : XOR2_X1 port map( A => A(16), B => B(16), Z => n228);
   U343 : XOR2_X1 port map( A => n228, B => n90, Z => SUM(16));
   U344 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => n229);
   U345 : NAND2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => n230);
   U346 : NAND2_X1 port map( A1 => B(16), A2 => carry_16_port, ZN => n231);
   U347 : NAND3_X1 port map( A1 => n231, A2 => n230, A3 => n229, ZN => 
                           carry_17_port);
   U348 : XOR2_X1 port map( A => A(17), B => B(17), Z => n232);
   U349 : XOR2_X1 port map( A => n232, B => n211, Z => SUM(17));
   U350 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n233);
   U351 : NAND2_X1 port map( A1 => carry_17_port, A2 => A(17), ZN => n234);
   U352 : NAND2_X1 port map( A1 => carry_17_port, A2 => B(17), ZN => n235);
   U353 : NAND3_X1 port map( A1 => n234, A2 => n233, A3 => n235, ZN => 
                           carry_18_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BOOTHMUL_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end BOOTHMUL_DW01_inc_0;

architecture SYN_rpl of BOOTHMUL_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_2_port, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => n7, CO => carry_9_port, S => SUM(8)
                           );
   U1_1_6 : HA_X1 port map( A => carry_6_port, B => A(6), CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => carry_4_port, B => A(4), CO => carry_5_port, S
                           => SUM(4));
   U1_1_1 : HA_X1 port map( A => A(0), B => A(1), CO => carry_2_port, S => 
                           SUM(1));
   U2 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U1 : BUF_X1 port map( A => carry_2_port, Z => n5);
   U3 : CLKBUF_X1 port map( A => A(0), Z => n2);
   U4 : AND2_X1 port map( A1 => carry_2_port, A2 => A(2), ZN => n3);
   U5 : XOR2_X1 port map( A => n3, B => A(3), Z => SUM(3));
   U6 : INV_X1 port map( A => n4, ZN => carry_4_port);
   U7 : NAND2_X1 port map( A1 => n3, A2 => A(3), ZN => n4);
   U8 : XOR2_X1 port map( A => n5, B => A(2), Z => SUM(2));
   U9 : AND2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => n6);
   U10 : AND2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => n7);
   U11 : XOR2_X1 port map( A => A(7), B => n6, Z => SUM(7));
   U12 : INV_X1 port map( A => n2, ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_1;

architecture SYN_BEHAVIORAL of RCA_NBIT64_1 is

   component RCA_NBIT64_1_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1045 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_1_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1045);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_2;

architecture SYN_BEHAVIORAL of RCA_NBIT64_2 is

   component RCA_NBIT64_2_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1046 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_2_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1046);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_3;

architecture SYN_BEHAVIORAL of RCA_NBIT64_3 is

   component RCA_NBIT64_3_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1047 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_3_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1047);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_4;

architecture SYN_BEHAVIORAL of RCA_NBIT64_4 is

   component RCA_NBIT64_4_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1048 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_4_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1048);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_5;

architecture SYN_BEHAVIORAL of RCA_NBIT64_5 is

   component RCA_NBIT64_5_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1049 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_5_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1049);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_6;

architecture SYN_BEHAVIORAL of RCA_NBIT64_6 is

   component RCA_NBIT64_6_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1050 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_6_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1050);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_7;

architecture SYN_BEHAVIORAL of RCA_NBIT64_7 is

   component RCA_NBIT64_7_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1051 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_7_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1051);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_8;

architecture SYN_BEHAVIORAL of RCA_NBIT64_8 is

   component RCA_NBIT64_8_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1052 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_8_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1052);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_9;

architecture SYN_BEHAVIORAL of RCA_NBIT64_9 is

   component RCA_NBIT64_9_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1053 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_9_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1053);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_10;

architecture SYN_BEHAVIORAL of RCA_NBIT64_10 is

   component RCA_NBIT64_10_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1054 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_10_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1054);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_11;

architecture SYN_BEHAVIORAL of RCA_NBIT64_11 is

   component RCA_NBIT64_11_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1055 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_11_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1055);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_12;

architecture SYN_BEHAVIORAL of RCA_NBIT64_12 is

   component RCA_NBIT64_12_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1056 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_12_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1056);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_13;

architecture SYN_BEHAVIORAL of RCA_NBIT64_13 is

   component RCA_NBIT64_13_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1057 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_13_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1057);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_14;

architecture SYN_BEHAVIORAL of RCA_NBIT64_14 is

   component RCA_NBIT64_14_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1058 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_14_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1058);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_0;

architecture SYN_BEHAVIORAL of RCA_NBIT64_0 is

   component RCA_NBIT64_0_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1059 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_53_2 : RCA_NBIT64_0_DW01_add_0 port map( A(64) => n2, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n2, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1059);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_0 is

   port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector (0 
         to 2);  Y : out std_logic_vector (0 to 63));

end MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_0;

architecture SYN_BEHAVIOR of MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_0 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, net15655, net15653, net15651, net15649, 
      net15647, net15645, net15853, net15849, net15847, net15845, net15843, 
      net15865, net15861, net15859, net15857, net15855, net15877, net15873, 
      net15871, net15869, net15867, net15889, net15887, net15885, net15883, 
      net15881, net15879, net18154, net25734, net25733, n18, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n112, A2 => n113, ZN => Y(19));
   U2 : NOR2_X1 port map( A1 => n160, A2 => n161, ZN => n136);
   U3 : NOR2_X1 port map( A1 => n162, A2 => n137, ZN => n33);
   U4 : INV_X2 port map( A => n136, ZN => n137);
   U5 : NAND2_X2 port map( A1 => n22, A2 => n23, ZN => Y(5));
   U6 : NAND2_X2 port map( A1 => n130, A2 => n131, ZN => Y(10));
   U7 : AND2_X1 port map( A1 => net15873, A2 => INPUT(186), ZN => n147);
   U8 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => Y(18));
   U9 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => Y(22));
   U10 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(9));
   U11 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => Y(15));
   U12 : BUF_X1 port map( A => n7, Z => net15887);
   U13 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => Y(2));
   U14 : NOR3_X1 port map( A1 => n156, A2 => n155, A3 => net15645, ZN => n7);
   U15 : AND2_X1 port map( A1 => n144, A2 => n145, ZN => n138);
   U16 : AND2_X1 port map( A1 => n146, A2 => n138, ZN => n139);
   U17 : OR2_X1 port map( A1 => n150, A2 => n153, ZN => n140);
   U18 : AND2_X1 port map( A1 => INPUT(123), A2 => n4, ZN => n141);
   U19 : AND2_X1 port map( A1 => INPUT(251), A2 => net25734, ZN => n142);
   U20 : AND2_X1 port map( A1 => INPUT(187), A2 => net15877, ZN => n143);
   U21 : NOR3_X1 port map( A1 => n141, A2 => n142, A3 => n143, ZN => n25);
   U22 : CLKBUF_X3 port map( A => n5, Z => net25734);
   U23 : NAND2_X1 port map( A1 => INPUT(121), A2 => net15853, ZN => n144);
   U24 : NAND2_X1 port map( A1 => INPUT(249), A2 => net25734, ZN => n145);
   U25 : NAND2_X1 port map( A1 => INPUT(185), A2 => net15867, ZN => n146);
   U26 : NOR2_X1 port map( A1 => n147, A2 => n140, ZN => n27);
   U27 : INV_X1 port map( A => net15849, ZN => n148);
   U28 : INV_X1 port map( A => INPUT(122), ZN => n149);
   U29 : NOR2_X1 port map( A1 => n148, A2 => n149, ZN => n150);
   U30 : INV_X1 port map( A => net25733, ZN => n151);
   U31 : INV_X1 port map( A => INPUT(250), ZN => n152);
   U32 : NOR2_X1 port map( A1 => n151, A2 => n152, ZN => n153);
   U33 : BUF_X2 port map( A => n5, Z => net15861);
   U34 : BUF_X2 port map( A => n6, Z => net15867);
   U35 : AND2_X2 port map( A1 => SEL(1), A2 => n154, ZN => n6);
   U36 : AND2_X2 port map( A1 => n155, A2 => SEL(1), ZN => n5);
   U37 : AOI22_X1 port map( A1 => INPUT(61), A2 => net15887, B1 => INPUT(317), 
                           B2 => net15653, ZN => n18);
   U38 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(61));
   U39 : BUF_X2 port map( A => SEL(0), Z => net15653);
   U40 : CLKBUF_X1 port map( A => SEL(0), Z => net15645);
   U41 : BUF_X1 port map( A => SEL(2), Z => n155);
   U42 : CLKBUF_X1 port map( A => SEL(1), Z => n156);
   U43 : INV_X1 port map( A => SEL(2), ZN => n154);
   U44 : NOR2_X1 port map( A1 => n154, A2 => SEL(1), ZN => n4);
   U45 : AND2_X1 port map( A1 => INPUT(120), A2 => net15847, ZN => n157);
   U46 : AND2_X1 port map( A1 => INPUT(248), A2 => net25733, ZN => n158);
   U47 : AND2_X1 port map( A1 => INPUT(184), A2 => net15869, ZN => n159);
   U48 : NOR3_X1 port map( A1 => n157, A2 => n158, A3 => n159, ZN => n31);
   U49 : AND2_X1 port map( A1 => INPUT(119), A2 => net15845, ZN => n160);
   U50 : AND2_X1 port map( A1 => INPUT(247), A2 => net25734, ZN => n161);
   U51 : AND2_X1 port map( A1 => INPUT(183), A2 => net15871, ZN => n162);
   U52 : BUF_X2 port map( A => n6, Z => net15871);
   U53 : BUF_X2 port map( A => n4, Z => net15849);
   U54 : BUF_X1 port map( A => net18154, Z => net15853);
   U55 : BUF_X2 port map( A => n5, Z => net25733);
   U56 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(60));
   U57 : BUF_X2 port map( A => n6, Z => net15873);
   U58 : CLKBUF_X1 port map( A => n4, Z => net18154);
   U59 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(59));
   U60 : CLKBUF_X1 port map( A => net18154, Z => net15847);
   U61 : CLKBUF_X1 port map( A => n5, Z => net15859);
   U62 : CLKBUF_X1 port map( A => net18154, Z => net15845);
   U63 : CLKBUF_X1 port map( A => n5, Z => net15857);
   U64 : CLKBUF_X1 port map( A => n6, Z => net15869);
   U65 : CLKBUF_X1 port map( A => net18154, Z => net15843);
   U66 : CLKBUF_X1 port map( A => n5, Z => net15855);
   U67 : CLKBUF_X1 port map( A => SEL(0), Z => net15651);
   U68 : CLKBUF_X1 port map( A => SEL(0), Z => net15649);
   U69 : CLKBUF_X1 port map( A => SEL(0), Z => net15647);
   U70 : AOI222_X1 port map( A1 => INPUT(113), A2 => net15849, B1 => INPUT(241)
                           , B2 => net15861, C1 => INPUT(177), C2 => net15873, 
                           ZN => n47);
   U71 : AOI222_X1 port map( A1 => INPUT(112), A2 => net15849, B1 => INPUT(240)
                           , B2 => net25734, C1 => INPUT(176), C2 => net15873, 
                           ZN => n49);
   U72 : AOI222_X1 port map( A1 => INPUT(111), A2 => net15849, B1 => INPUT(239)
                           , B2 => net25733, C1 => INPUT(175), C2 => net15873, 
                           ZN => n51);
   U73 : AOI222_X1 port map( A1 => INPUT(110), A2 => net15849, B1 => INPUT(238)
                           , B2 => net25734, C1 => INPUT(174), C2 => net15873, 
                           ZN => n53);
   U74 : AOI222_X1 port map( A1 => INPUT(124), A2 => net18154, B1 => INPUT(252)
                           , B2 => net15861, C1 => INPUT(188), C2 => n6, ZN => 
                           n21);
   U75 : AOI222_X1 port map( A1 => INPUT(118), A2 => net15843, B1 => INPUT(246)
                           , B2 => net25733, C1 => INPUT(182), C2 => net15871, 
                           ZN => n35);
   U76 : AOI222_X1 port map( A1 => INPUT(117), A2 => net15843, B1 => INPUT(245)
                           , B2 => net15865, C1 => INPUT(181), C2 => net15871, 
                           ZN => n37);
   U77 : AND3_X1 port map( A1 => n163, A2 => n164, A3 => n165, ZN => n19);
   U78 : NAND2_X1 port map( A1 => INPUT(189), A2 => n6, ZN => n163);
   U79 : NAND2_X1 port map( A1 => INPUT(253), A2 => n5, ZN => n164);
   U80 : NAND2_X1 port map( A1 => INPUT(125), A2 => n4, ZN => n165);
   U81 : AOI222_X1 port map( A1 => INPUT(109), A2 => net15849, B1 => INPUT(237)
                           , B2 => net25733, C1 => INPUT(173), C2 => net15873, 
                           ZN => n55);
   U82 : AOI222_X1 port map( A1 => INPUT(108), A2 => net15849, B1 => INPUT(236)
                           , B2 => net15865, C1 => INPUT(172), C2 => net15873, 
                           ZN => n57);
   U83 : AOI222_X1 port map( A1 => INPUT(107), A2 => net15849, B1 => INPUT(235)
                           , B2 => net15855, C1 => INPUT(171), C2 => net15873, 
                           ZN => n59);
   U84 : AOI222_X1 port map( A1 => INPUT(106), A2 => net15849, B1 => INPUT(234)
                           , B2 => net15857, C1 => INPUT(170), C2 => net15873, 
                           ZN => n61);
   U85 : AOI222_X1 port map( A1 => INPUT(96), A2 => net15847, B1 => INPUT(224),
                           B2 => net25733, C1 => INPUT(160), C2 => net15871, ZN
                           => n83);
   U86 : AOI222_X1 port map( A1 => INPUT(97), A2 => net15847, B1 => INPUT(225),
                           B2 => net25734, C1 => INPUT(161), C2 => net15871, ZN
                           => n81);
   U87 : AOI222_X1 port map( A1 => INPUT(98), A2 => net15847, B1 => INPUT(226),
                           B2 => net25733, C1 => INPUT(162), C2 => net15871, ZN
                           => n79);
   U88 : AOI222_X1 port map( A1 => INPUT(99), A2 => net15847, B1 => INPUT(227),
                           B2 => net25733, C1 => INPUT(163), C2 => net15871, ZN
                           => n77);
   U89 : AOI222_X1 port map( A1 => INPUT(100), A2 => net15847, B1 => INPUT(228)
                           , B2 => net25733, C1 => INPUT(164), C2 => net15871, 
                           ZN => n75);
   U90 : AOI222_X1 port map( A1 => INPUT(101), A2 => net15847, B1 => INPUT(229)
                           , B2 => net25734, C1 => INPUT(165), C2 => net15871, 
                           ZN => n73);
   U91 : AOI222_X1 port map( A1 => INPUT(105), A2 => net15847, B1 => INPUT(233)
                           , B2 => net15859, C1 => INPUT(169), C2 => net15871, 
                           ZN => n63);
   U92 : AOI222_X1 port map( A1 => INPUT(104), A2 => net15847, B1 => INPUT(232)
                           , B2 => net15861, C1 => INPUT(168), C2 => net15871, 
                           ZN => n65);
   U93 : AOI222_X1 port map( A1 => INPUT(103), A2 => net15847, B1 => INPUT(231)
                           , B2 => net25734, C1 => INPUT(167), C2 => net15871, 
                           ZN => n69);
   U94 : AOI222_X1 port map( A1 => INPUT(102), A2 => net15847, B1 => INPUT(230)
                           , B2 => net25734, C1 => INPUT(166), C2 => net15871, 
                           ZN => n71);
   U95 : AOI222_X1 port map( A1 => INPUT(95), A2 => net15847, B1 => INPUT(223),
                           B2 => net25734, C1 => INPUT(159), C2 => net15871, ZN
                           => n85);
   U96 : AOI222_X1 port map( A1 => INPUT(83), A2 => net15843, B1 => INPUT(211),
                           B2 => net15855, C1 => INPUT(147), C2 => net15867, ZN
                           => n113);
   U97 : AOI222_X1 port map( A1 => INPUT(82), A2 => net15843, B1 => INPUT(210),
                           B2 => net15857, C1 => INPUT(146), C2 => net15867, ZN
                           => n115);
   U98 : AOI222_X1 port map( A1 => INPUT(81), A2 => net15843, B1 => INPUT(209),
                           B2 => net15859, C1 => INPUT(145), C2 => net15867, ZN
                           => n117);
   U99 : AOI222_X1 port map( A1 => INPUT(67), A2 => net15847, B1 => INPUT(195),
                           B2 => net25733, C1 => INPUT(131), C2 => net15871, ZN
                           => n67);
   U100 : AOI222_X1 port map( A1 => INPUT(66), A2 => net15845, B1 => INPUT(194)
                           , B2 => net15865, C1 => INPUT(130), C2 => net15869, 
                           ZN => n89);
   U101 : AOI222_X1 port map( A1 => INPUT(65), A2 => net15843, B1 => INPUT(193)
                           , B2 => net15855, C1 => INPUT(129), C2 => net15867, 
                           ZN => n111);
   U102 : AOI222_X1 port map( A1 => INPUT(64), A2 => net15843, B1 => INPUT(192)
                           , B2 => net15861, C1 => INPUT(128), C2 => net15867, 
                           ZN => n133);
   U103 : AOI222_X1 port map( A1 => INPUT(126), A2 => net15843, B1 => 
                           INPUT(254), B2 => net15857, C1 => INPUT(190), C2 => 
                           net15871, ZN => n17);
   U104 : BUF_X1 port map( A => n7, Z => net15885);
   U105 : BUF_X1 port map( A => n7, Z => net15883);
   U106 : BUF_X1 port map( A => n7, Z => net15881);
   U107 : BUF_X1 port map( A => n7, Z => net15879);
   U108 : AOI222_X1 port map( A1 => INPUT(115), A2 => net15849, B1 => 
                           INPUT(243), B2 => net15857, C1 => INPUT(179), C2 => 
                           net15873, ZN => n41);
   U109 : AOI222_X1 port map( A1 => INPUT(114), A2 => net15849, B1 => 
                           INPUT(242), B2 => net15859, C1 => INPUT(178), C2 => 
                           net15873, ZN => n43);
   U110 : AOI222_X1 port map( A1 => INPUT(116), A2 => net15849, B1 => 
                           INPUT(244), B2 => net15855, C1 => INPUT(180), C2 => 
                           net15873, ZN => n39);
   U111 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(7));
   U112 : AOI222_X1 port map( A1 => INPUT(71), A2 => net15853, B1 => INPUT(199)
                           , B2 => net15857, C1 => INPUT(135), C2 => net15877, 
                           ZN => n11);
   U113 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(6));
   U114 : AOI222_X1 port map( A1 => INPUT(70), A2 => net15853, B1 => INPUT(198)
                           , B2 => net15859, C1 => INPUT(134), C2 => net15877, 
                           ZN => n13);
   U115 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(4));
   U116 : AOI222_X1 port map( A1 => INPUT(68), A2 => net15849, B1 => INPUT(196)
                           , B2 => net25734, C1 => INPUT(132), C2 => net15873, 
                           ZN => n45);
   U117 : AOI222_X1 port map( A1 => INPUT(69), A2 => net15843, B1 => INPUT(197)
                           , B2 => net15861, C1 => INPUT(133), C2 => net15871, 
                           ZN => n23);
   U118 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => Y(29));
   U119 : AOI222_X1 port map( A1 => INPUT(93), A2 => net15845, B1 => INPUT(221)
                           , B2 => net15865, C1 => INPUT(157), C2 => net15869, 
                           ZN => n91);
   U120 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => Y(28));
   U121 : AOI222_X1 port map( A1 => INPUT(92), A2 => net15845, B1 => INPUT(220)
                           , B2 => net15855, C1 => INPUT(156), C2 => net15869, 
                           ZN => n93);
   U122 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => Y(27));
   U123 : AOI222_X1 port map( A1 => INPUT(91), A2 => net15845, B1 => INPUT(219)
                           , B2 => net15857, C1 => INPUT(155), C2 => net15869, 
                           ZN => n95);
   U124 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => Y(26));
   U125 : AOI222_X1 port map( A1 => INPUT(90), A2 => net15845, B1 => INPUT(218)
                           , B2 => net15859, C1 => INPUT(154), C2 => net15869, 
                           ZN => n97);
   U126 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => Y(25));
   U127 : AOI222_X1 port map( A1 => INPUT(89), A2 => net15845, B1 => INPUT(217)
                           , B2 => net15861, C1 => INPUT(153), C2 => net15869, 
                           ZN => n99);
   U128 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => Y(24));
   U129 : AOI222_X1 port map( A1 => INPUT(88), A2 => net15845, B1 => INPUT(216)
                           , B2 => net25734, C1 => INPUT(152), C2 => net15869, 
                           ZN => n101);
   U130 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => Y(23));
   U131 : AOI222_X1 port map( A1 => INPUT(87), A2 => net15845, B1 => INPUT(215)
                           , B2 => net25733, C1 => INPUT(151), C2 => net15869, 
                           ZN => n103);
   U132 : AOI222_X1 port map( A1 => INPUT(86), A2 => net15845, B1 => INPUT(214)
                           , B2 => net25734, C1 => INPUT(150), C2 => net15869, 
                           ZN => n105);
   U133 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => Y(21));
   U134 : AOI222_X1 port map( A1 => INPUT(85), A2 => net15845, B1 => INPUT(213)
                           , B2 => net25733, C1 => INPUT(149), C2 => net15869, 
                           ZN => n107);
   U135 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => Y(30));
   U136 : AOI222_X1 port map( A1 => INPUT(94), A2 => net15845, B1 => INPUT(222)
                           , B2 => net25733, C1 => INPUT(158), C2 => net15869, 
                           ZN => n87);
   U137 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => Y(20));
   U138 : AOI222_X1 port map( A1 => INPUT(84), A2 => net15845, B1 => INPUT(212)
                           , B2 => net15865, C1 => INPUT(148), C2 => net15869, 
                           ZN => n109);
   U139 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => Y(16));
   U140 : AOI222_X1 port map( A1 => INPUT(80), A2 => net15843, B1 => INPUT(208)
                           , B2 => net15861, C1 => INPUT(144), C2 => net15867, 
                           ZN => n119);
   U141 : AOI222_X1 port map( A1 => INPUT(79), A2 => net15843, B1 => INPUT(207)
                           , B2 => net25734, C1 => INPUT(143), C2 => net15867, 
                           ZN => n121);
   U142 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => Y(14));
   U143 : AOI222_X1 port map( A1 => INPUT(78), A2 => net15843, B1 => INPUT(206)
                           , B2 => net25733, C1 => INPUT(142), C2 => net15867, 
                           ZN => n123);
   U144 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => Y(13));
   U145 : AOI222_X1 port map( A1 => INPUT(77), A2 => net15843, B1 => INPUT(205)
                           , B2 => net25734, C1 => INPUT(141), C2 => net15867, 
                           ZN => n125);
   U146 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => Y(12));
   U147 : AOI222_X1 port map( A1 => INPUT(76), A2 => net15843, B1 => INPUT(204)
                           , B2 => net25733, C1 => INPUT(140), C2 => net15867, 
                           ZN => n127);
   U148 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => Y(11));
   U149 : AOI222_X1 port map( A1 => INPUT(75), A2 => net15843, B1 => INPUT(203)
                           , B2 => net25734, C1 => INPUT(139), C2 => net15867, 
                           ZN => n129);
   U150 : AOI222_X1 port map( A1 => INPUT(74), A2 => net15843, B1 => INPUT(202)
                           , B2 => net25733, C1 => INPUT(138), C2 => net15867, 
                           ZN => n131);
   U151 : AOI222_X1 port map( A1 => INPUT(73), A2 => net15853, B1 => INPUT(201)
                           , B2 => net15865, C1 => INPUT(137), C2 => net15877, 
                           ZN => n3);
   U152 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(8));
   U153 : AOI222_X1 port map( A1 => INPUT(72), A2 => net15853, B1 => INPUT(200)
                           , B2 => net15855, C1 => INPUT(136), C2 => net15877, 
                           ZN => n9);
   U154 : AOI22_X1 port map( A1 => INPUT(51), A2 => net15885, B1 => INPUT(307),
                           B2 => net15651, ZN => n40);
   U155 : AOI22_X1 port map( A1 => INPUT(52), A2 => net15885, B1 => INPUT(308),
                           B2 => net15653, ZN => n38);
   U156 : AOI22_X1 port map( A1 => INPUT(59), A2 => net15887, B1 => INPUT(315),
                           B2 => net15653, ZN => n24);
   U157 : AOI22_X1 port map( A1 => INPUT(58), A2 => net15887, B1 => INPUT(314),
                           B2 => net15653, ZN => n26);
   U158 : AOI22_X1 port map( A1 => INPUT(57), A2 => net15887, B1 => INPUT(313),
                           B2 => net15653, ZN => n28);
   U159 : AOI22_X1 port map( A1 => INPUT(56), A2 => net15887, B1 => INPUT(312),
                           B2 => net15653, ZN => n30);
   U160 : AOI22_X1 port map( A1 => INPUT(55), A2 => net15887, B1 => INPUT(311),
                           B2 => net15653, ZN => n32);
   U161 : AOI22_X1 port map( A1 => INPUT(54), A2 => net15887, B1 => INPUT(310),
                           B2 => net15653, ZN => n34);
   U162 : AOI22_X1 port map( A1 => INPUT(50), A2 => net15885, B1 => INPUT(306),
                           B2 => net15651, ZN => n42);
   U163 : AOI22_X1 port map( A1 => INPUT(49), A2 => net15885, B1 => INPUT(305),
                           B2 => net15651, ZN => n46);
   U164 : AOI22_X1 port map( A1 => INPUT(53), A2 => net15887, B1 => INPUT(309),
                           B2 => net15653, ZN => n36);
   U165 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(3));
   U166 : AOI22_X1 port map( A1 => INPUT(3), A2 => net15883, B1 => INPUT(259), 
                           B2 => net15649, ZN => n66);
   U167 : AOI22_X1 port map( A1 => INPUT(2), A2 => net15881, B1 => INPUT(258), 
                           B2 => net15647, ZN => n88);
   U168 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => Y(1));
   U169 : AOI22_X1 port map( A1 => INPUT(1), A2 => net15879, B1 => INPUT(257), 
                           B2 => net15647, ZN => n110);
   U170 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => Y(0));
   U171 : AOI22_X1 port map( A1 => INPUT(0), A2 => net15879, B1 => INPUT(256), 
                           B2 => net15645, ZN => n132);
   U172 : AOI22_X1 port map( A1 => INPUT(19), A2 => net15879, B1 => INPUT(275),
                           B2 => net15645, ZN => n112);
   U173 : AOI22_X1 port map( A1 => INPUT(18), A2 => net15879, B1 => INPUT(274),
                           B2 => net15645, ZN => n114);
   U174 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => Y(17));
   U175 : AOI22_X1 port map( A1 => INPUT(17), A2 => net15879, B1 => INPUT(273),
                           B2 => net15645, ZN => n116);
   U176 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => Y(31));
   U177 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => Y(32));
   U178 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => Y(33));
   U179 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => Y(34));
   U180 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => Y(35));
   U181 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => Y(36));
   U182 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => Y(37));
   U183 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => Y(38));
   U184 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(39));
   U185 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(42));
   U186 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(41));
   U187 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(40));
   U188 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(56));
   U189 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(55));
   U190 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(54));
   U191 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(51));
   U192 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(50));
   U193 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(49));
   U194 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(48));
   U195 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(47));
   U196 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(46));
   U197 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(45));
   U198 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(44));
   U199 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(43));
   U200 : NAND2_X1 port map( A1 => n28, A2 => n139, ZN => Y(57));
   U201 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(58));
   U202 : AOI22_X1 port map( A1 => INPUT(31), A2 => net15883, B1 => INPUT(287),
                           B2 => net15649, ZN => n84);
   U203 : AOI22_X1 port map( A1 => INPUT(32), A2 => net15883, B1 => INPUT(288),
                           B2 => net15649, ZN => n82);
   U204 : AOI22_X1 port map( A1 => INPUT(33), A2 => net15883, B1 => INPUT(289),
                           B2 => net15649, ZN => n80);
   U205 : AOI22_X1 port map( A1 => INPUT(34), A2 => net15883, B1 => INPUT(290),
                           B2 => net15649, ZN => n78);
   U206 : AOI22_X1 port map( A1 => INPUT(35), A2 => net15883, B1 => INPUT(291),
                           B2 => net15649, ZN => n76);
   U207 : AOI22_X1 port map( A1 => INPUT(36), A2 => net15883, B1 => INPUT(292),
                           B2 => net15649, ZN => n74);
   U208 : AOI22_X1 port map( A1 => INPUT(37), A2 => net15883, B1 => INPUT(293),
                           B2 => net15649, ZN => n72);
   U209 : AOI22_X1 port map( A1 => INPUT(48), A2 => net15885, B1 => INPUT(304),
                           B2 => net15651, ZN => n48);
   U210 : AOI22_X1 port map( A1 => INPUT(47), A2 => net15885, B1 => INPUT(303),
                           B2 => net15651, ZN => n50);
   U211 : AOI22_X1 port map( A1 => INPUT(46), A2 => net15885, B1 => INPUT(302),
                           B2 => net15651, ZN => n52);
   U212 : AOI22_X1 port map( A1 => INPUT(45), A2 => net15885, B1 => INPUT(301),
                           B2 => net15651, ZN => n54);
   U213 : AOI22_X1 port map( A1 => INPUT(44), A2 => net15885, B1 => INPUT(300),
                           B2 => net15651, ZN => n56);
   U214 : AOI22_X1 port map( A1 => INPUT(43), A2 => net15885, B1 => INPUT(299),
                           B2 => net15651, ZN => n58);
   U215 : AOI22_X1 port map( A1 => INPUT(42), A2 => net15885, B1 => INPUT(298),
                           B2 => net15651, ZN => n60);
   U216 : AOI22_X1 port map( A1 => INPUT(41), A2 => net15883, B1 => INPUT(297),
                           B2 => net15651, ZN => n62);
   U217 : AOI22_X1 port map( A1 => INPUT(40), A2 => net15883, B1 => INPUT(296),
                           B2 => net15649, ZN => n64);
   U218 : AOI22_X1 port map( A1 => INPUT(39), A2 => net15883, B1 => INPUT(295),
                           B2 => net15649, ZN => n68);
   U219 : AOI22_X1 port map( A1 => INPUT(38), A2 => net15883, B1 => INPUT(294),
                           B2 => net15649, ZN => n70);
   U220 : AOI22_X1 port map( A1 => INPUT(28), A2 => net15881, B1 => INPUT(284),
                           B2 => net15647, ZN => n92);
   U221 : AOI22_X1 port map( A1 => INPUT(27), A2 => net15881, B1 => INPUT(283),
                           B2 => net15647, ZN => n94);
   U222 : AOI22_X1 port map( A1 => INPUT(26), A2 => net15881, B1 => INPUT(282),
                           B2 => net15647, ZN => n96);
   U223 : AOI22_X1 port map( A1 => INPUT(24), A2 => net15881, B1 => INPUT(280),
                           B2 => net15647, ZN => n100);
   U224 : AOI22_X1 port map( A1 => INPUT(23), A2 => net15881, B1 => INPUT(279),
                           B2 => net15647, ZN => n102);
   U225 : AOI22_X1 port map( A1 => INPUT(22), A2 => net15881, B1 => INPUT(278),
                           B2 => net15647, ZN => n104);
   U226 : AOI22_X1 port map( A1 => INPUT(20), A2 => net15881, B1 => INPUT(276),
                           B2 => net15647, ZN => n108);
   U227 : AOI22_X1 port map( A1 => INPUT(25), A2 => net15881, B1 => INPUT(281),
                           B2 => net15647, ZN => n98);
   U228 : AOI22_X1 port map( A1 => INPUT(29), A2 => net15881, B1 => INPUT(285),
                           B2 => net15647, ZN => n90);
   U229 : AOI22_X1 port map( A1 => INPUT(21), A2 => net15881, B1 => INPUT(277),
                           B2 => net15647, ZN => n106);
   U230 : AOI22_X1 port map( A1 => INPUT(30), A2 => net15881, B1 => INPUT(286),
                           B2 => net15649, ZN => n86);
   U231 : AOI22_X1 port map( A1 => INPUT(9), A2 => net15889, B1 => net15655, B2
                           => INPUT(265), ZN => n2);
   U232 : AOI22_X1 port map( A1 => INPUT(11), A2 => net15879, B1 => INPUT(267),
                           B2 => net15645, ZN => n128);
   U233 : AOI22_X1 port map( A1 => INPUT(10), A2 => net15879, B1 => INPUT(266),
                           B2 => net15645, ZN => n130);
   U234 : AOI22_X1 port map( A1 => INPUT(13), A2 => net15879, B1 => INPUT(269),
                           B2 => net15645, ZN => n124);
   U235 : AOI22_X1 port map( A1 => INPUT(12), A2 => net15879, B1 => INPUT(268),
                           B2 => net15645, ZN => n126);
   U236 : AOI22_X1 port map( A1 => INPUT(15), A2 => net15879, B1 => INPUT(271),
                           B2 => net15645, ZN => n120);
   U237 : AOI22_X1 port map( A1 => INPUT(14), A2 => net15879, B1 => INPUT(270),
                           B2 => net15645, ZN => n122);
   U238 : AOI22_X1 port map( A1 => INPUT(16), A2 => net15879, B1 => INPUT(272),
                           B2 => net15645, ZN => n118);
   U239 : AOI22_X1 port map( A1 => INPUT(7), A2 => net15889, B1 => INPUT(263), 
                           B2 => net15655, ZN => n10);
   U240 : AOI22_X1 port map( A1 => INPUT(5), A2 => net15887, B1 => INPUT(261), 
                           B2 => net15653, ZN => n22);
   U241 : AOI22_X1 port map( A1 => INPUT(4), A2 => net15885, B1 => INPUT(260), 
                           B2 => net15651, ZN => n44);
   U242 : AOI22_X1 port map( A1 => INPUT(8), A2 => net15889, B1 => INPUT(264), 
                           B2 => net15655, ZN => n8);
   U243 : AOI22_X1 port map( A1 => INPUT(6), A2 => net15889, B1 => INPUT(262), 
                           B2 => net15655, ZN => n12);
   U244 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(63));
   U245 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(62));
   U246 : AOI22_X1 port map( A1 => INPUT(63), A2 => net15887, B1 => INPUT(319),
                           B2 => net15655, ZN => n14);
   U247 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(52));
   U248 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(53));
   U249 : AOI22_X1 port map( A1 => INPUT(62), A2 => net15887, B1 => INPUT(318),
                           B2 => net15653, ZN => n16);
   U250 : AOI222_X1 port map( A1 => INPUT(127), A2 => net15843, B1 => 
                           INPUT(255), B2 => net15859, C1 => INPUT(191), C2 => 
                           net15871, ZN => n15);
   U251 : AOI22_X1 port map( A1 => INPUT(60), A2 => net15887, B1 => INPUT(316),
                           B2 => net15653, ZN => n20);
   U252 : CLKBUF_X1 port map( A => n7, Z => net15889);
   U253 : CLKBUF_X1 port map( A => n6, Z => net15877);
   U254 : CLKBUF_X1 port map( A => n5, Z => net15865);
   U255 : CLKBUF_X1 port map( A => SEL(0), Z => net15655);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_15 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_15;

architecture SYN_Behavior of Shifter_NBIT64_15 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_16 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_16;

architecture SYN_Behavior of Shifter_NBIT64_16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Shifter_NBIT64_0 is

   port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
         std_logic_vector (127 downto 0));

end Shifter_NBIT64_0;

architecture SYN_Behavior of Shifter_NBIT64_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, RESULT_1_48_port : std_logic;

begin
   RESULT <= ( TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port, X_Logic0_port, 
      TO_SHIFT(62), TO_SHIFT(61), TO_SHIFT(60), TO_SHIFT(59), TO_SHIFT(58), 
      TO_SHIFT(57), TO_SHIFT(56), TO_SHIFT(55), TO_SHIFT(54), TO_SHIFT(53), 
      TO_SHIFT(52), TO_SHIFT(51), TO_SHIFT(50), TO_SHIFT(49), TO_SHIFT(48), 
      TO_SHIFT(47), RESULT_1_48_port, TO_SHIFT(45), TO_SHIFT(44), TO_SHIFT(43),
      TO_SHIFT(42), TO_SHIFT(41), TO_SHIFT(40), TO_SHIFT(39), TO_SHIFT(38), 
      TO_SHIFT(37), TO_SHIFT(36), TO_SHIFT(35), TO_SHIFT(34), TO_SHIFT(33), 
      TO_SHIFT(32), TO_SHIFT(31), TO_SHIFT(30), TO_SHIFT(29), TO_SHIFT(28), 
      TO_SHIFT(27), TO_SHIFT(26), TO_SHIFT(25), TO_SHIFT(24), TO_SHIFT(23), 
      TO_SHIFT(22), TO_SHIFT(21), TO_SHIFT(20), TO_SHIFT(19), TO_SHIFT(18), 
      TO_SHIFT(17), TO_SHIFT(16), TO_SHIFT(15), TO_SHIFT(14), TO_SHIFT(13), 
      TO_SHIFT(12), TO_SHIFT(11), TO_SHIFT(10), TO_SHIFT(9), TO_SHIFT(8), 
      TO_SHIFT(7), TO_SHIFT(6), TO_SHIFT(5), TO_SHIFT(4), TO_SHIFT(3), 
      TO_SHIFT(2), TO_SHIFT(1), TO_SHIFT(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => TO_SHIFT(46), Z => RESULT_1_48_port);

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity Booth_Encoder_0 is

   port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
         std_logic_vector (2 downto 0));

end Booth_Encoder_0;

architecture SYN_Behavior of Booth_Encoder_0 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n3);
   U2 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n3, ZN => n5);
   U3 : OAI22_X1 port map( A1 => n5, A2 => n6, B1 => B(2), B2 => n3, ZN => 
                           OUT_TO_MUX(1));
   U4 : INV_X1 port map( A => B(2), ZN => n6);
   U5 : AOI21_X1 port map( B1 => n2, B2 => n3, A => B(2), ZN => OUT_TO_MUX(0));
   U6 : OAI21_X1 port map( B1 => B(1), B2 => B(0), A => n3, ZN => n2);
   U7 : AND3_X1 port map( A1 => B(2), A2 => n3, A3 => n5, ZN => OUT_TO_MUX(2));

end SYN_Behavior;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BOOTHMUL is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL;

architecture SYN_STRUCTURAL of BOOTHMUL is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component RCA_NBIT64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_1
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_2
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_3
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_4
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_5
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_6
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_7
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_8
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_9
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_10
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_11
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_12
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_13
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_14
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_15
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_0
      port( INPUT : in std_logic_vector (0 to 319);  SEL : in std_logic_vector 
            (0 to 2);  Y : out std_logic_vector (0 to 63));
   end component;
   
   component Shifter_NBIT64_1
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_2
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_3
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_4
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_5
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_6
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_7
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_8
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_9
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_10
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_11
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_12
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_13
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_14
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_15
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_16
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_17
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_18
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_19
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_20
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_21
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_22
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_23
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_24
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_25
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_26
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_27
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_28
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_29
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_30
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_31
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Shifter_NBIT64_0
      port( TO_SHIFT : in std_logic_vector (63 downto 0);  RESULT : out 
            std_logic_vector (127 downto 0));
   end component;
   
   component Booth_Encoder_1
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_2
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_3
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_4
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_5
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_6
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_7
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_8
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_9
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_10
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_11
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_12
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_13
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_14
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_15
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component Booth_Encoder_0
      port( B : in std_logic_vector (2 downto 0);  OUT_TO_MUX : out 
            std_logic_vector (2 downto 0));
   end component;
   
   signal X_Logic0_port, A_neg_tmp_63_port, A_neg_tmp_31_port, 
      A_neg_tmp_30_port, A_neg_tmp_29_port, A_neg_tmp_28_port, 
      A_neg_tmp_27_port, A_neg_tmp_26_port, A_neg_tmp_25_port, 
      A_neg_tmp_24_port, A_neg_tmp_23_port, A_neg_tmp_22_port, 
      A_neg_tmp_21_port, A_neg_tmp_20_port, A_neg_tmp_19_port, 
      A_neg_tmp_18_port, A_neg_tmp_17_port, A_neg_tmp_16_port, 
      A_neg_tmp_15_port, A_neg_tmp_14_port, A_neg_tmp_13_port, 
      A_neg_tmp_12_port, A_neg_tmp_11_port, A_neg_tmp_10_port, A_neg_tmp_9_port
      , A_neg_tmp_8_port, A_neg_tmp_7_port, A_neg_tmp_6_port, A_neg_tmp_5_port,
      A_neg_tmp_4_port, A_neg_tmp_3_port, A_neg_tmp_2_port, A_neg_tmp_1_port, 
      A_neg_tmp_0_port, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, 
      N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91
      , N92, N93, N94, N95, N96, N97, selection_signal_0_2_port, 
      selection_signal_0_1_port, selection_signal_0_0_port, 
      selection_signal_1_2_port, selection_signal_1_1_port, 
      selection_signal_1_0_port, selection_signal_2_2_port, 
      selection_signal_2_1_port, selection_signal_2_0_port, 
      selection_signal_3_2_port, selection_signal_3_1_port, 
      selection_signal_3_0_port, selection_signal_4_2_port, 
      selection_signal_4_1_port, selection_signal_4_0_port, 
      selection_signal_5_2_port, selection_signal_5_1_port, 
      selection_signal_5_0_port, selection_signal_6_2_port, 
      selection_signal_6_1_port, selection_signal_6_0_port, 
      selection_signal_7_2_port, selection_signal_7_1_port, 
      selection_signal_7_0_port, selection_signal_8_2_port, 
      selection_signal_8_1_port, selection_signal_8_0_port, 
      selection_signal_9_2_port, selection_signal_9_1_port, 
      selection_signal_9_0_port, selection_signal_10_2_port, 
      selection_signal_10_1_port, selection_signal_10_0_port, 
      selection_signal_11_2_port, selection_signal_11_1_port, 
      selection_signal_11_0_port, selection_signal_12_2_port, 
      selection_signal_12_1_port, selection_signal_12_0_port, 
      selection_signal_13_2_port, selection_signal_13_1_port, 
      selection_signal_13_0_port, selection_signal_14_2_port, 
      selection_signal_14_1_port, selection_signal_14_0_port, 
      selection_signal_15_2_port, selection_signal_15_1_port, 
      selection_signal_15_0_port, A_pos_shifted_by1_0_63_port, 
      A_pos_shifted_by1_0_62_port, A_pos_shifted_by1_0_61_port, 
      A_pos_shifted_by1_0_60_port, A_pos_shifted_by1_0_59_port, 
      A_pos_shifted_by1_0_58_port, A_pos_shifted_by1_0_57_port, 
      A_pos_shifted_by1_0_56_port, A_pos_shifted_by1_0_55_port, 
      A_pos_shifted_by1_0_54_port, A_pos_shifted_by1_0_53_port, 
      A_pos_shifted_by1_0_52_port, A_pos_shifted_by1_0_51_port, 
      A_pos_shifted_by1_0_50_port, A_pos_shifted_by1_0_49_port, 
      A_pos_shifted_by1_0_48_port, A_pos_shifted_by1_0_47_port, 
      A_pos_shifted_by1_0_46_port, A_pos_shifted_by1_0_45_port, 
      A_pos_shifted_by1_0_44_port, A_pos_shifted_by1_0_43_port, 
      A_pos_shifted_by1_0_42_port, A_pos_shifted_by1_0_41_port, 
      A_pos_shifted_by1_0_40_port, A_pos_shifted_by1_0_39_port, 
      A_pos_shifted_by1_0_38_port, A_pos_shifted_by1_0_37_port, 
      A_pos_shifted_by1_0_36_port, A_pos_shifted_by1_0_35_port, 
      A_pos_shifted_by1_0_34_port, A_pos_shifted_by1_0_33_port, 
      A_pos_shifted_by1_0_32_port, A_pos_shifted_by1_0_31_port, 
      A_pos_shifted_by1_0_30_port, A_pos_shifted_by1_0_29_port, 
      A_pos_shifted_by1_0_28_port, A_pos_shifted_by1_0_27_port, 
      A_pos_shifted_by1_0_26_port, A_pos_shifted_by1_0_25_port, 
      A_pos_shifted_by1_0_24_port, A_pos_shifted_by1_0_23_port, 
      A_pos_shifted_by1_0_22_port, A_pos_shifted_by1_0_21_port, 
      A_pos_shifted_by1_0_20_port, A_pos_shifted_by1_0_19_port, 
      A_pos_shifted_by1_0_18_port, A_pos_shifted_by1_0_17_port, 
      A_pos_shifted_by1_0_16_port, A_pos_shifted_by1_0_15_port, 
      A_pos_shifted_by1_0_14_port, A_pos_shifted_by1_0_13_port, 
      A_pos_shifted_by1_0_12_port, A_pos_shifted_by1_0_11_port, 
      A_pos_shifted_by1_0_10_port, A_pos_shifted_by1_0_9_port, 
      A_pos_shifted_by1_0_8_port, A_pos_shifted_by1_0_7_port, 
      A_pos_shifted_by1_0_6_port, A_pos_shifted_by1_0_5_port, 
      A_pos_shifted_by1_0_4_port, A_pos_shifted_by1_0_3_port, 
      A_pos_shifted_by1_0_2_port, A_pos_shifted_by1_0_1_port, 
      A_pos_shifted_by1_0_0_port, A_pos_shifted_by1_1_63_port, 
      A_pos_shifted_by1_1_62_port, A_pos_shifted_by1_1_61_port, 
      A_pos_shifted_by1_1_60_port, A_pos_shifted_by1_1_59_port, 
      A_pos_shifted_by1_1_58_port, A_pos_shifted_by1_1_57_port, 
      A_pos_shifted_by1_1_56_port, A_pos_shifted_by1_1_55_port, 
      A_pos_shifted_by1_1_54_port, A_pos_shifted_by1_1_53_port, 
      A_pos_shifted_by1_1_52_port, A_pos_shifted_by1_1_51_port, 
      A_pos_shifted_by1_1_50_port, A_pos_shifted_by1_1_49_port, 
      A_pos_shifted_by1_1_48_port, A_pos_shifted_by1_1_47_port, 
      A_pos_shifted_by1_1_46_port, A_pos_shifted_by1_1_45_port, 
      A_pos_shifted_by1_1_44_port, A_pos_shifted_by1_1_43_port, 
      A_pos_shifted_by1_1_42_port, A_pos_shifted_by1_1_41_port, 
      A_pos_shifted_by1_1_40_port, A_pos_shifted_by1_1_39_port, 
      A_pos_shifted_by1_1_38_port, A_pos_shifted_by1_1_37_port, 
      A_pos_shifted_by1_1_36_port, A_pos_shifted_by1_1_35_port, 
      A_pos_shifted_by1_1_34_port, A_pos_shifted_by1_1_33_port, 
      A_pos_shifted_by1_1_32_port, A_pos_shifted_by1_1_31_port, 
      A_pos_shifted_by1_1_30_port, A_pos_shifted_by1_1_29_port, 
      A_pos_shifted_by1_1_28_port, A_pos_shifted_by1_1_27_port, 
      A_pos_shifted_by1_1_26_port, A_pos_shifted_by1_1_25_port, 
      A_pos_shifted_by1_1_24_port, A_pos_shifted_by1_1_23_port, 
      A_pos_shifted_by1_1_22_port, A_pos_shifted_by1_1_21_port, 
      A_pos_shifted_by1_1_20_port, A_pos_shifted_by1_1_19_port, 
      A_pos_shifted_by1_1_18_port, A_pos_shifted_by1_1_17_port, 
      A_pos_shifted_by1_1_16_port, A_pos_shifted_by1_1_15_port, 
      A_pos_shifted_by1_1_14_port, A_pos_shifted_by1_1_13_port, 
      A_pos_shifted_by1_1_12_port, A_pos_shifted_by1_1_11_port, 
      A_pos_shifted_by1_1_10_port, A_pos_shifted_by1_1_9_port, 
      A_pos_shifted_by1_1_8_port, A_pos_shifted_by1_1_7_port, 
      A_pos_shifted_by1_1_6_port, A_pos_shifted_by1_1_5_port, 
      A_pos_shifted_by1_1_4_port, A_pos_shifted_by1_1_3_port, 
      A_pos_shifted_by1_1_2_port, A_pos_shifted_by1_1_1_port, 
      A_pos_shifted_by1_1_0_port, A_pos_shifted_by1_2_63_port, 
      A_pos_shifted_by1_2_62_port, A_pos_shifted_by1_2_61_port, 
      A_pos_shifted_by1_2_60_port, A_pos_shifted_by1_2_59_port, 
      A_pos_shifted_by1_2_58_port, A_pos_shifted_by1_2_57_port, 
      A_pos_shifted_by1_2_56_port, A_pos_shifted_by1_2_55_port, 
      A_pos_shifted_by1_2_54_port, A_pos_shifted_by1_2_53_port, 
      A_pos_shifted_by1_2_52_port, A_pos_shifted_by1_2_51_port, 
      A_pos_shifted_by1_2_50_port, A_pos_shifted_by1_2_49_port, 
      A_pos_shifted_by1_2_48_port, A_pos_shifted_by1_2_47_port, 
      A_pos_shifted_by1_2_46_port, A_pos_shifted_by1_2_45_port, 
      A_pos_shifted_by1_2_44_port, A_pos_shifted_by1_2_43_port, 
      A_pos_shifted_by1_2_42_port, A_pos_shifted_by1_2_41_port, 
      A_pos_shifted_by1_2_40_port, A_pos_shifted_by1_2_39_port, 
      A_pos_shifted_by1_2_38_port, A_pos_shifted_by1_2_37_port, 
      A_pos_shifted_by1_2_36_port, A_pos_shifted_by1_2_35_port, 
      A_pos_shifted_by1_2_34_port, A_pos_shifted_by1_2_33_port, 
      A_pos_shifted_by1_2_32_port, A_pos_shifted_by1_2_31_port, 
      A_pos_shifted_by1_2_30_port, A_pos_shifted_by1_2_29_port, 
      A_pos_shifted_by1_2_28_port, A_pos_shifted_by1_2_27_port, 
      A_pos_shifted_by1_2_26_port, A_pos_shifted_by1_2_25_port, 
      A_pos_shifted_by1_2_24_port, A_pos_shifted_by1_2_23_port, 
      A_pos_shifted_by1_2_22_port, A_pos_shifted_by1_2_21_port, 
      A_pos_shifted_by1_2_20_port, A_pos_shifted_by1_2_19_port, 
      A_pos_shifted_by1_2_18_port, A_pos_shifted_by1_2_17_port, 
      A_pos_shifted_by1_2_16_port, A_pos_shifted_by1_2_15_port, 
      A_pos_shifted_by1_2_14_port, A_pos_shifted_by1_2_13_port, 
      A_pos_shifted_by1_2_12_port, A_pos_shifted_by1_2_11_port, 
      A_pos_shifted_by1_2_10_port, A_pos_shifted_by1_2_9_port, 
      A_pos_shifted_by1_2_8_port, A_pos_shifted_by1_2_7_port, 
      A_pos_shifted_by1_2_6_port, A_pos_shifted_by1_2_5_port, 
      A_pos_shifted_by1_2_4_port, A_pos_shifted_by1_2_3_port, 
      A_pos_shifted_by1_2_2_port, A_pos_shifted_by1_2_1_port, 
      A_pos_shifted_by1_2_0_port, A_pos_shifted_by1_3_63_port, 
      A_pos_shifted_by1_3_62_port, A_pos_shifted_by1_3_61_port, 
      A_pos_shifted_by1_3_60_port, A_pos_shifted_by1_3_59_port, 
      A_pos_shifted_by1_3_58_port, A_pos_shifted_by1_3_57_port, 
      A_pos_shifted_by1_3_56_port, A_pos_shifted_by1_3_55_port, 
      A_pos_shifted_by1_3_54_port, A_pos_shifted_by1_3_53_port, 
      A_pos_shifted_by1_3_52_port, A_pos_shifted_by1_3_51_port, 
      A_pos_shifted_by1_3_50_port, A_pos_shifted_by1_3_49_port, 
      A_pos_shifted_by1_3_48_port, A_pos_shifted_by1_3_47_port, 
      A_pos_shifted_by1_3_46_port, A_pos_shifted_by1_3_45_port, 
      A_pos_shifted_by1_3_44_port, A_pos_shifted_by1_3_43_port, 
      A_pos_shifted_by1_3_42_port, A_pos_shifted_by1_3_41_port, 
      A_pos_shifted_by1_3_40_port, A_pos_shifted_by1_3_39_port, 
      A_pos_shifted_by1_3_38_port, A_pos_shifted_by1_3_37_port, 
      A_pos_shifted_by1_3_36_port, A_pos_shifted_by1_3_35_port, 
      A_pos_shifted_by1_3_34_port, A_pos_shifted_by1_3_33_port, 
      A_pos_shifted_by1_3_32_port, A_pos_shifted_by1_3_31_port, 
      A_pos_shifted_by1_3_30_port, A_pos_shifted_by1_3_29_port, 
      A_pos_shifted_by1_3_28_port, A_pos_shifted_by1_3_27_port, 
      A_pos_shifted_by1_3_26_port, A_pos_shifted_by1_3_25_port, 
      A_pos_shifted_by1_3_24_port, A_pos_shifted_by1_3_23_port, 
      A_pos_shifted_by1_3_22_port, A_pos_shifted_by1_3_21_port, 
      A_pos_shifted_by1_3_20_port, A_pos_shifted_by1_3_19_port, 
      A_pos_shifted_by1_3_18_port, A_pos_shifted_by1_3_17_port, 
      A_pos_shifted_by1_3_16_port, A_pos_shifted_by1_3_15_port, 
      A_pos_shifted_by1_3_14_port, A_pos_shifted_by1_3_13_port, 
      A_pos_shifted_by1_3_12_port, A_pos_shifted_by1_3_11_port, 
      A_pos_shifted_by1_3_10_port, A_pos_shifted_by1_3_9_port, 
      A_pos_shifted_by1_3_8_port, A_pos_shifted_by1_3_7_port, 
      A_pos_shifted_by1_3_6_port, A_pos_shifted_by1_3_5_port, 
      A_pos_shifted_by1_3_4_port, A_pos_shifted_by1_3_3_port, 
      A_pos_shifted_by1_3_2_port, A_pos_shifted_by1_3_1_port, 
      A_pos_shifted_by1_3_0_port, A_pos_shifted_by1_4_63_port, 
      A_pos_shifted_by1_4_62_port, A_pos_shifted_by1_4_61_port, 
      A_pos_shifted_by1_4_60_port, A_pos_shifted_by1_4_59_port, 
      A_pos_shifted_by1_4_58_port, A_pos_shifted_by1_4_57_port, 
      A_pos_shifted_by1_4_56_port, A_pos_shifted_by1_4_55_port, 
      A_pos_shifted_by1_4_54_port, A_pos_shifted_by1_4_53_port, 
      A_pos_shifted_by1_4_52_port, A_pos_shifted_by1_4_51_port, 
      A_pos_shifted_by1_4_50_port, A_pos_shifted_by1_4_49_port, 
      A_pos_shifted_by1_4_48_port, A_pos_shifted_by1_4_47_port, 
      A_pos_shifted_by1_4_46_port, A_pos_shifted_by1_4_45_port, 
      A_pos_shifted_by1_4_44_port, A_pos_shifted_by1_4_43_port, 
      A_pos_shifted_by1_4_42_port, A_pos_shifted_by1_4_41_port, 
      A_pos_shifted_by1_4_40_port, A_pos_shifted_by1_4_39_port, 
      A_pos_shifted_by1_4_38_port, A_pos_shifted_by1_4_37_port, 
      A_pos_shifted_by1_4_36_port, A_pos_shifted_by1_4_35_port, 
      A_pos_shifted_by1_4_34_port, A_pos_shifted_by1_4_33_port, 
      A_pos_shifted_by1_4_32_port, A_pos_shifted_by1_4_31_port, 
      A_pos_shifted_by1_4_30_port, A_pos_shifted_by1_4_29_port, 
      A_pos_shifted_by1_4_28_port, A_pos_shifted_by1_4_27_port, 
      A_pos_shifted_by1_4_26_port, A_pos_shifted_by1_4_25_port, 
      A_pos_shifted_by1_4_24_port, A_pos_shifted_by1_4_23_port, 
      A_pos_shifted_by1_4_22_port, A_pos_shifted_by1_4_21_port, 
      A_pos_shifted_by1_4_20_port, A_pos_shifted_by1_4_19_port, 
      A_pos_shifted_by1_4_18_port, A_pos_shifted_by1_4_17_port, 
      A_pos_shifted_by1_4_16_port, A_pos_shifted_by1_4_15_port, 
      A_pos_shifted_by1_4_14_port, A_pos_shifted_by1_4_13_port, 
      A_pos_shifted_by1_4_12_port, A_pos_shifted_by1_4_11_port, 
      A_pos_shifted_by1_4_10_port, A_pos_shifted_by1_4_9_port, 
      A_pos_shifted_by1_4_8_port, A_pos_shifted_by1_4_7_port, 
      A_pos_shifted_by1_4_6_port, A_pos_shifted_by1_4_5_port, 
      A_pos_shifted_by1_4_4_port, A_pos_shifted_by1_4_3_port, 
      A_pos_shifted_by1_4_2_port, A_pos_shifted_by1_4_1_port, 
      A_pos_shifted_by1_4_0_port, A_pos_shifted_by1_5_63_port, 
      A_pos_shifted_by1_5_62_port, A_pos_shifted_by1_5_61_port, 
      A_pos_shifted_by1_5_60_port, A_pos_shifted_by1_5_59_port, 
      A_pos_shifted_by1_5_58_port, A_pos_shifted_by1_5_57_port, 
      A_pos_shifted_by1_5_56_port, A_pos_shifted_by1_5_55_port, 
      A_pos_shifted_by1_5_54_port, A_pos_shifted_by1_5_53_port, 
      A_pos_shifted_by1_5_52_port, A_pos_shifted_by1_5_51_port, 
      A_pos_shifted_by1_5_50_port, A_pos_shifted_by1_5_49_port, 
      A_pos_shifted_by1_5_48_port, A_pos_shifted_by1_5_47_port, 
      A_pos_shifted_by1_5_46_port, A_pos_shifted_by1_5_45_port, 
      A_pos_shifted_by1_5_44_port, A_pos_shifted_by1_5_43_port, 
      A_pos_shifted_by1_5_42_port, A_pos_shifted_by1_5_41_port, 
      A_pos_shifted_by1_5_40_port, A_pos_shifted_by1_5_39_port, 
      A_pos_shifted_by1_5_38_port, A_pos_shifted_by1_5_37_port, 
      A_pos_shifted_by1_5_36_port, A_pos_shifted_by1_5_35_port, 
      A_pos_shifted_by1_5_34_port, A_pos_shifted_by1_5_33_port, 
      A_pos_shifted_by1_5_32_port, A_pos_shifted_by1_5_31_port, 
      A_pos_shifted_by1_5_30_port, A_pos_shifted_by1_5_29_port, 
      A_pos_shifted_by1_5_28_port, A_pos_shifted_by1_5_27_port, 
      A_pos_shifted_by1_5_26_port, A_pos_shifted_by1_5_25_port, 
      A_pos_shifted_by1_5_24_port, A_pos_shifted_by1_5_23_port, 
      A_pos_shifted_by1_5_22_port, A_pos_shifted_by1_5_21_port, 
      A_pos_shifted_by1_5_20_port, A_pos_shifted_by1_5_19_port, 
      A_pos_shifted_by1_5_18_port, A_pos_shifted_by1_5_17_port, 
      A_pos_shifted_by1_5_16_port, A_pos_shifted_by1_5_15_port, 
      A_pos_shifted_by1_5_14_port, A_pos_shifted_by1_5_13_port, 
      A_pos_shifted_by1_5_12_port, A_pos_shifted_by1_5_11_port, 
      A_pos_shifted_by1_5_10_port, A_pos_shifted_by1_5_9_port, 
      A_pos_shifted_by1_5_8_port, A_pos_shifted_by1_5_7_port, 
      A_pos_shifted_by1_5_6_port, A_pos_shifted_by1_5_5_port, 
      A_pos_shifted_by1_5_4_port, A_pos_shifted_by1_5_3_port, 
      A_pos_shifted_by1_5_2_port, A_pos_shifted_by1_5_1_port, 
      A_pos_shifted_by1_5_0_port, A_pos_shifted_by1_6_63_port, 
      A_pos_shifted_by1_6_62_port, A_pos_shifted_by1_6_61_port, 
      A_pos_shifted_by1_6_60_port, A_pos_shifted_by1_6_59_port, 
      A_pos_shifted_by1_6_58_port, A_pos_shifted_by1_6_57_port, 
      A_pos_shifted_by1_6_56_port, A_pos_shifted_by1_6_55_port, 
      A_pos_shifted_by1_6_54_port, A_pos_shifted_by1_6_53_port, 
      A_pos_shifted_by1_6_52_port, A_pos_shifted_by1_6_51_port, 
      A_pos_shifted_by1_6_50_port, A_pos_shifted_by1_6_49_port, 
      A_pos_shifted_by1_6_48_port, A_pos_shifted_by1_6_47_port, 
      A_pos_shifted_by1_6_46_port, A_pos_shifted_by1_6_45_port, 
      A_pos_shifted_by1_6_44_port, A_pos_shifted_by1_6_43_port, 
      A_pos_shifted_by1_6_42_port, A_pos_shifted_by1_6_41_port, 
      A_pos_shifted_by1_6_40_port, A_pos_shifted_by1_6_39_port, 
      A_pos_shifted_by1_6_38_port, A_pos_shifted_by1_6_37_port, 
      A_pos_shifted_by1_6_36_port, A_pos_shifted_by1_6_35_port, 
      A_pos_shifted_by1_6_34_port, A_pos_shifted_by1_6_33_port, 
      A_pos_shifted_by1_6_32_port, A_pos_shifted_by1_6_31_port, 
      A_pos_shifted_by1_6_30_port, A_pos_shifted_by1_6_29_port, 
      A_pos_shifted_by1_6_28_port, A_pos_shifted_by1_6_27_port, 
      A_pos_shifted_by1_6_26_port, A_pos_shifted_by1_6_25_port, 
      A_pos_shifted_by1_6_24_port, A_pos_shifted_by1_6_23_port, 
      A_pos_shifted_by1_6_22_port, A_pos_shifted_by1_6_21_port, 
      A_pos_shifted_by1_6_20_port, A_pos_shifted_by1_6_19_port, 
      A_pos_shifted_by1_6_18_port, A_pos_shifted_by1_6_17_port, 
      A_pos_shifted_by1_6_16_port, A_pos_shifted_by1_6_15_port, 
      A_pos_shifted_by1_6_14_port, A_pos_shifted_by1_6_13_port, 
      A_pos_shifted_by1_6_12_port, A_pos_shifted_by1_6_11_port, 
      A_pos_shifted_by1_6_10_port, A_pos_shifted_by1_6_9_port, 
      A_pos_shifted_by1_6_8_port, A_pos_shifted_by1_6_7_port, 
      A_pos_shifted_by1_6_6_port, A_pos_shifted_by1_6_5_port, 
      A_pos_shifted_by1_6_4_port, A_pos_shifted_by1_6_3_port, 
      A_pos_shifted_by1_6_2_port, A_pos_shifted_by1_6_1_port, 
      A_pos_shifted_by1_6_0_port, A_pos_shifted_by1_7_63_port, 
      A_pos_shifted_by1_7_62_port, A_pos_shifted_by1_7_61_port, 
      A_pos_shifted_by1_7_60_port, A_pos_shifted_by1_7_59_port, 
      A_pos_shifted_by1_7_58_port, A_pos_shifted_by1_7_57_port, 
      A_pos_shifted_by1_7_56_port, A_pos_shifted_by1_7_55_port, 
      A_pos_shifted_by1_7_54_port, A_pos_shifted_by1_7_53_port, 
      A_pos_shifted_by1_7_52_port, A_pos_shifted_by1_7_51_port, 
      A_pos_shifted_by1_7_50_port, A_pos_shifted_by1_7_49_port, 
      A_pos_shifted_by1_7_48_port, A_pos_shifted_by1_7_47_port, 
      A_pos_shifted_by1_7_46_port, A_pos_shifted_by1_7_45_port, 
      A_pos_shifted_by1_7_44_port, A_pos_shifted_by1_7_43_port, 
      A_pos_shifted_by1_7_42_port, A_pos_shifted_by1_7_41_port, 
      A_pos_shifted_by1_7_40_port, A_pos_shifted_by1_7_39_port, 
      A_pos_shifted_by1_7_38_port, A_pos_shifted_by1_7_37_port, 
      A_pos_shifted_by1_7_36_port, A_pos_shifted_by1_7_35_port, 
      A_pos_shifted_by1_7_34_port, A_pos_shifted_by1_7_33_port, 
      A_pos_shifted_by1_7_32_port, A_pos_shifted_by1_7_31_port, 
      A_pos_shifted_by1_7_30_port, A_pos_shifted_by1_7_29_port, 
      A_pos_shifted_by1_7_28_port, A_pos_shifted_by1_7_27_port, 
      A_pos_shifted_by1_7_26_port, A_pos_shifted_by1_7_25_port, 
      A_pos_shifted_by1_7_24_port, A_pos_shifted_by1_7_23_port, 
      A_pos_shifted_by1_7_22_port, A_pos_shifted_by1_7_21_port, 
      A_pos_shifted_by1_7_20_port, A_pos_shifted_by1_7_19_port, 
      A_pos_shifted_by1_7_18_port, A_pos_shifted_by1_7_17_port, 
      A_pos_shifted_by1_7_16_port, A_pos_shifted_by1_7_15_port, 
      A_pos_shifted_by1_7_14_port, A_pos_shifted_by1_7_13_port, 
      A_pos_shifted_by1_7_12_port, A_pos_shifted_by1_7_11_port, 
      A_pos_shifted_by1_7_10_port, A_pos_shifted_by1_7_9_port, 
      A_pos_shifted_by1_7_8_port, A_pos_shifted_by1_7_7_port, 
      A_pos_shifted_by1_7_6_port, A_pos_shifted_by1_7_5_port, 
      A_pos_shifted_by1_7_4_port, A_pos_shifted_by1_7_3_port, 
      A_pos_shifted_by1_7_2_port, A_pos_shifted_by1_7_1_port, 
      A_pos_shifted_by1_7_0_port, A_pos_shifted_by2_0_63_port, 
      A_pos_shifted_by2_0_62_port, A_pos_shifted_by2_0_61_port, 
      A_pos_shifted_by2_0_60_port, A_pos_shifted_by2_0_59_port, 
      A_pos_shifted_by2_0_58_port, A_pos_shifted_by2_0_57_port, 
      A_pos_shifted_by2_0_56_port, A_pos_shifted_by2_0_55_port, 
      A_pos_shifted_by2_0_54_port, A_pos_shifted_by2_0_53_port, 
      A_pos_shifted_by2_0_52_port, A_pos_shifted_by2_0_51_port, 
      A_pos_shifted_by2_0_50_port, A_pos_shifted_by2_0_49_port, 
      A_pos_shifted_by2_0_48_port, A_pos_shifted_by2_0_47_port, 
      A_pos_shifted_by2_0_46_port, A_pos_shifted_by2_0_45_port, 
      A_pos_shifted_by2_0_44_port, A_pos_shifted_by2_0_43_port, 
      A_pos_shifted_by2_0_42_port, A_pos_shifted_by2_0_41_port, 
      A_pos_shifted_by2_0_40_port, A_pos_shifted_by2_0_39_port, 
      A_pos_shifted_by2_0_38_port, A_pos_shifted_by2_0_37_port, 
      A_pos_shifted_by2_0_36_port, A_pos_shifted_by2_0_35_port, 
      A_pos_shifted_by2_0_34_port, A_pos_shifted_by2_0_33_port, 
      A_pos_shifted_by2_0_32_port, A_pos_shifted_by2_0_31_port, 
      A_pos_shifted_by2_0_30_port, A_pos_shifted_by2_0_29_port, 
      A_pos_shifted_by2_0_28_port, A_pos_shifted_by2_0_27_port, 
      A_pos_shifted_by2_0_26_port, A_pos_shifted_by2_0_25_port, 
      A_pos_shifted_by2_0_24_port, A_pos_shifted_by2_0_23_port, 
      A_pos_shifted_by2_0_22_port, A_pos_shifted_by2_0_21_port, 
      A_pos_shifted_by2_0_20_port, A_pos_shifted_by2_0_19_port, 
      A_pos_shifted_by2_0_18_port, A_pos_shifted_by2_0_17_port, 
      A_pos_shifted_by2_0_16_port, A_pos_shifted_by2_0_15_port, 
      A_pos_shifted_by2_0_14_port, A_pos_shifted_by2_0_13_port, 
      A_pos_shifted_by2_0_12_port, A_pos_shifted_by2_0_11_port, 
      A_pos_shifted_by2_0_10_port, A_pos_shifted_by2_0_9_port, 
      A_pos_shifted_by2_0_8_port, A_pos_shifted_by2_0_7_port, 
      A_pos_shifted_by2_0_6_port, A_pos_shifted_by2_0_5_port, 
      A_pos_shifted_by2_0_4_port, A_pos_shifted_by2_0_3_port, 
      A_pos_shifted_by2_0_2_port, A_pos_shifted_by2_0_1_port, 
      A_pos_shifted_by2_0_0_port, A_pos_shifted_by2_1_63_port, 
      A_pos_shifted_by2_1_62_port, A_pos_shifted_by2_1_61_port, 
      A_pos_shifted_by2_1_60_port, A_pos_shifted_by2_1_59_port, 
      A_pos_shifted_by2_1_58_port, A_pos_shifted_by2_1_57_port, 
      A_pos_shifted_by2_1_56_port, A_pos_shifted_by2_1_55_port, 
      A_pos_shifted_by2_1_54_port, A_pos_shifted_by2_1_53_port, 
      A_pos_shifted_by2_1_52_port, A_pos_shifted_by2_1_51_port, 
      A_pos_shifted_by2_1_50_port, A_pos_shifted_by2_1_49_port, 
      A_pos_shifted_by2_1_48_port, A_pos_shifted_by2_1_47_port, 
      A_pos_shifted_by2_1_46_port, A_pos_shifted_by2_1_45_port, 
      A_pos_shifted_by2_1_44_port, A_pos_shifted_by2_1_43_port, 
      A_pos_shifted_by2_1_42_port, A_pos_shifted_by2_1_41_port, 
      A_pos_shifted_by2_1_40_port, A_pos_shifted_by2_1_39_port, 
      A_pos_shifted_by2_1_38_port, A_pos_shifted_by2_1_37_port, 
      A_pos_shifted_by2_1_36_port, A_pos_shifted_by2_1_35_port, 
      A_pos_shifted_by2_1_34_port, A_pos_shifted_by2_1_33_port, 
      A_pos_shifted_by2_1_32_port, A_pos_shifted_by2_1_31_port, 
      A_pos_shifted_by2_1_30_port, A_pos_shifted_by2_1_29_port, 
      A_pos_shifted_by2_1_28_port, A_pos_shifted_by2_1_27_port, 
      A_pos_shifted_by2_1_26_port, A_pos_shifted_by2_1_25_port, 
      A_pos_shifted_by2_1_24_port, A_pos_shifted_by2_1_23_port, 
      A_pos_shifted_by2_1_22_port, A_pos_shifted_by2_1_21_port, 
      A_pos_shifted_by2_1_20_port, A_pos_shifted_by2_1_19_port, 
      A_pos_shifted_by2_1_18_port, A_pos_shifted_by2_1_17_port, 
      A_pos_shifted_by2_1_16_port, A_pos_shifted_by2_1_15_port, 
      A_pos_shifted_by2_1_14_port, A_pos_shifted_by2_1_13_port, 
      A_pos_shifted_by2_1_12_port, A_pos_shifted_by2_1_11_port, 
      A_pos_shifted_by2_1_10_port, A_pos_shifted_by2_1_9_port, 
      A_pos_shifted_by2_1_8_port, A_pos_shifted_by2_1_7_port, 
      A_pos_shifted_by2_1_6_port, A_pos_shifted_by2_1_5_port, 
      A_pos_shifted_by2_1_4_port, A_pos_shifted_by2_1_3_port, 
      A_pos_shifted_by2_1_2_port, A_pos_shifted_by2_1_1_port, 
      A_pos_shifted_by2_1_0_port, A_pos_shifted_by2_2_63_port, 
      A_pos_shifted_by2_2_62_port, A_pos_shifted_by2_2_61_port, 
      A_pos_shifted_by2_2_60_port, A_pos_shifted_by2_2_59_port, 
      A_pos_shifted_by2_2_58_port, A_pos_shifted_by2_2_57_port, 
      A_pos_shifted_by2_2_56_port, A_pos_shifted_by2_2_55_port, 
      A_pos_shifted_by2_2_54_port, A_pos_shifted_by2_2_53_port, 
      A_pos_shifted_by2_2_52_port, A_pos_shifted_by2_2_51_port, 
      A_pos_shifted_by2_2_50_port, A_pos_shifted_by2_2_49_port, 
      A_pos_shifted_by2_2_48_port, A_pos_shifted_by2_2_47_port, 
      A_pos_shifted_by2_2_46_port, A_pos_shifted_by2_2_45_port, 
      A_pos_shifted_by2_2_44_port, A_pos_shifted_by2_2_43_port, 
      A_pos_shifted_by2_2_42_port, A_pos_shifted_by2_2_41_port, 
      A_pos_shifted_by2_2_40_port, A_pos_shifted_by2_2_39_port, 
      A_pos_shifted_by2_2_38_port, A_pos_shifted_by2_2_37_port, 
      A_pos_shifted_by2_2_36_port, A_pos_shifted_by2_2_35_port, 
      A_pos_shifted_by2_2_34_port, A_pos_shifted_by2_2_33_port, 
      A_pos_shifted_by2_2_32_port, A_pos_shifted_by2_2_31_port, 
      A_pos_shifted_by2_2_30_port, A_pos_shifted_by2_2_29_port, 
      A_pos_shifted_by2_2_28_port, A_pos_shifted_by2_2_27_port, 
      A_pos_shifted_by2_2_26_port, A_pos_shifted_by2_2_25_port, 
      A_pos_shifted_by2_2_24_port, A_pos_shifted_by2_2_23_port, 
      A_pos_shifted_by2_2_22_port, A_pos_shifted_by2_2_21_port, 
      A_pos_shifted_by2_2_20_port, A_pos_shifted_by2_2_19_port, 
      A_pos_shifted_by2_2_18_port, A_pos_shifted_by2_2_17_port, 
      A_pos_shifted_by2_2_16_port, A_pos_shifted_by2_2_15_port, 
      A_pos_shifted_by2_2_14_port, A_pos_shifted_by2_2_13_port, 
      A_pos_shifted_by2_2_12_port, A_pos_shifted_by2_2_11_port, 
      A_pos_shifted_by2_2_10_port, A_pos_shifted_by2_2_9_port, 
      A_pos_shifted_by2_2_8_port, A_pos_shifted_by2_2_7_port, 
      A_pos_shifted_by2_2_6_port, A_pos_shifted_by2_2_5_port, 
      A_pos_shifted_by2_2_4_port, A_pos_shifted_by2_2_3_port, 
      A_pos_shifted_by2_2_2_port, A_pos_shifted_by2_2_1_port, 
      A_pos_shifted_by2_2_0_port, A_pos_shifted_by2_3_63_port, 
      A_pos_shifted_by2_3_62_port, A_pos_shifted_by2_3_61_port, 
      A_pos_shifted_by2_3_60_port, A_pos_shifted_by2_3_59_port, 
      A_pos_shifted_by2_3_58_port, A_pos_shifted_by2_3_57_port, 
      A_pos_shifted_by2_3_56_port, A_pos_shifted_by2_3_55_port, 
      A_pos_shifted_by2_3_54_port, A_pos_shifted_by2_3_53_port, 
      A_pos_shifted_by2_3_52_port, A_pos_shifted_by2_3_51_port, 
      A_pos_shifted_by2_3_50_port, A_pos_shifted_by2_3_49_port, 
      A_pos_shifted_by2_3_48_port, A_pos_shifted_by2_3_47_port, 
      A_pos_shifted_by2_3_46_port, A_pos_shifted_by2_3_45_port, 
      A_pos_shifted_by2_3_44_port, A_pos_shifted_by2_3_43_port, 
      A_pos_shifted_by2_3_42_port, A_pos_shifted_by2_3_41_port, 
      A_pos_shifted_by2_3_40_port, A_pos_shifted_by2_3_39_port, 
      A_pos_shifted_by2_3_38_port, A_pos_shifted_by2_3_37_port, 
      A_pos_shifted_by2_3_36_port, A_pos_shifted_by2_3_35_port, 
      A_pos_shifted_by2_3_34_port, A_pos_shifted_by2_3_33_port, 
      A_pos_shifted_by2_3_32_port, A_pos_shifted_by2_3_31_port, 
      A_pos_shifted_by2_3_30_port, A_pos_shifted_by2_3_29_port, 
      A_pos_shifted_by2_3_28_port, A_pos_shifted_by2_3_27_port, 
      A_pos_shifted_by2_3_26_port, A_pos_shifted_by2_3_25_port, 
      A_pos_shifted_by2_3_24_port, A_pos_shifted_by2_3_23_port, 
      A_pos_shifted_by2_3_22_port, A_pos_shifted_by2_3_21_port, 
      A_pos_shifted_by2_3_20_port, A_pos_shifted_by2_3_19_port, 
      A_pos_shifted_by2_3_18_port, A_pos_shifted_by2_3_17_port, 
      A_pos_shifted_by2_3_16_port, A_pos_shifted_by2_3_15_port, 
      A_pos_shifted_by2_3_14_port, A_pos_shifted_by2_3_13_port, 
      A_pos_shifted_by2_3_12_port, A_pos_shifted_by2_3_11_port, 
      A_pos_shifted_by2_3_10_port, A_pos_shifted_by2_3_9_port, 
      A_pos_shifted_by2_3_8_port, A_pos_shifted_by2_3_7_port, 
      A_pos_shifted_by2_3_6_port, A_pos_shifted_by2_3_5_port, 
      A_pos_shifted_by2_3_4_port, A_pos_shifted_by2_3_3_port, 
      A_pos_shifted_by2_3_2_port, A_pos_shifted_by2_3_1_port, 
      A_pos_shifted_by2_3_0_port, A_pos_shifted_by2_4_63_port, 
      A_pos_shifted_by2_4_62_port, A_pos_shifted_by2_4_61_port, 
      A_pos_shifted_by2_4_60_port, A_pos_shifted_by2_4_59_port, 
      A_pos_shifted_by2_4_58_port, A_pos_shifted_by2_4_57_port, 
      A_pos_shifted_by2_4_56_port, A_pos_shifted_by2_4_55_port, 
      A_pos_shifted_by2_4_54_port, A_pos_shifted_by2_4_53_port, 
      A_pos_shifted_by2_4_52_port, A_pos_shifted_by2_4_51_port, 
      A_pos_shifted_by2_4_50_port, A_pos_shifted_by2_4_49_port, 
      A_pos_shifted_by2_4_48_port, A_pos_shifted_by2_4_47_port, 
      A_pos_shifted_by2_4_46_port, A_pos_shifted_by2_4_45_port, 
      A_pos_shifted_by2_4_44_port, A_pos_shifted_by2_4_43_port, 
      A_pos_shifted_by2_4_42_port, A_pos_shifted_by2_4_41_port, 
      A_pos_shifted_by2_4_40_port, A_pos_shifted_by2_4_39_port, 
      A_pos_shifted_by2_4_38_port, A_pos_shifted_by2_4_37_port, 
      A_pos_shifted_by2_4_36_port, A_pos_shifted_by2_4_35_port, 
      A_pos_shifted_by2_4_34_port, A_pos_shifted_by2_4_33_port, 
      A_pos_shifted_by2_4_32_port, A_pos_shifted_by2_4_31_port, 
      A_pos_shifted_by2_4_30_port, A_pos_shifted_by2_4_29_port, 
      A_pos_shifted_by2_4_28_port, A_pos_shifted_by2_4_27_port, 
      A_pos_shifted_by2_4_26_port, A_pos_shifted_by2_4_25_port, 
      A_pos_shifted_by2_4_24_port, A_pos_shifted_by2_4_23_port, 
      A_pos_shifted_by2_4_22_port, A_pos_shifted_by2_4_21_port, 
      A_pos_shifted_by2_4_20_port, A_pos_shifted_by2_4_19_port, 
      A_pos_shifted_by2_4_18_port, A_pos_shifted_by2_4_17_port, 
      A_pos_shifted_by2_4_16_port, A_pos_shifted_by2_4_15_port, 
      A_pos_shifted_by2_4_14_port, A_pos_shifted_by2_4_13_port, 
      A_pos_shifted_by2_4_12_port, A_pos_shifted_by2_4_11_port, 
      A_pos_shifted_by2_4_10_port, A_pos_shifted_by2_4_9_port, 
      A_pos_shifted_by2_4_8_port, A_pos_shifted_by2_4_7_port, 
      A_pos_shifted_by2_4_6_port, A_pos_shifted_by2_4_5_port, 
      A_pos_shifted_by2_4_4_port, A_pos_shifted_by2_4_3_port, 
      A_pos_shifted_by2_4_2_port, A_pos_shifted_by2_4_1_port, 
      A_pos_shifted_by2_4_0_port, A_pos_shifted_by2_5_63_port, 
      A_pos_shifted_by2_5_62_port, A_pos_shifted_by2_5_61_port, 
      A_pos_shifted_by2_5_60_port, A_pos_shifted_by2_5_59_port, 
      A_pos_shifted_by2_5_58_port, A_pos_shifted_by2_5_57_port, 
      A_pos_shifted_by2_5_56_port, A_pos_shifted_by2_5_55_port, 
      A_pos_shifted_by2_5_54_port, A_pos_shifted_by2_5_53_port, 
      A_pos_shifted_by2_5_52_port, A_pos_shifted_by2_5_51_port, 
      A_pos_shifted_by2_5_50_port, A_pos_shifted_by2_5_49_port, 
      A_pos_shifted_by2_5_48_port, A_pos_shifted_by2_5_47_port, 
      A_pos_shifted_by2_5_46_port, A_pos_shifted_by2_5_45_port, 
      A_pos_shifted_by2_5_44_port, A_pos_shifted_by2_5_43_port, 
      A_pos_shifted_by2_5_42_port, A_pos_shifted_by2_5_41_port, 
      A_pos_shifted_by2_5_40_port, A_pos_shifted_by2_5_39_port, 
      A_pos_shifted_by2_5_38_port, A_pos_shifted_by2_5_37_port, 
      A_pos_shifted_by2_5_36_port, A_pos_shifted_by2_5_35_port, 
      A_pos_shifted_by2_5_34_port, A_pos_shifted_by2_5_33_port, 
      A_pos_shifted_by2_5_32_port, A_pos_shifted_by2_5_31_port, 
      A_pos_shifted_by2_5_30_port, A_pos_shifted_by2_5_29_port, 
      A_pos_shifted_by2_5_28_port, A_pos_shifted_by2_5_27_port, 
      A_pos_shifted_by2_5_26_port, A_pos_shifted_by2_5_25_port, 
      A_pos_shifted_by2_5_24_port, A_pos_shifted_by2_5_23_port, 
      A_pos_shifted_by2_5_22_port, A_pos_shifted_by2_5_21_port, 
      A_pos_shifted_by2_5_20_port, A_pos_shifted_by2_5_19_port, 
      A_pos_shifted_by2_5_18_port, A_pos_shifted_by2_5_17_port, 
      A_pos_shifted_by2_5_16_port, A_pos_shifted_by2_5_15_port, 
      A_pos_shifted_by2_5_14_port, A_pos_shifted_by2_5_13_port, 
      A_pos_shifted_by2_5_12_port, A_pos_shifted_by2_5_11_port, 
      A_pos_shifted_by2_5_10_port, A_pos_shifted_by2_5_9_port, 
      A_pos_shifted_by2_5_8_port, A_pos_shifted_by2_5_7_port, 
      A_pos_shifted_by2_5_6_port, A_pos_shifted_by2_5_5_port, 
      A_pos_shifted_by2_5_4_port, A_pos_shifted_by2_5_3_port, 
      A_pos_shifted_by2_5_2_port, A_pos_shifted_by2_5_1_port, 
      A_pos_shifted_by2_5_0_port, A_pos_shifted_by2_6_63_port, 
      A_pos_shifted_by2_6_62_port, A_pos_shifted_by2_6_61_port, 
      A_pos_shifted_by2_6_60_port, A_pos_shifted_by2_6_59_port, 
      A_pos_shifted_by2_6_58_port, A_pos_shifted_by2_6_57_port, 
      A_pos_shifted_by2_6_56_port, A_pos_shifted_by2_6_55_port, 
      A_pos_shifted_by2_6_54_port, A_pos_shifted_by2_6_53_port, 
      A_pos_shifted_by2_6_52_port, A_pos_shifted_by2_6_51_port, 
      A_pos_shifted_by2_6_50_port, A_pos_shifted_by2_6_49_port, 
      A_pos_shifted_by2_6_48_port, A_pos_shifted_by2_6_47_port, 
      A_pos_shifted_by2_6_46_port, A_pos_shifted_by2_6_45_port, 
      A_pos_shifted_by2_6_44_port, A_pos_shifted_by2_6_43_port, 
      A_pos_shifted_by2_6_42_port, A_pos_shifted_by2_6_41_port, 
      A_pos_shifted_by2_6_40_port, A_pos_shifted_by2_6_39_port, 
      A_pos_shifted_by2_6_38_port, A_pos_shifted_by2_6_37_port, 
      A_pos_shifted_by2_6_36_port, A_pos_shifted_by2_6_35_port, 
      A_pos_shifted_by2_6_34_port, A_pos_shifted_by2_6_33_port, 
      A_pos_shifted_by2_6_32_port, A_pos_shifted_by2_6_31_port, 
      A_pos_shifted_by2_6_30_port, A_pos_shifted_by2_6_29_port, 
      A_pos_shifted_by2_6_28_port, A_pos_shifted_by2_6_27_port, 
      A_pos_shifted_by2_6_26_port, A_pos_shifted_by2_6_25_port, 
      A_pos_shifted_by2_6_24_port, A_pos_shifted_by2_6_23_port, 
      A_pos_shifted_by2_6_22_port, A_pos_shifted_by2_6_21_port, 
      A_pos_shifted_by2_6_20_port, A_pos_shifted_by2_6_19_port, 
      A_pos_shifted_by2_6_18_port, A_pos_shifted_by2_6_17_port, 
      A_pos_shifted_by2_6_16_port, A_pos_shifted_by2_6_15_port, 
      A_pos_shifted_by2_6_14_port, A_pos_shifted_by2_6_13_port, 
      A_pos_shifted_by2_6_12_port, A_pos_shifted_by2_6_11_port, 
      A_pos_shifted_by2_6_10_port, A_pos_shifted_by2_6_9_port, 
      A_pos_shifted_by2_6_8_port, A_pos_shifted_by2_6_7_port, 
      A_pos_shifted_by2_6_6_port, A_pos_shifted_by2_6_5_port, 
      A_pos_shifted_by2_6_4_port, A_pos_shifted_by2_6_3_port, 
      A_pos_shifted_by2_6_2_port, A_pos_shifted_by2_6_1_port, 
      A_pos_shifted_by2_6_0_port, A_pos_shifted_by2_7_63_port, 
      A_pos_shifted_by2_7_62_port, A_pos_shifted_by2_7_61_port, 
      A_pos_shifted_by2_7_60_port, A_pos_shifted_by2_7_59_port, 
      A_pos_shifted_by2_7_58_port, A_pos_shifted_by2_7_57_port, 
      A_pos_shifted_by2_7_56_port, A_pos_shifted_by2_7_55_port, 
      A_pos_shifted_by2_7_54_port, A_pos_shifted_by2_7_53_port, 
      A_pos_shifted_by2_7_52_port, A_pos_shifted_by2_7_51_port, 
      A_pos_shifted_by2_7_50_port, A_pos_shifted_by2_7_49_port, 
      A_pos_shifted_by2_7_48_port, A_pos_shifted_by2_7_47_port, 
      A_pos_shifted_by2_7_46_port, A_pos_shifted_by2_7_45_port, 
      A_pos_shifted_by2_7_44_port, A_pos_shifted_by2_7_43_port, 
      A_pos_shifted_by2_7_42_port, A_pos_shifted_by2_7_41_port, 
      A_pos_shifted_by2_7_40_port, A_pos_shifted_by2_7_39_port, 
      A_pos_shifted_by2_7_38_port, A_pos_shifted_by2_7_37_port, 
      A_pos_shifted_by2_7_36_port, A_pos_shifted_by2_7_35_port, 
      A_pos_shifted_by2_7_34_port, A_pos_shifted_by2_7_33_port, 
      A_pos_shifted_by2_7_32_port, A_pos_shifted_by2_7_31_port, 
      A_pos_shifted_by2_7_30_port, A_pos_shifted_by2_7_29_port, 
      A_pos_shifted_by2_7_28_port, A_pos_shifted_by2_7_27_port, 
      A_pos_shifted_by2_7_26_port, A_pos_shifted_by2_7_25_port, 
      A_pos_shifted_by2_7_24_port, A_pos_shifted_by2_7_23_port, 
      A_pos_shifted_by2_7_22_port, A_pos_shifted_by2_7_21_port, 
      A_pos_shifted_by2_7_20_port, A_pos_shifted_by2_7_19_port, 
      A_pos_shifted_by2_7_18_port, A_pos_shifted_by2_7_17_port, 
      A_pos_shifted_by2_7_16_port, A_pos_shifted_by2_7_15_port, 
      A_pos_shifted_by2_7_14_port, A_pos_shifted_by2_7_13_port, 
      A_pos_shifted_by2_7_12_port, A_pos_shifted_by2_7_11_port, 
      A_pos_shifted_by2_7_10_port, A_pos_shifted_by2_7_9_port, 
      A_pos_shifted_by2_7_8_port, A_pos_shifted_by2_7_7_port, 
      A_pos_shifted_by2_7_6_port, A_pos_shifted_by2_7_5_port, 
      A_pos_shifted_by2_7_4_port, A_pos_shifted_by2_7_3_port, 
      A_pos_shifted_by2_7_2_port, A_pos_shifted_by2_7_1_port, 
      A_pos_shifted_by2_7_0_port, A_pos_shifted_by1_8_63_port, 
      A_pos_shifted_by1_8_62_port, A_pos_shifted_by1_8_61_port, 
      A_pos_shifted_by1_8_60_port, A_pos_shifted_by1_8_59_port, 
      A_pos_shifted_by1_8_58_port, A_pos_shifted_by1_8_57_port, 
      A_pos_shifted_by1_8_56_port, A_pos_shifted_by1_8_55_port, 
      A_pos_shifted_by1_8_54_port, A_pos_shifted_by1_8_53_port, 
      A_pos_shifted_by1_8_52_port, A_pos_shifted_by1_8_51_port, 
      A_pos_shifted_by1_8_50_port, A_pos_shifted_by1_8_49_port, 
      A_pos_shifted_by1_8_48_port, A_pos_shifted_by1_8_47_port, 
      A_pos_shifted_by1_8_46_port, A_pos_shifted_by1_8_45_port, 
      A_pos_shifted_by1_8_44_port, A_pos_shifted_by1_8_43_port, 
      A_pos_shifted_by1_8_42_port, A_pos_shifted_by1_8_41_port, 
      A_pos_shifted_by1_8_40_port, A_pos_shifted_by1_8_39_port, 
      A_pos_shifted_by1_8_38_port, A_pos_shifted_by1_8_37_port, 
      A_pos_shifted_by1_8_36_port, A_pos_shifted_by1_8_35_port, 
      A_pos_shifted_by1_8_34_port, A_pos_shifted_by1_8_33_port, 
      A_pos_shifted_by1_8_32_port, A_pos_shifted_by1_8_31_port, 
      A_pos_shifted_by1_8_30_port, A_pos_shifted_by1_8_29_port, 
      A_pos_shifted_by1_8_28_port, A_pos_shifted_by1_8_27_port, 
      A_pos_shifted_by1_8_26_port, A_pos_shifted_by1_8_25_port, 
      A_pos_shifted_by1_8_24_port, A_pos_shifted_by1_8_23_port, 
      A_pos_shifted_by1_8_22_port, A_pos_shifted_by1_8_21_port, 
      A_pos_shifted_by1_8_20_port, A_pos_shifted_by1_8_19_port, 
      A_pos_shifted_by1_8_18_port, A_pos_shifted_by1_8_17_port, 
      A_pos_shifted_by1_8_16_port, A_pos_shifted_by1_8_15_port, 
      A_pos_shifted_by1_8_14_port, A_pos_shifted_by1_8_13_port, 
      A_pos_shifted_by1_8_12_port, A_pos_shifted_by1_8_11_port, 
      A_pos_shifted_by1_8_10_port, A_pos_shifted_by1_8_9_port, 
      A_pos_shifted_by1_8_8_port, A_pos_shifted_by1_8_7_port, 
      A_pos_shifted_by1_8_6_port, A_pos_shifted_by1_8_5_port, 
      A_pos_shifted_by1_8_4_port, A_pos_shifted_by1_8_3_port, 
      A_pos_shifted_by1_8_2_port, A_pos_shifted_by1_8_1_port, 
      A_pos_shifted_by1_8_0_port, A_pos_shifted_by1_9_63_port, 
      A_pos_shifted_by1_9_62_port, A_pos_shifted_by1_9_61_port, 
      A_pos_shifted_by1_9_60_port, A_pos_shifted_by1_9_59_port, 
      A_pos_shifted_by1_9_58_port, A_pos_shifted_by1_9_57_port, 
      A_pos_shifted_by1_9_56_port, A_pos_shifted_by1_9_55_port, 
      A_pos_shifted_by1_9_54_port, A_pos_shifted_by1_9_53_port, 
      A_pos_shifted_by1_9_52_port, A_pos_shifted_by1_9_51_port, 
      A_pos_shifted_by1_9_50_port, A_pos_shifted_by1_9_49_port, 
      A_pos_shifted_by1_9_48_port, A_pos_shifted_by1_9_47_port, 
      A_pos_shifted_by1_9_46_port, A_pos_shifted_by1_9_45_port, 
      A_pos_shifted_by1_9_44_port, A_pos_shifted_by1_9_43_port, 
      A_pos_shifted_by1_9_42_port, A_pos_shifted_by1_9_41_port, 
      A_pos_shifted_by1_9_40_port, A_pos_shifted_by1_9_39_port, 
      A_pos_shifted_by1_9_38_port, A_pos_shifted_by1_9_37_port, 
      A_pos_shifted_by1_9_36_port, A_pos_shifted_by1_9_35_port, 
      A_pos_shifted_by1_9_34_port, A_pos_shifted_by1_9_33_port, 
      A_pos_shifted_by1_9_32_port, A_pos_shifted_by1_9_31_port, 
      A_pos_shifted_by1_9_30_port, A_pos_shifted_by1_9_29_port, 
      A_pos_shifted_by1_9_28_port, A_pos_shifted_by1_9_27_port, 
      A_pos_shifted_by1_9_26_port, A_pos_shifted_by1_9_25_port, 
      A_pos_shifted_by1_9_24_port, A_pos_shifted_by1_9_23_port, 
      A_pos_shifted_by1_9_22_port, A_pos_shifted_by1_9_21_port, 
      A_pos_shifted_by1_9_20_port, A_pos_shifted_by1_9_19_port, 
      A_pos_shifted_by1_9_18_port, A_pos_shifted_by1_9_17_port, 
      A_pos_shifted_by1_9_16_port, A_pos_shifted_by1_9_15_port, 
      A_pos_shifted_by1_9_14_port, A_pos_shifted_by1_9_13_port, 
      A_pos_shifted_by1_9_12_port, A_pos_shifted_by1_9_11_port, 
      A_pos_shifted_by1_9_10_port, A_pos_shifted_by1_9_9_port, 
      A_pos_shifted_by1_9_8_port, A_pos_shifted_by1_9_7_port, 
      A_pos_shifted_by1_9_6_port, A_pos_shifted_by1_9_5_port, 
      A_pos_shifted_by1_9_4_port, A_pos_shifted_by1_9_3_port, 
      A_pos_shifted_by1_9_2_port, A_pos_shifted_by1_9_1_port, 
      A_pos_shifted_by1_9_0_port, A_pos_shifted_by1_10_63_port, 
      A_pos_shifted_by1_10_62_port, A_pos_shifted_by1_10_61_port, 
      A_pos_shifted_by1_10_60_port, A_pos_shifted_by1_10_59_port, 
      A_pos_shifted_by1_10_58_port, A_pos_shifted_by1_10_57_port, 
      A_pos_shifted_by1_10_56_port, A_pos_shifted_by1_10_55_port, 
      A_pos_shifted_by1_10_54_port, A_pos_shifted_by1_10_53_port, 
      A_pos_shifted_by1_10_52_port, A_pos_shifted_by1_10_51_port, 
      A_pos_shifted_by1_10_50_port, A_pos_shifted_by1_10_49_port, 
      A_pos_shifted_by1_10_48_port, A_pos_shifted_by1_10_47_port, 
      A_pos_shifted_by1_10_46_port, A_pos_shifted_by1_10_45_port, 
      A_pos_shifted_by1_10_44_port, A_pos_shifted_by1_10_43_port, 
      A_pos_shifted_by1_10_42_port, A_pos_shifted_by1_10_41_port, 
      A_pos_shifted_by1_10_40_port, A_pos_shifted_by1_10_39_port, 
      A_pos_shifted_by1_10_38_port, A_pos_shifted_by1_10_37_port, 
      A_pos_shifted_by1_10_36_port, A_pos_shifted_by1_10_35_port, 
      A_pos_shifted_by1_10_34_port, A_pos_shifted_by1_10_33_port, 
      A_pos_shifted_by1_10_32_port, A_pos_shifted_by1_10_31_port, 
      A_pos_shifted_by1_10_30_port, A_pos_shifted_by1_10_29_port, 
      A_pos_shifted_by1_10_28_port, A_pos_shifted_by1_10_27_port, 
      A_pos_shifted_by1_10_26_port, A_pos_shifted_by1_10_25_port, 
      A_pos_shifted_by1_10_24_port, A_pos_shifted_by1_10_23_port, 
      A_pos_shifted_by1_10_22_port, A_pos_shifted_by1_10_21_port, 
      A_pos_shifted_by1_10_20_port, A_pos_shifted_by1_10_19_port, 
      A_pos_shifted_by1_10_18_port, A_pos_shifted_by1_10_17_port, 
      A_pos_shifted_by1_10_16_port, A_pos_shifted_by1_10_15_port, 
      A_pos_shifted_by1_10_14_port, A_pos_shifted_by1_10_13_port, 
      A_pos_shifted_by1_10_12_port, A_pos_shifted_by1_10_11_port, 
      A_pos_shifted_by1_10_10_port, A_pos_shifted_by1_10_9_port, 
      A_pos_shifted_by1_10_8_port, A_pos_shifted_by1_10_7_port, 
      A_pos_shifted_by1_10_6_port, A_pos_shifted_by1_10_5_port, 
      A_pos_shifted_by1_10_4_port, A_pos_shifted_by1_10_3_port, 
      A_pos_shifted_by1_10_2_port, A_pos_shifted_by1_10_1_port, 
      A_pos_shifted_by1_10_0_port, A_pos_shifted_by1_11_63_port, 
      A_pos_shifted_by1_11_62_port, A_pos_shifted_by1_11_61_port, 
      A_pos_shifted_by1_11_60_port, A_pos_shifted_by1_11_59_port, 
      A_pos_shifted_by1_11_58_port, A_pos_shifted_by1_11_57_port, 
      A_pos_shifted_by1_11_56_port, A_pos_shifted_by1_11_55_port, 
      A_pos_shifted_by1_11_54_port, A_pos_shifted_by1_11_53_port, 
      A_pos_shifted_by1_11_52_port, A_pos_shifted_by1_11_51_port, 
      A_pos_shifted_by1_11_50_port, A_pos_shifted_by1_11_49_port, 
      A_pos_shifted_by1_11_48_port, A_pos_shifted_by1_11_47_port, 
      A_pos_shifted_by1_11_46_port, A_pos_shifted_by1_11_45_port, 
      A_pos_shifted_by1_11_44_port, A_pos_shifted_by1_11_43_port, 
      A_pos_shifted_by1_11_42_port, A_pos_shifted_by1_11_41_port, 
      A_pos_shifted_by1_11_40_port, A_pos_shifted_by1_11_39_port, 
      A_pos_shifted_by1_11_38_port, A_pos_shifted_by1_11_37_port, 
      A_pos_shifted_by1_11_36_port, A_pos_shifted_by1_11_35_port, 
      A_pos_shifted_by1_11_34_port, A_pos_shifted_by1_11_33_port, 
      A_pos_shifted_by1_11_32_port, A_pos_shifted_by1_11_31_port, 
      A_pos_shifted_by1_11_30_port, A_pos_shifted_by1_11_29_port, 
      A_pos_shifted_by1_11_28_port, A_pos_shifted_by1_11_27_port, 
      A_pos_shifted_by1_11_26_port, A_pos_shifted_by1_11_25_port, 
      A_pos_shifted_by1_11_24_port, A_pos_shifted_by1_11_23_port, 
      A_pos_shifted_by1_11_22_port, A_pos_shifted_by1_11_21_port, 
      A_pos_shifted_by1_11_20_port, A_pos_shifted_by1_11_19_port, 
      A_pos_shifted_by1_11_18_port, A_pos_shifted_by1_11_17_port, 
      A_pos_shifted_by1_11_16_port, A_pos_shifted_by1_11_15_port, 
      A_pos_shifted_by1_11_14_port, A_pos_shifted_by1_11_13_port, 
      A_pos_shifted_by1_11_12_port, A_pos_shifted_by1_11_11_port, 
      A_pos_shifted_by1_11_10_port, A_pos_shifted_by1_11_9_port, 
      A_pos_shifted_by1_11_8_port, A_pos_shifted_by1_11_7_port, 
      A_pos_shifted_by1_11_6_port, A_pos_shifted_by1_11_5_port, 
      A_pos_shifted_by1_11_4_port, A_pos_shifted_by1_11_3_port, 
      A_pos_shifted_by1_11_2_port, A_pos_shifted_by1_11_1_port, 
      A_pos_shifted_by1_11_0_port, A_pos_shifted_by1_12_63_port, 
      A_pos_shifted_by1_12_62_port, A_pos_shifted_by1_12_61_port, 
      A_pos_shifted_by1_12_60_port, A_pos_shifted_by1_12_59_port, 
      A_pos_shifted_by1_12_58_port, A_pos_shifted_by1_12_57_port, 
      A_pos_shifted_by1_12_56_port, A_pos_shifted_by1_12_55_port, 
      A_pos_shifted_by1_12_54_port, A_pos_shifted_by1_12_53_port, 
      A_pos_shifted_by1_12_52_port, A_pos_shifted_by1_12_51_port, 
      A_pos_shifted_by1_12_50_port, A_pos_shifted_by1_12_49_port, 
      A_pos_shifted_by1_12_48_port, A_pos_shifted_by1_12_47_port, 
      A_pos_shifted_by1_12_46_port, A_pos_shifted_by1_12_45_port, 
      A_pos_shifted_by1_12_44_port, A_pos_shifted_by1_12_43_port, 
      A_pos_shifted_by1_12_42_port, A_pos_shifted_by1_12_41_port, 
      A_pos_shifted_by1_12_40_port, A_pos_shifted_by1_12_39_port, 
      A_pos_shifted_by1_12_38_port, A_pos_shifted_by1_12_37_port, 
      A_pos_shifted_by1_12_36_port, A_pos_shifted_by1_12_35_port, 
      A_pos_shifted_by1_12_34_port, A_pos_shifted_by1_12_33_port, 
      A_pos_shifted_by1_12_32_port, A_pos_shifted_by1_12_31_port, 
      A_pos_shifted_by1_12_30_port, A_pos_shifted_by1_12_29_port, 
      A_pos_shifted_by1_12_28_port, A_pos_shifted_by1_12_27_port, 
      A_pos_shifted_by1_12_26_port, A_pos_shifted_by1_12_25_port, 
      A_pos_shifted_by1_12_24_port, A_pos_shifted_by1_12_23_port, 
      A_pos_shifted_by1_12_22_port, A_pos_shifted_by1_12_21_port, 
      A_pos_shifted_by1_12_20_port, A_pos_shifted_by1_12_19_port, 
      A_pos_shifted_by1_12_18_port, A_pos_shifted_by1_12_17_port, 
      A_pos_shifted_by1_12_16_port, A_pos_shifted_by1_12_15_port, 
      A_pos_shifted_by1_12_14_port, A_pos_shifted_by1_12_13_port, 
      A_pos_shifted_by1_12_12_port, A_pos_shifted_by1_12_11_port, 
      A_pos_shifted_by1_12_10_port, A_pos_shifted_by1_12_9_port, 
      A_pos_shifted_by1_12_8_port, A_pos_shifted_by1_12_7_port, 
      A_pos_shifted_by1_12_6_port, A_pos_shifted_by1_12_5_port, 
      A_pos_shifted_by1_12_4_port, A_pos_shifted_by1_12_3_port, 
      A_pos_shifted_by1_12_2_port, A_pos_shifted_by1_12_1_port, 
      A_pos_shifted_by1_12_0_port, A_pos_shifted_by1_13_63_port, 
      A_pos_shifted_by1_13_62_port, A_pos_shifted_by1_13_61_port, 
      A_pos_shifted_by1_13_60_port, A_pos_shifted_by1_13_59_port, 
      A_pos_shifted_by1_13_58_port, A_pos_shifted_by1_13_57_port, 
      A_pos_shifted_by1_13_56_port, A_pos_shifted_by1_13_55_port, 
      A_pos_shifted_by1_13_54_port, A_pos_shifted_by1_13_53_port, 
      A_pos_shifted_by1_13_52_port, A_pos_shifted_by1_13_51_port, 
      A_pos_shifted_by1_13_50_port, A_pos_shifted_by1_13_49_port, 
      A_pos_shifted_by1_13_48_port, A_pos_shifted_by1_13_47_port, 
      A_pos_shifted_by1_13_46_port, A_pos_shifted_by1_13_45_port, 
      A_pos_shifted_by1_13_44_port, A_pos_shifted_by1_13_43_port, 
      A_pos_shifted_by1_13_42_port, A_pos_shifted_by1_13_41_port, 
      A_pos_shifted_by1_13_40_port, A_pos_shifted_by1_13_39_port, 
      A_pos_shifted_by1_13_38_port, A_pos_shifted_by1_13_37_port, 
      A_pos_shifted_by1_13_36_port, A_pos_shifted_by1_13_35_port, 
      A_pos_shifted_by1_13_34_port, A_pos_shifted_by1_13_33_port, 
      A_pos_shifted_by1_13_32_port, A_pos_shifted_by1_13_31_port, 
      A_pos_shifted_by1_13_30_port, A_pos_shifted_by1_13_29_port, 
      A_pos_shifted_by1_13_28_port, A_pos_shifted_by1_13_27_port, 
      A_pos_shifted_by1_13_26_port, A_pos_shifted_by1_13_25_port, 
      A_pos_shifted_by1_13_24_port, A_pos_shifted_by1_13_23_port, 
      A_pos_shifted_by1_13_22_port, A_pos_shifted_by1_13_21_port, 
      A_pos_shifted_by1_13_20_port, A_pos_shifted_by1_13_19_port, 
      A_pos_shifted_by1_13_18_port, A_pos_shifted_by1_13_17_port, 
      A_pos_shifted_by1_13_16_port, A_pos_shifted_by1_13_15_port, 
      A_pos_shifted_by1_13_14_port, A_pos_shifted_by1_13_13_port, 
      A_pos_shifted_by1_13_12_port, A_pos_shifted_by1_13_11_port, 
      A_pos_shifted_by1_13_10_port, A_pos_shifted_by1_13_9_port, 
      A_pos_shifted_by1_13_8_port, A_pos_shifted_by1_13_7_port, 
      A_pos_shifted_by1_13_6_port, A_pos_shifted_by1_13_5_port, 
      A_pos_shifted_by1_13_4_port, A_pos_shifted_by1_13_3_port, 
      A_pos_shifted_by1_13_2_port, A_pos_shifted_by1_13_1_port, 
      A_pos_shifted_by1_13_0_port, A_pos_shifted_by1_14_63_port, 
      A_pos_shifted_by1_14_62_port, A_pos_shifted_by1_14_61_port, 
      A_pos_shifted_by1_14_60_port, A_pos_shifted_by1_14_59_port, 
      A_pos_shifted_by1_14_58_port, A_pos_shifted_by1_14_57_port, 
      A_pos_shifted_by1_14_56_port, A_pos_shifted_by1_14_55_port, 
      A_pos_shifted_by1_14_54_port, A_pos_shifted_by1_14_53_port, 
      A_pos_shifted_by1_14_52_port, A_pos_shifted_by1_14_51_port, 
      A_pos_shifted_by1_14_50_port, A_pos_shifted_by1_14_49_port, 
      A_pos_shifted_by1_14_48_port, A_pos_shifted_by1_14_47_port, 
      A_pos_shifted_by1_14_46_port, A_pos_shifted_by1_14_45_port, 
      A_pos_shifted_by1_14_44_port, A_pos_shifted_by1_14_43_port, 
      A_pos_shifted_by1_14_42_port, A_pos_shifted_by1_14_41_port, 
      A_pos_shifted_by1_14_40_port, A_pos_shifted_by1_14_39_port, 
      A_pos_shifted_by1_14_38_port, A_pos_shifted_by1_14_37_port, 
      A_pos_shifted_by1_14_36_port, A_pos_shifted_by1_14_35_port, 
      A_pos_shifted_by1_14_34_port, A_pos_shifted_by1_14_33_port, 
      A_pos_shifted_by1_14_32_port, A_pos_shifted_by1_14_31_port, 
      A_pos_shifted_by1_14_30_port, A_pos_shifted_by1_14_29_port, 
      A_pos_shifted_by1_14_28_port, A_pos_shifted_by1_14_27_port, 
      A_pos_shifted_by1_14_26_port, A_pos_shifted_by1_14_25_port, 
      A_pos_shifted_by1_14_24_port, A_pos_shifted_by1_14_23_port, 
      A_pos_shifted_by1_14_22_port, A_pos_shifted_by1_14_21_port, 
      A_pos_shifted_by1_14_20_port, A_pos_shifted_by1_14_19_port, 
      A_pos_shifted_by1_14_18_port, A_pos_shifted_by1_14_17_port, 
      A_pos_shifted_by1_14_16_port, A_pos_shifted_by1_14_15_port, 
      A_pos_shifted_by1_14_14_port, A_pos_shifted_by1_14_13_port, 
      A_pos_shifted_by1_14_12_port, A_pos_shifted_by1_14_11_port, 
      A_pos_shifted_by1_14_10_port, A_pos_shifted_by1_14_9_port, 
      A_pos_shifted_by1_14_8_port, A_pos_shifted_by1_14_7_port, 
      A_pos_shifted_by1_14_6_port, A_pos_shifted_by1_14_5_port, 
      A_pos_shifted_by1_14_4_port, A_pos_shifted_by1_14_3_port, 
      A_pos_shifted_by1_14_2_port, A_pos_shifted_by1_14_1_port, 
      A_pos_shifted_by1_14_0_port, A_pos_shifted_by1_15_63_port, 
      A_pos_shifted_by1_15_62_port, A_pos_shifted_by1_15_61_port, 
      A_pos_shifted_by1_15_60_port, A_pos_shifted_by1_15_59_port, 
      A_pos_shifted_by1_15_58_port, A_pos_shifted_by1_15_57_port, 
      A_pos_shifted_by1_15_56_port, A_pos_shifted_by1_15_55_port, 
      A_pos_shifted_by1_15_54_port, A_pos_shifted_by1_15_53_port, 
      A_pos_shifted_by1_15_52_port, A_pos_shifted_by1_15_51_port, 
      A_pos_shifted_by1_15_50_port, A_pos_shifted_by1_15_49_port, 
      A_pos_shifted_by1_15_48_port, A_pos_shifted_by1_15_47_port, 
      A_pos_shifted_by1_15_46_port, A_pos_shifted_by1_15_45_port, 
      A_pos_shifted_by1_15_44_port, A_pos_shifted_by1_15_43_port, 
      A_pos_shifted_by1_15_42_port, A_pos_shifted_by1_15_41_port, 
      A_pos_shifted_by1_15_40_port, A_pos_shifted_by1_15_39_port, 
      A_pos_shifted_by1_15_38_port, A_pos_shifted_by1_15_37_port, 
      A_pos_shifted_by1_15_36_port, A_pos_shifted_by1_15_35_port, 
      A_pos_shifted_by1_15_34_port, A_pos_shifted_by1_15_33_port, 
      A_pos_shifted_by1_15_32_port, A_pos_shifted_by1_15_31_port, 
      A_pos_shifted_by1_15_30_port, A_pos_shifted_by1_15_29_port, 
      A_pos_shifted_by1_15_28_port, A_pos_shifted_by1_15_27_port, 
      A_pos_shifted_by1_15_26_port, A_pos_shifted_by1_15_25_port, 
      A_pos_shifted_by1_15_24_port, A_pos_shifted_by1_15_23_port, 
      A_pos_shifted_by1_15_22_port, A_pos_shifted_by1_15_21_port, 
      A_pos_shifted_by1_15_20_port, A_pos_shifted_by1_15_19_port, 
      A_pos_shifted_by1_15_18_port, A_pos_shifted_by1_15_17_port, 
      A_pos_shifted_by1_15_16_port, A_pos_shifted_by1_15_15_port, 
      A_pos_shifted_by1_15_14_port, A_pos_shifted_by1_15_13_port, 
      A_pos_shifted_by1_15_12_port, A_pos_shifted_by1_15_11_port, 
      A_pos_shifted_by1_15_10_port, A_pos_shifted_by1_15_9_port, 
      A_pos_shifted_by1_15_8_port, A_pos_shifted_by1_15_7_port, 
      A_pos_shifted_by1_15_6_port, A_pos_shifted_by1_15_5_port, 
      A_pos_shifted_by1_15_4_port, A_pos_shifted_by1_15_3_port, 
      A_pos_shifted_by1_15_2_port, A_pos_shifted_by1_15_1_port, 
      A_pos_shifted_by1_15_0_port, A_pos_shifted_by2_8_63_port, 
      A_pos_shifted_by2_8_62_port, A_pos_shifted_by2_8_61_port, 
      A_pos_shifted_by2_8_60_port, A_pos_shifted_by2_8_59_port, 
      A_pos_shifted_by2_8_58_port, A_pos_shifted_by2_8_57_port, 
      A_pos_shifted_by2_8_56_port, A_pos_shifted_by2_8_55_port, 
      A_pos_shifted_by2_8_54_port, A_pos_shifted_by2_8_53_port, 
      A_pos_shifted_by2_8_52_port, A_pos_shifted_by2_8_51_port, 
      A_pos_shifted_by2_8_50_port, A_pos_shifted_by2_8_49_port, 
      A_pos_shifted_by2_8_48_port, A_pos_shifted_by2_8_47_port, 
      A_pos_shifted_by2_8_46_port, A_pos_shifted_by2_8_45_port, 
      A_pos_shifted_by2_8_44_port, A_pos_shifted_by2_8_43_port, 
      A_pos_shifted_by2_8_42_port, A_pos_shifted_by2_8_41_port, 
      A_pos_shifted_by2_8_40_port, A_pos_shifted_by2_8_39_port, 
      A_pos_shifted_by2_8_38_port, A_pos_shifted_by2_8_37_port, 
      A_pos_shifted_by2_8_36_port, A_pos_shifted_by2_8_35_port, 
      A_pos_shifted_by2_8_34_port, A_pos_shifted_by2_8_33_port, 
      A_pos_shifted_by2_8_32_port, A_pos_shifted_by2_8_31_port, 
      A_pos_shifted_by2_8_30_port, A_pos_shifted_by2_8_29_port, 
      A_pos_shifted_by2_8_28_port, A_pos_shifted_by2_8_27_port, 
      A_pos_shifted_by2_8_26_port, A_pos_shifted_by2_8_25_port, 
      A_pos_shifted_by2_8_24_port, A_pos_shifted_by2_8_23_port, 
      A_pos_shifted_by2_8_22_port, A_pos_shifted_by2_8_21_port, 
      A_pos_shifted_by2_8_20_port, A_pos_shifted_by2_8_19_port, 
      A_pos_shifted_by2_8_18_port, A_pos_shifted_by2_8_17_port, 
      A_pos_shifted_by2_8_16_port, A_pos_shifted_by2_8_15_port, 
      A_pos_shifted_by2_8_14_port, A_pos_shifted_by2_8_13_port, 
      A_pos_shifted_by2_8_12_port, A_pos_shifted_by2_8_11_port, 
      A_pos_shifted_by2_8_10_port, A_pos_shifted_by2_8_9_port, 
      A_pos_shifted_by2_8_8_port, A_pos_shifted_by2_8_7_port, 
      A_pos_shifted_by2_8_6_port, A_pos_shifted_by2_8_5_port, 
      A_pos_shifted_by2_8_4_port, A_pos_shifted_by2_8_3_port, 
      A_pos_shifted_by2_8_2_port, A_pos_shifted_by2_8_1_port, 
      A_pos_shifted_by2_8_0_port, A_pos_shifted_by2_9_63_port, 
      A_pos_shifted_by2_9_62_port, A_pos_shifted_by2_9_61_port, 
      A_pos_shifted_by2_9_60_port, A_pos_shifted_by2_9_59_port, 
      A_pos_shifted_by2_9_58_port, A_pos_shifted_by2_9_57_port, 
      A_pos_shifted_by2_9_56_port, A_pos_shifted_by2_9_55_port, 
      A_pos_shifted_by2_9_54_port, A_pos_shifted_by2_9_53_port, 
      A_pos_shifted_by2_9_52_port, A_pos_shifted_by2_9_51_port, 
      A_pos_shifted_by2_9_50_port, A_pos_shifted_by2_9_49_port, 
      A_pos_shifted_by2_9_48_port, A_pos_shifted_by2_9_47_port, 
      A_pos_shifted_by2_9_46_port, A_pos_shifted_by2_9_45_port, 
      A_pos_shifted_by2_9_44_port, A_pos_shifted_by2_9_43_port, 
      A_pos_shifted_by2_9_42_port, A_pos_shifted_by2_9_41_port, 
      A_pos_shifted_by2_9_40_port, A_pos_shifted_by2_9_39_port, 
      A_pos_shifted_by2_9_38_port, A_pos_shifted_by2_9_37_port, 
      A_pos_shifted_by2_9_36_port, A_pos_shifted_by2_9_35_port, 
      A_pos_shifted_by2_9_34_port, A_pos_shifted_by2_9_33_port, 
      A_pos_shifted_by2_9_32_port, A_pos_shifted_by2_9_31_port, 
      A_pos_shifted_by2_9_30_port, A_pos_shifted_by2_9_29_port, 
      A_pos_shifted_by2_9_28_port, A_pos_shifted_by2_9_27_port, 
      A_pos_shifted_by2_9_26_port, A_pos_shifted_by2_9_25_port, 
      A_pos_shifted_by2_9_24_port, A_pos_shifted_by2_9_23_port, 
      A_pos_shifted_by2_9_22_port, A_pos_shifted_by2_9_21_port, 
      A_pos_shifted_by2_9_20_port, A_pos_shifted_by2_9_19_port, 
      A_pos_shifted_by2_9_18_port, A_pos_shifted_by2_9_17_port, 
      A_pos_shifted_by2_9_16_port, A_pos_shifted_by2_9_15_port, 
      A_pos_shifted_by2_9_14_port, A_pos_shifted_by2_9_13_port, 
      A_pos_shifted_by2_9_12_port, A_pos_shifted_by2_9_11_port, 
      A_pos_shifted_by2_9_10_port, A_pos_shifted_by2_9_9_port, 
      A_pos_shifted_by2_9_8_port, A_pos_shifted_by2_9_7_port, 
      A_pos_shifted_by2_9_6_port, A_pos_shifted_by2_9_5_port, 
      A_pos_shifted_by2_9_4_port, A_pos_shifted_by2_9_3_port, 
      A_pos_shifted_by2_9_2_port, A_pos_shifted_by2_9_1_port, 
      A_pos_shifted_by2_9_0_port, A_pos_shifted_by2_10_63_port, 
      A_pos_shifted_by2_10_62_port, A_pos_shifted_by2_10_61_port, 
      A_pos_shifted_by2_10_60_port, A_pos_shifted_by2_10_59_port, 
      A_pos_shifted_by2_10_58_port, A_pos_shifted_by2_10_57_port, 
      A_pos_shifted_by2_10_56_port, A_pos_shifted_by2_10_55_port, 
      A_pos_shifted_by2_10_54_port, A_pos_shifted_by2_10_53_port, 
      A_pos_shifted_by2_10_52_port, A_pos_shifted_by2_10_51_port, 
      A_pos_shifted_by2_10_50_port, A_pos_shifted_by2_10_49_port, 
      A_pos_shifted_by2_10_48_port, A_pos_shifted_by2_10_47_port, 
      A_pos_shifted_by2_10_46_port, A_pos_shifted_by2_10_45_port, 
      A_pos_shifted_by2_10_44_port, A_pos_shifted_by2_10_43_port, 
      A_pos_shifted_by2_10_42_port, A_pos_shifted_by2_10_41_port, 
      A_pos_shifted_by2_10_40_port, A_pos_shifted_by2_10_39_port, 
      A_pos_shifted_by2_10_38_port, A_pos_shifted_by2_10_37_port, 
      A_pos_shifted_by2_10_36_port, A_pos_shifted_by2_10_35_port, 
      A_pos_shifted_by2_10_34_port, A_pos_shifted_by2_10_33_port, 
      A_pos_shifted_by2_10_32_port, A_pos_shifted_by2_10_31_port, 
      A_pos_shifted_by2_10_30_port, A_pos_shifted_by2_10_29_port, 
      A_pos_shifted_by2_10_28_port, A_pos_shifted_by2_10_27_port, 
      A_pos_shifted_by2_10_26_port, A_pos_shifted_by2_10_25_port, 
      A_pos_shifted_by2_10_24_port, A_pos_shifted_by2_10_23_port, 
      A_pos_shifted_by2_10_22_port, A_pos_shifted_by2_10_21_port, 
      A_pos_shifted_by2_10_20_port, A_pos_shifted_by2_10_19_port, 
      A_pos_shifted_by2_10_18_port, A_pos_shifted_by2_10_17_port, 
      A_pos_shifted_by2_10_16_port, A_pos_shifted_by2_10_15_port, 
      A_pos_shifted_by2_10_14_port, A_pos_shifted_by2_10_13_port, 
      A_pos_shifted_by2_10_12_port, A_pos_shifted_by2_10_11_port, 
      A_pos_shifted_by2_10_10_port, A_pos_shifted_by2_10_9_port, 
      A_pos_shifted_by2_10_8_port, A_pos_shifted_by2_10_7_port, 
      A_pos_shifted_by2_10_6_port, A_pos_shifted_by2_10_5_port, 
      A_pos_shifted_by2_10_4_port, A_pos_shifted_by2_10_3_port, 
      A_pos_shifted_by2_10_2_port, A_pos_shifted_by2_10_1_port, 
      A_pos_shifted_by2_10_0_port, A_pos_shifted_by2_11_63_port, 
      A_pos_shifted_by2_11_62_port, A_pos_shifted_by2_11_61_port, 
      A_pos_shifted_by2_11_60_port, A_pos_shifted_by2_11_59_port, 
      A_pos_shifted_by2_11_58_port, A_pos_shifted_by2_11_57_port, 
      A_pos_shifted_by2_11_56_port, A_pos_shifted_by2_11_55_port, 
      A_pos_shifted_by2_11_54_port, A_pos_shifted_by2_11_53_port, 
      A_pos_shifted_by2_11_52_port, A_pos_shifted_by2_11_51_port, 
      A_pos_shifted_by2_11_50_port, A_pos_shifted_by2_11_49_port, 
      A_pos_shifted_by2_11_48_port, A_pos_shifted_by2_11_47_port, 
      A_pos_shifted_by2_11_46_port, A_pos_shifted_by2_11_45_port, 
      A_pos_shifted_by2_11_44_port, A_pos_shifted_by2_11_43_port, 
      A_pos_shifted_by2_11_42_port, A_pos_shifted_by2_11_41_port, 
      A_pos_shifted_by2_11_40_port, A_pos_shifted_by2_11_39_port, 
      A_pos_shifted_by2_11_38_port, A_pos_shifted_by2_11_37_port, 
      A_pos_shifted_by2_11_36_port, A_pos_shifted_by2_11_35_port, 
      A_pos_shifted_by2_11_34_port, A_pos_shifted_by2_11_33_port, 
      A_pos_shifted_by2_11_32_port, A_pos_shifted_by2_11_31_port, 
      A_pos_shifted_by2_11_30_port, A_pos_shifted_by2_11_29_port, 
      A_pos_shifted_by2_11_28_port, A_pos_shifted_by2_11_27_port, 
      A_pos_shifted_by2_11_26_port, A_pos_shifted_by2_11_25_port, 
      A_pos_shifted_by2_11_24_port, A_pos_shifted_by2_11_23_port, 
      A_pos_shifted_by2_11_22_port, A_pos_shifted_by2_11_21_port, 
      A_pos_shifted_by2_11_20_port, A_pos_shifted_by2_11_19_port, 
      A_pos_shifted_by2_11_18_port, A_pos_shifted_by2_11_17_port, 
      A_pos_shifted_by2_11_16_port, A_pos_shifted_by2_11_15_port, 
      A_pos_shifted_by2_11_14_port, A_pos_shifted_by2_11_13_port, 
      A_pos_shifted_by2_11_12_port, A_pos_shifted_by2_11_11_port, 
      A_pos_shifted_by2_11_10_port, A_pos_shifted_by2_11_9_port, 
      A_pos_shifted_by2_11_8_port, A_pos_shifted_by2_11_7_port, 
      A_pos_shifted_by2_11_6_port, A_pos_shifted_by2_11_5_port, 
      A_pos_shifted_by2_11_4_port, A_pos_shifted_by2_11_3_port, 
      A_pos_shifted_by2_11_2_port, A_pos_shifted_by2_11_1_port, 
      A_pos_shifted_by2_11_0_port, A_pos_shifted_by2_12_63_port, 
      A_pos_shifted_by2_12_62_port, A_pos_shifted_by2_12_61_port, 
      A_pos_shifted_by2_12_60_port, A_pos_shifted_by2_12_59_port, 
      A_pos_shifted_by2_12_58_port, A_pos_shifted_by2_12_57_port, 
      A_pos_shifted_by2_12_56_port, A_pos_shifted_by2_12_55_port, 
      A_pos_shifted_by2_12_54_port, A_pos_shifted_by2_12_53_port, 
      A_pos_shifted_by2_12_52_port, A_pos_shifted_by2_12_51_port, 
      A_pos_shifted_by2_12_50_port, A_pos_shifted_by2_12_49_port, 
      A_pos_shifted_by2_12_48_port, A_pos_shifted_by2_12_47_port, 
      A_pos_shifted_by2_12_46_port, A_pos_shifted_by2_12_45_port, 
      A_pos_shifted_by2_12_44_port, A_pos_shifted_by2_12_43_port, 
      A_pos_shifted_by2_12_42_port, A_pos_shifted_by2_12_41_port, 
      A_pos_shifted_by2_12_40_port, A_pos_shifted_by2_12_39_port, 
      A_pos_shifted_by2_12_38_port, A_pos_shifted_by2_12_37_port, 
      A_pos_shifted_by2_12_36_port, A_pos_shifted_by2_12_35_port, 
      A_pos_shifted_by2_12_34_port, A_pos_shifted_by2_12_33_port, 
      A_pos_shifted_by2_12_32_port, A_pos_shifted_by2_12_31_port, 
      A_pos_shifted_by2_12_30_port, A_pos_shifted_by2_12_29_port, 
      A_pos_shifted_by2_12_28_port, A_pos_shifted_by2_12_27_port, 
      A_pos_shifted_by2_12_26_port, A_pos_shifted_by2_12_25_port, 
      A_pos_shifted_by2_12_24_port, A_pos_shifted_by2_12_23_port, 
      A_pos_shifted_by2_12_22_port, A_pos_shifted_by2_12_21_port, 
      A_pos_shifted_by2_12_20_port, A_pos_shifted_by2_12_19_port, 
      A_pos_shifted_by2_12_18_port, A_pos_shifted_by2_12_17_port, 
      A_pos_shifted_by2_12_16_port, A_pos_shifted_by2_12_15_port, 
      A_pos_shifted_by2_12_14_port, A_pos_shifted_by2_12_13_port, 
      A_pos_shifted_by2_12_12_port, A_pos_shifted_by2_12_11_port, 
      A_pos_shifted_by2_12_10_port, A_pos_shifted_by2_12_9_port, 
      A_pos_shifted_by2_12_8_port, A_pos_shifted_by2_12_7_port, 
      A_pos_shifted_by2_12_6_port, A_pos_shifted_by2_12_5_port, 
      A_pos_shifted_by2_12_4_port, A_pos_shifted_by2_12_3_port, 
      A_pos_shifted_by2_12_2_port, A_pos_shifted_by2_12_1_port, 
      A_pos_shifted_by2_12_0_port, A_pos_shifted_by2_13_63_port, 
      A_pos_shifted_by2_13_62_port, A_pos_shifted_by2_13_61_port, 
      A_pos_shifted_by2_13_60_port, A_pos_shifted_by2_13_59_port, 
      A_pos_shifted_by2_13_58_port, A_pos_shifted_by2_13_57_port, 
      A_pos_shifted_by2_13_56_port, A_pos_shifted_by2_13_55_port, 
      A_pos_shifted_by2_13_54_port, A_pos_shifted_by2_13_53_port, 
      A_pos_shifted_by2_13_52_port, A_pos_shifted_by2_13_51_port, 
      A_pos_shifted_by2_13_50_port, A_pos_shifted_by2_13_49_port, 
      A_pos_shifted_by2_13_48_port, A_pos_shifted_by2_13_47_port, 
      A_pos_shifted_by2_13_46_port, A_pos_shifted_by2_13_45_port, 
      A_pos_shifted_by2_13_44_port, A_pos_shifted_by2_13_43_port, 
      A_pos_shifted_by2_13_42_port, A_pos_shifted_by2_13_41_port, 
      A_pos_shifted_by2_13_40_port, A_pos_shifted_by2_13_39_port, 
      A_pos_shifted_by2_13_38_port, A_pos_shifted_by2_13_37_port, 
      A_pos_shifted_by2_13_36_port, A_pos_shifted_by2_13_35_port, 
      A_pos_shifted_by2_13_34_port, A_pos_shifted_by2_13_33_port, 
      A_pos_shifted_by2_13_32_port, A_pos_shifted_by2_13_31_port, 
      A_pos_shifted_by2_13_30_port, A_pos_shifted_by2_13_29_port, 
      A_pos_shifted_by2_13_28_port, A_pos_shifted_by2_13_27_port, 
      A_pos_shifted_by2_13_26_port, A_pos_shifted_by2_13_25_port, 
      A_pos_shifted_by2_13_24_port, A_pos_shifted_by2_13_23_port, 
      A_pos_shifted_by2_13_22_port, A_pos_shifted_by2_13_21_port, 
      A_pos_shifted_by2_13_20_port, A_pos_shifted_by2_13_19_port, 
      A_pos_shifted_by2_13_18_port, A_pos_shifted_by2_13_17_port, 
      A_pos_shifted_by2_13_16_port, A_pos_shifted_by2_13_15_port, 
      A_pos_shifted_by2_13_14_port, A_pos_shifted_by2_13_13_port, 
      A_pos_shifted_by2_13_12_port, A_pos_shifted_by2_13_11_port, 
      A_pos_shifted_by2_13_10_port, A_pos_shifted_by2_13_9_port, 
      A_pos_shifted_by2_13_8_port, A_pos_shifted_by2_13_7_port, 
      A_pos_shifted_by2_13_6_port, A_pos_shifted_by2_13_5_port, 
      A_pos_shifted_by2_13_4_port, A_pos_shifted_by2_13_3_port, 
      A_pos_shifted_by2_13_2_port, A_pos_shifted_by2_13_1_port, 
      A_pos_shifted_by2_13_0_port, A_pos_shifted_by2_14_63_port, 
      A_pos_shifted_by2_14_62_port, A_pos_shifted_by2_14_61_port, 
      A_pos_shifted_by2_14_60_port, A_pos_shifted_by2_14_59_port, 
      A_pos_shifted_by2_14_58_port, A_pos_shifted_by2_14_57_port, 
      A_pos_shifted_by2_14_56_port, A_pos_shifted_by2_14_55_port, 
      A_pos_shifted_by2_14_54_port, A_pos_shifted_by2_14_53_port, 
      A_pos_shifted_by2_14_52_port, A_pos_shifted_by2_14_51_port, 
      A_pos_shifted_by2_14_50_port, A_pos_shifted_by2_14_49_port, 
      A_pos_shifted_by2_14_48_port, A_pos_shifted_by2_14_47_port, 
      A_pos_shifted_by2_14_46_port, A_pos_shifted_by2_14_45_port, 
      A_pos_shifted_by2_14_44_port, A_pos_shifted_by2_14_43_port, 
      A_pos_shifted_by2_14_42_port, A_pos_shifted_by2_14_41_port, 
      A_pos_shifted_by2_14_40_port, A_pos_shifted_by2_14_39_port, 
      A_pos_shifted_by2_14_38_port, A_pos_shifted_by2_14_37_port, 
      A_pos_shifted_by2_14_36_port, A_pos_shifted_by2_14_35_port, 
      A_pos_shifted_by2_14_34_port, A_pos_shifted_by2_14_33_port, 
      A_pos_shifted_by2_14_32_port, A_pos_shifted_by2_14_31_port, 
      A_pos_shifted_by2_14_30_port, A_pos_shifted_by2_14_29_port, 
      A_pos_shifted_by2_14_28_port, A_pos_shifted_by2_14_27_port, 
      A_pos_shifted_by2_14_26_port, A_pos_shifted_by2_14_25_port, 
      A_pos_shifted_by2_14_24_port, A_pos_shifted_by2_14_23_port, 
      A_pos_shifted_by2_14_22_port, A_pos_shifted_by2_14_21_port, 
      A_pos_shifted_by2_14_20_port, A_pos_shifted_by2_14_19_port, 
      A_pos_shifted_by2_14_18_port, A_pos_shifted_by2_14_17_port, 
      A_pos_shifted_by2_14_16_port, A_pos_shifted_by2_14_15_port, 
      A_pos_shifted_by2_14_14_port, A_pos_shifted_by2_14_13_port, 
      A_pos_shifted_by2_14_12_port, A_pos_shifted_by2_14_11_port, 
      A_pos_shifted_by2_14_10_port, A_pos_shifted_by2_14_9_port, 
      A_pos_shifted_by2_14_8_port, A_pos_shifted_by2_14_7_port, 
      A_pos_shifted_by2_14_6_port, A_pos_shifted_by2_14_5_port, 
      A_pos_shifted_by2_14_4_port, A_pos_shifted_by2_14_3_port, 
      A_pos_shifted_by2_14_2_port, A_pos_shifted_by2_14_1_port, 
      A_pos_shifted_by2_14_0_port, A_neg_shifted_by1_0_63_port, 
      A_neg_shifted_by1_0_62_port, A_neg_shifted_by1_0_61_port, 
      A_neg_shifted_by1_0_60_port, A_neg_shifted_by1_0_59_port, 
      A_neg_shifted_by1_0_58_port, A_neg_shifted_by1_0_57_port, 
      A_neg_shifted_by1_0_56_port, A_neg_shifted_by1_0_55_port, 
      A_neg_shifted_by1_0_54_port, A_neg_shifted_by1_0_53_port, 
      A_neg_shifted_by1_0_52_port, A_neg_shifted_by1_0_51_port, 
      A_neg_shifted_by1_0_50_port, A_neg_shifted_by1_0_49_port, 
      A_neg_shifted_by1_0_48_port, A_neg_shifted_by1_0_47_port, 
      A_neg_shifted_by1_0_46_port, A_neg_shifted_by1_0_45_port, 
      A_neg_shifted_by1_0_44_port, A_neg_shifted_by1_0_43_port, 
      A_neg_shifted_by1_0_42_port, A_neg_shifted_by1_0_41_port, 
      A_neg_shifted_by1_0_40_port, A_neg_shifted_by1_0_39_port, 
      A_neg_shifted_by1_0_38_port, A_neg_shifted_by1_0_37_port, 
      A_neg_shifted_by1_0_36_port, A_neg_shifted_by1_0_35_port, 
      A_neg_shifted_by1_0_34_port, A_neg_shifted_by1_0_33_port, 
      A_neg_shifted_by1_0_32_port, A_neg_shifted_by1_0_31_port, 
      A_neg_shifted_by1_0_30_port, A_neg_shifted_by1_0_29_port, 
      A_neg_shifted_by1_0_28_port, A_neg_shifted_by1_0_27_port, 
      A_neg_shifted_by1_0_26_port, A_neg_shifted_by1_0_25_port, 
      A_neg_shifted_by1_0_24_port, A_neg_shifted_by1_0_23_port, 
      A_neg_shifted_by1_0_22_port, A_neg_shifted_by1_0_21_port, 
      A_neg_shifted_by1_0_20_port, A_neg_shifted_by1_0_19_port, 
      A_neg_shifted_by1_0_18_port, A_neg_shifted_by1_0_17_port, 
      A_neg_shifted_by1_0_16_port, A_neg_shifted_by1_0_15_port, 
      A_neg_shifted_by1_0_14_port, A_neg_shifted_by1_0_13_port, 
      A_neg_shifted_by1_0_12_port, A_neg_shifted_by1_0_11_port, 
      A_neg_shifted_by1_0_10_port, A_neg_shifted_by1_0_9_port, 
      A_neg_shifted_by1_0_8_port, A_neg_shifted_by1_0_7_port, 
      A_neg_shifted_by1_0_6_port, A_neg_shifted_by1_0_5_port, 
      A_neg_shifted_by1_0_4_port, A_neg_shifted_by1_0_3_port, 
      A_neg_shifted_by1_0_2_port, A_neg_shifted_by1_0_1_port, 
      A_neg_shifted_by1_0_0_port, A_neg_shifted_by1_1_63_port, 
      A_neg_shifted_by1_1_62_port, A_neg_shifted_by1_1_61_port, 
      A_neg_shifted_by1_1_60_port, A_neg_shifted_by1_1_59_port, 
      A_neg_shifted_by1_1_58_port, A_neg_shifted_by1_1_57_port, 
      A_neg_shifted_by1_1_56_port, A_neg_shifted_by1_1_55_port, 
      A_neg_shifted_by1_1_54_port, A_neg_shifted_by1_1_53_port, 
      A_neg_shifted_by1_1_52_port, A_neg_shifted_by1_1_51_port, 
      A_neg_shifted_by1_1_50_port, A_neg_shifted_by1_1_49_port, 
      A_neg_shifted_by1_1_48_port, A_neg_shifted_by1_1_47_port, 
      A_neg_shifted_by1_1_46_port, A_neg_shifted_by1_1_45_port, 
      A_neg_shifted_by1_1_44_port, A_neg_shifted_by1_1_43_port, 
      A_neg_shifted_by1_1_42_port, A_neg_shifted_by1_1_41_port, 
      A_neg_shifted_by1_1_40_port, A_neg_shifted_by1_1_39_port, 
      A_neg_shifted_by1_1_38_port, A_neg_shifted_by1_1_37_port, 
      A_neg_shifted_by1_1_36_port, A_neg_shifted_by1_1_35_port, 
      A_neg_shifted_by1_1_34_port, A_neg_shifted_by1_1_33_port, 
      A_neg_shifted_by1_1_32_port, A_neg_shifted_by1_1_31_port, 
      A_neg_shifted_by1_1_30_port, A_neg_shifted_by1_1_29_port, 
      A_neg_shifted_by1_1_28_port, A_neg_shifted_by1_1_27_port, 
      A_neg_shifted_by1_1_26_port, A_neg_shifted_by1_1_25_port, 
      A_neg_shifted_by1_1_24_port, A_neg_shifted_by1_1_23_port, 
      A_neg_shifted_by1_1_22_port, A_neg_shifted_by1_1_21_port, 
      A_neg_shifted_by1_1_20_port, A_neg_shifted_by1_1_19_port, 
      A_neg_shifted_by1_1_18_port, A_neg_shifted_by1_1_17_port, 
      A_neg_shifted_by1_1_16_port, A_neg_shifted_by1_1_15_port, 
      A_neg_shifted_by1_1_14_port, A_neg_shifted_by1_1_13_port, 
      A_neg_shifted_by1_1_12_port, A_neg_shifted_by1_1_11_port, 
      A_neg_shifted_by1_1_10_port, A_neg_shifted_by1_1_9_port, 
      A_neg_shifted_by1_1_8_port, A_neg_shifted_by1_1_7_port, 
      A_neg_shifted_by1_1_6_port, A_neg_shifted_by1_1_5_port, 
      A_neg_shifted_by1_1_4_port, A_neg_shifted_by1_1_3_port, 
      A_neg_shifted_by1_1_2_port, A_neg_shifted_by1_1_1_port, 
      A_neg_shifted_by1_1_0_port, A_neg_shifted_by1_2_63_port, 
      A_neg_shifted_by1_2_62_port, A_neg_shifted_by1_2_61_port, 
      A_neg_shifted_by1_2_60_port, A_neg_shifted_by1_2_59_port, 
      A_neg_shifted_by1_2_58_port, A_neg_shifted_by1_2_57_port, 
      A_neg_shifted_by1_2_56_port, A_neg_shifted_by1_2_55_port, 
      A_neg_shifted_by1_2_54_port, A_neg_shifted_by1_2_53_port, 
      A_neg_shifted_by1_2_52_port, A_neg_shifted_by1_2_51_port, 
      A_neg_shifted_by1_2_50_port, A_neg_shifted_by1_2_49_port, 
      A_neg_shifted_by1_2_48_port, A_neg_shifted_by1_2_47_port, 
      A_neg_shifted_by1_2_46_port, A_neg_shifted_by1_2_45_port, 
      A_neg_shifted_by1_2_44_port, A_neg_shifted_by1_2_43_port, 
      A_neg_shifted_by1_2_42_port, A_neg_shifted_by1_2_41_port, 
      A_neg_shifted_by1_2_40_port, A_neg_shifted_by1_2_39_port, 
      A_neg_shifted_by1_2_38_port, A_neg_shifted_by1_2_37_port, 
      A_neg_shifted_by1_2_36_port, A_neg_shifted_by1_2_35_port, 
      A_neg_shifted_by1_2_34_port, A_neg_shifted_by1_2_33_port, 
      A_neg_shifted_by1_2_32_port, A_neg_shifted_by1_2_31_port, 
      A_neg_shifted_by1_2_30_port, A_neg_shifted_by1_2_29_port, 
      A_neg_shifted_by1_2_28_port, A_neg_shifted_by1_2_27_port, 
      A_neg_shifted_by1_2_26_port, A_neg_shifted_by1_2_25_port, 
      A_neg_shifted_by1_2_24_port, A_neg_shifted_by1_2_23_port, 
      A_neg_shifted_by1_2_22_port, A_neg_shifted_by1_2_21_port, 
      A_neg_shifted_by1_2_20_port, A_neg_shifted_by1_2_19_port, 
      A_neg_shifted_by1_2_18_port, A_neg_shifted_by1_2_17_port, 
      A_neg_shifted_by1_2_16_port, A_neg_shifted_by1_2_15_port, 
      A_neg_shifted_by1_2_14_port, A_neg_shifted_by1_2_13_port, 
      A_neg_shifted_by1_2_12_port, A_neg_shifted_by1_2_11_port, 
      A_neg_shifted_by1_2_10_port, A_neg_shifted_by1_2_9_port, 
      A_neg_shifted_by1_2_8_port, A_neg_shifted_by1_2_7_port, 
      A_neg_shifted_by1_2_6_port, A_neg_shifted_by1_2_5_port, 
      A_neg_shifted_by1_2_4_port, A_neg_shifted_by1_2_3_port, 
      A_neg_shifted_by1_2_2_port, A_neg_shifted_by1_2_1_port, 
      A_neg_shifted_by1_2_0_port, A_neg_shifted_by1_3_63_port, 
      A_neg_shifted_by1_3_62_port, A_neg_shifted_by1_3_61_port, 
      A_neg_shifted_by1_3_60_port, A_neg_shifted_by1_3_59_port, 
      A_neg_shifted_by1_3_58_port, A_neg_shifted_by1_3_57_port, 
      A_neg_shifted_by1_3_56_port, A_neg_shifted_by1_3_55_port, 
      A_neg_shifted_by1_3_54_port, A_neg_shifted_by1_3_53_port, 
      A_neg_shifted_by1_3_52_port, A_neg_shifted_by1_3_51_port, 
      A_neg_shifted_by1_3_50_port, A_neg_shifted_by1_3_49_port, 
      A_neg_shifted_by1_3_48_port, A_neg_shifted_by1_3_47_port, 
      A_neg_shifted_by1_3_46_port, A_neg_shifted_by1_3_45_port, 
      A_neg_shifted_by1_3_44_port, A_neg_shifted_by1_3_43_port, 
      A_neg_shifted_by1_3_42_port, A_neg_shifted_by1_3_41_port, 
      A_neg_shifted_by1_3_40_port, A_neg_shifted_by1_3_39_port, 
      A_neg_shifted_by1_3_38_port, A_neg_shifted_by1_3_37_port, 
      A_neg_shifted_by1_3_36_port, A_neg_shifted_by1_3_35_port, 
      A_neg_shifted_by1_3_34_port, A_neg_shifted_by1_3_33_port, 
      A_neg_shifted_by1_3_32_port, A_neg_shifted_by1_3_31_port, 
      A_neg_shifted_by1_3_30_port, A_neg_shifted_by1_3_29_port, 
      A_neg_shifted_by1_3_28_port, A_neg_shifted_by1_3_27_port, 
      A_neg_shifted_by1_3_26_port, A_neg_shifted_by1_3_25_port, 
      A_neg_shifted_by1_3_24_port, A_neg_shifted_by1_3_23_port, 
      A_neg_shifted_by1_3_22_port, A_neg_shifted_by1_3_21_port, 
      A_neg_shifted_by1_3_20_port, A_neg_shifted_by1_3_19_port, 
      A_neg_shifted_by1_3_18_port, A_neg_shifted_by1_3_17_port, 
      A_neg_shifted_by1_3_16_port, A_neg_shifted_by1_3_15_port, 
      A_neg_shifted_by1_3_14_port, A_neg_shifted_by1_3_13_port, 
      A_neg_shifted_by1_3_12_port, A_neg_shifted_by1_3_11_port, 
      A_neg_shifted_by1_3_10_port, A_neg_shifted_by1_3_9_port, 
      A_neg_shifted_by1_3_8_port, A_neg_shifted_by1_3_7_port, 
      A_neg_shifted_by1_3_6_port, A_neg_shifted_by1_3_5_port, 
      A_neg_shifted_by1_3_4_port, A_neg_shifted_by1_3_3_port, 
      A_neg_shifted_by1_3_2_port, A_neg_shifted_by1_3_1_port, 
      A_neg_shifted_by1_3_0_port, A_neg_shifted_by1_4_63_port, 
      A_neg_shifted_by1_4_62_port, A_neg_shifted_by1_4_61_port, 
      A_neg_shifted_by1_4_60_port, A_neg_shifted_by1_4_59_port, 
      A_neg_shifted_by1_4_58_port, A_neg_shifted_by1_4_57_port, 
      A_neg_shifted_by1_4_56_port, A_neg_shifted_by1_4_55_port, 
      A_neg_shifted_by1_4_54_port, A_neg_shifted_by1_4_53_port, 
      A_neg_shifted_by1_4_52_port, A_neg_shifted_by1_4_51_port, 
      A_neg_shifted_by1_4_50_port, A_neg_shifted_by1_4_49_port, 
      A_neg_shifted_by1_4_48_port, A_neg_shifted_by1_4_47_port, 
      A_neg_shifted_by1_4_46_port, A_neg_shifted_by1_4_45_port, 
      A_neg_shifted_by1_4_44_port, A_neg_shifted_by1_4_43_port, 
      A_neg_shifted_by1_4_42_port, A_neg_shifted_by1_4_41_port, 
      A_neg_shifted_by1_4_40_port, A_neg_shifted_by1_4_39_port, 
      A_neg_shifted_by1_4_38_port, A_neg_shifted_by1_4_37_port, 
      A_neg_shifted_by1_4_36_port, A_neg_shifted_by1_4_35_port, 
      A_neg_shifted_by1_4_34_port, A_neg_shifted_by1_4_33_port, 
      A_neg_shifted_by1_4_32_port, A_neg_shifted_by1_4_31_port, 
      A_neg_shifted_by1_4_30_port, A_neg_shifted_by1_4_29_port, 
      A_neg_shifted_by1_4_28_port, A_neg_shifted_by1_4_27_port, 
      A_neg_shifted_by1_4_26_port, A_neg_shifted_by1_4_25_port, 
      A_neg_shifted_by1_4_24_port, A_neg_shifted_by1_4_23_port, 
      A_neg_shifted_by1_4_22_port, A_neg_shifted_by1_4_21_port, 
      A_neg_shifted_by1_4_20_port, A_neg_shifted_by1_4_19_port, 
      A_neg_shifted_by1_4_18_port, A_neg_shifted_by1_4_17_port, 
      A_neg_shifted_by1_4_16_port, A_neg_shifted_by1_4_15_port, 
      A_neg_shifted_by1_4_14_port, A_neg_shifted_by1_4_13_port, 
      A_neg_shifted_by1_4_12_port, A_neg_shifted_by1_4_11_port, 
      A_neg_shifted_by1_4_10_port, A_neg_shifted_by1_4_9_port, 
      A_neg_shifted_by1_4_8_port, A_neg_shifted_by1_4_7_port, 
      A_neg_shifted_by1_4_6_port, A_neg_shifted_by1_4_5_port, 
      A_neg_shifted_by1_4_4_port, A_neg_shifted_by1_4_3_port, 
      A_neg_shifted_by1_4_2_port, A_neg_shifted_by1_4_1_port, 
      A_neg_shifted_by1_4_0_port, A_neg_shifted_by1_5_63_port, 
      A_neg_shifted_by1_5_62_port, A_neg_shifted_by1_5_61_port, 
      A_neg_shifted_by1_5_60_port, A_neg_shifted_by1_5_59_port, 
      A_neg_shifted_by1_5_58_port, A_neg_shifted_by1_5_57_port, 
      A_neg_shifted_by1_5_56_port, A_neg_shifted_by1_5_55_port, 
      A_neg_shifted_by1_5_54_port, A_neg_shifted_by1_5_53_port, 
      A_neg_shifted_by1_5_52_port, A_neg_shifted_by1_5_51_port, 
      A_neg_shifted_by1_5_50_port, A_neg_shifted_by1_5_49_port, 
      A_neg_shifted_by1_5_48_port, A_neg_shifted_by1_5_47_port, 
      A_neg_shifted_by1_5_46_port, A_neg_shifted_by1_5_45_port, 
      A_neg_shifted_by1_5_44_port, A_neg_shifted_by1_5_43_port, 
      A_neg_shifted_by1_5_42_port, A_neg_shifted_by1_5_41_port, 
      A_neg_shifted_by1_5_40_port, A_neg_shifted_by1_5_39_port, 
      A_neg_shifted_by1_5_38_port, A_neg_shifted_by1_5_37_port, 
      A_neg_shifted_by1_5_36_port, A_neg_shifted_by1_5_35_port, 
      A_neg_shifted_by1_5_34_port, A_neg_shifted_by1_5_33_port, 
      A_neg_shifted_by1_5_32_port, A_neg_shifted_by1_5_31_port, 
      A_neg_shifted_by1_5_30_port, A_neg_shifted_by1_5_29_port, 
      A_neg_shifted_by1_5_28_port, A_neg_shifted_by1_5_27_port, 
      A_neg_shifted_by1_5_26_port, A_neg_shifted_by1_5_25_port, 
      A_neg_shifted_by1_5_24_port, A_neg_shifted_by1_5_23_port, 
      A_neg_shifted_by1_5_22_port, A_neg_shifted_by1_5_21_port, 
      A_neg_shifted_by1_5_20_port, A_neg_shifted_by1_5_19_port, 
      A_neg_shifted_by1_5_18_port, A_neg_shifted_by1_5_17_port, 
      A_neg_shifted_by1_5_16_port, A_neg_shifted_by1_5_15_port, 
      A_neg_shifted_by1_5_14_port, A_neg_shifted_by1_5_13_port, 
      A_neg_shifted_by1_5_12_port, A_neg_shifted_by1_5_11_port, 
      A_neg_shifted_by1_5_10_port, A_neg_shifted_by1_5_9_port, 
      A_neg_shifted_by1_5_8_port, A_neg_shifted_by1_5_7_port, 
      A_neg_shifted_by1_5_6_port, A_neg_shifted_by1_5_5_port, 
      A_neg_shifted_by1_5_4_port, A_neg_shifted_by1_5_3_port, 
      A_neg_shifted_by1_5_2_port, A_neg_shifted_by1_5_1_port, 
      A_neg_shifted_by1_5_0_port, A_neg_shifted_by1_6_63_port, 
      A_neg_shifted_by1_6_62_port, A_neg_shifted_by1_6_61_port, 
      A_neg_shifted_by1_6_60_port, A_neg_shifted_by1_6_59_port, 
      A_neg_shifted_by1_6_58_port, A_neg_shifted_by1_6_57_port, 
      A_neg_shifted_by1_6_56_port, A_neg_shifted_by1_6_55_port, 
      A_neg_shifted_by1_6_54_port, A_neg_shifted_by1_6_53_port, 
      A_neg_shifted_by1_6_52_port, A_neg_shifted_by1_6_51_port, 
      A_neg_shifted_by1_6_50_port, A_neg_shifted_by1_6_49_port, 
      A_neg_shifted_by1_6_48_port, A_neg_shifted_by1_6_47_port, 
      A_neg_shifted_by1_6_46_port, A_neg_shifted_by1_6_45_port, 
      A_neg_shifted_by1_6_44_port, A_neg_shifted_by1_6_43_port, 
      A_neg_shifted_by1_6_42_port, A_neg_shifted_by1_6_41_port, 
      A_neg_shifted_by1_6_40_port, A_neg_shifted_by1_6_39_port, 
      A_neg_shifted_by1_6_38_port, A_neg_shifted_by1_6_37_port, 
      A_neg_shifted_by1_6_36_port, A_neg_shifted_by1_6_35_port, 
      A_neg_shifted_by1_6_34_port, A_neg_shifted_by1_6_33_port, 
      A_neg_shifted_by1_6_32_port, A_neg_shifted_by1_6_31_port, 
      A_neg_shifted_by1_6_30_port, A_neg_shifted_by1_6_29_port, 
      A_neg_shifted_by1_6_28_port, A_neg_shifted_by1_6_27_port, 
      A_neg_shifted_by1_6_26_port, A_neg_shifted_by1_6_25_port, 
      A_neg_shifted_by1_6_24_port, A_neg_shifted_by1_6_23_port, 
      A_neg_shifted_by1_6_22_port, A_neg_shifted_by1_6_21_port, 
      A_neg_shifted_by1_6_20_port, A_neg_shifted_by1_6_19_port, 
      A_neg_shifted_by1_6_18_port, A_neg_shifted_by1_6_17_port, 
      A_neg_shifted_by1_6_16_port, A_neg_shifted_by1_6_15_port, 
      A_neg_shifted_by1_6_14_port, A_neg_shifted_by1_6_13_port, 
      A_neg_shifted_by1_6_12_port, A_neg_shifted_by1_6_11_port, 
      A_neg_shifted_by1_6_10_port, A_neg_shifted_by1_6_9_port, 
      A_neg_shifted_by1_6_8_port, A_neg_shifted_by1_6_7_port, 
      A_neg_shifted_by1_6_6_port, A_neg_shifted_by1_6_5_port, 
      A_neg_shifted_by1_6_4_port, A_neg_shifted_by1_6_3_port, 
      A_neg_shifted_by1_6_2_port, A_neg_shifted_by1_6_1_port, 
      A_neg_shifted_by1_6_0_port, A_neg_shifted_by1_7_63_port, 
      A_neg_shifted_by1_7_62_port, A_neg_shifted_by1_7_61_port, 
      A_neg_shifted_by1_7_60_port, A_neg_shifted_by1_7_59_port, 
      A_neg_shifted_by1_7_58_port, A_neg_shifted_by1_7_57_port, 
      A_neg_shifted_by1_7_56_port, A_neg_shifted_by1_7_55_port, 
      A_neg_shifted_by1_7_54_port, A_neg_shifted_by1_7_53_port, 
      A_neg_shifted_by1_7_52_port, A_neg_shifted_by1_7_51_port, 
      A_neg_shifted_by1_7_50_port, A_neg_shifted_by1_7_49_port, 
      A_neg_shifted_by1_7_48_port, A_neg_shifted_by1_7_47_port, 
      A_neg_shifted_by1_7_46_port, A_neg_shifted_by1_7_45_port, 
      A_neg_shifted_by1_7_44_port, A_neg_shifted_by1_7_43_port, 
      A_neg_shifted_by1_7_42_port, A_neg_shifted_by1_7_41_port, 
      A_neg_shifted_by1_7_40_port, A_neg_shifted_by1_7_39_port, 
      A_neg_shifted_by1_7_38_port, A_neg_shifted_by1_7_37_port, 
      A_neg_shifted_by1_7_36_port, A_neg_shifted_by1_7_35_port, 
      A_neg_shifted_by1_7_34_port, A_neg_shifted_by1_7_33_port, 
      A_neg_shifted_by1_7_32_port, A_neg_shifted_by1_7_31_port, 
      A_neg_shifted_by1_7_30_port, A_neg_shifted_by1_7_29_port, 
      A_neg_shifted_by1_7_28_port, A_neg_shifted_by1_7_27_port, 
      A_neg_shifted_by1_7_26_port, A_neg_shifted_by1_7_25_port, 
      A_neg_shifted_by1_7_24_port, A_neg_shifted_by1_7_23_port, 
      A_neg_shifted_by1_7_22_port, A_neg_shifted_by1_7_21_port, 
      A_neg_shifted_by1_7_20_port, A_neg_shifted_by1_7_19_port, 
      A_neg_shifted_by1_7_18_port, A_neg_shifted_by1_7_17_port, 
      A_neg_shifted_by1_7_16_port, A_neg_shifted_by1_7_15_port, 
      A_neg_shifted_by1_7_14_port, A_neg_shifted_by1_7_13_port, 
      A_neg_shifted_by1_7_12_port, A_neg_shifted_by1_7_11_port, 
      A_neg_shifted_by1_7_10_port, A_neg_shifted_by1_7_9_port, 
      A_neg_shifted_by1_7_8_port, A_neg_shifted_by1_7_7_port, 
      A_neg_shifted_by1_7_6_port, A_neg_shifted_by1_7_5_port, 
      A_neg_shifted_by1_7_4_port, A_neg_shifted_by1_7_3_port, 
      A_neg_shifted_by1_7_2_port, A_neg_shifted_by1_7_1_port, 
      A_neg_shifted_by1_7_0_port, A_neg_shifted_by2_0_63_port, 
      A_neg_shifted_by2_0_62_port, A_neg_shifted_by2_0_61_port, 
      A_neg_shifted_by2_0_60_port, A_neg_shifted_by2_0_59_port, 
      A_neg_shifted_by2_0_58_port, A_neg_shifted_by2_0_57_port, 
      A_neg_shifted_by2_0_56_port, A_neg_shifted_by2_0_55_port, 
      A_neg_shifted_by2_0_54_port, A_neg_shifted_by2_0_53_port, 
      A_neg_shifted_by2_0_52_port, A_neg_shifted_by2_0_51_port, 
      A_neg_shifted_by2_0_50_port, A_neg_shifted_by2_0_49_port, 
      A_neg_shifted_by2_0_48_port, A_neg_shifted_by2_0_47_port, 
      A_neg_shifted_by2_0_46_port, A_neg_shifted_by2_0_45_port, 
      A_neg_shifted_by2_0_44_port, A_neg_shifted_by2_0_43_port, 
      A_neg_shifted_by2_0_42_port, A_neg_shifted_by2_0_41_port, 
      A_neg_shifted_by2_0_40_port, A_neg_shifted_by2_0_39_port, 
      A_neg_shifted_by2_0_38_port, A_neg_shifted_by2_0_37_port, 
      A_neg_shifted_by2_0_36_port, A_neg_shifted_by2_0_35_port, 
      A_neg_shifted_by2_0_34_port, A_neg_shifted_by2_0_33_port, 
      A_neg_shifted_by2_0_32_port, A_neg_shifted_by2_0_31_port, 
      A_neg_shifted_by2_0_30_port, A_neg_shifted_by2_0_29_port, 
      A_neg_shifted_by2_0_28_port, A_neg_shifted_by2_0_27_port, 
      A_neg_shifted_by2_0_26_port, A_neg_shifted_by2_0_25_port, 
      A_neg_shifted_by2_0_24_port, A_neg_shifted_by2_0_23_port, 
      A_neg_shifted_by2_0_22_port, A_neg_shifted_by2_0_21_port, 
      A_neg_shifted_by2_0_20_port, A_neg_shifted_by2_0_19_port, 
      A_neg_shifted_by2_0_18_port, A_neg_shifted_by2_0_17_port, 
      A_neg_shifted_by2_0_16_port, A_neg_shifted_by2_0_15_port, 
      A_neg_shifted_by2_0_14_port, A_neg_shifted_by2_0_13_port, 
      A_neg_shifted_by2_0_12_port, A_neg_shifted_by2_0_11_port, 
      A_neg_shifted_by2_0_10_port, A_neg_shifted_by2_0_9_port, 
      A_neg_shifted_by2_0_8_port, A_neg_shifted_by2_0_7_port, 
      A_neg_shifted_by2_0_6_port, A_neg_shifted_by2_0_5_port, 
      A_neg_shifted_by2_0_4_port, A_neg_shifted_by2_0_3_port, 
      A_neg_shifted_by2_0_2_port, A_neg_shifted_by2_0_1_port, 
      A_neg_shifted_by2_0_0_port, A_neg_shifted_by2_1_63_port, 
      A_neg_shifted_by2_1_62_port, A_neg_shifted_by2_1_61_port, 
      A_neg_shifted_by2_1_60_port, A_neg_shifted_by2_1_59_port, 
      A_neg_shifted_by2_1_58_port, A_neg_shifted_by2_1_57_port, 
      A_neg_shifted_by2_1_56_port, A_neg_shifted_by2_1_55_port, 
      A_neg_shifted_by2_1_54_port, A_neg_shifted_by2_1_53_port, 
      A_neg_shifted_by2_1_52_port, A_neg_shifted_by2_1_51_port, 
      A_neg_shifted_by2_1_50_port, A_neg_shifted_by2_1_49_port, 
      A_neg_shifted_by2_1_48_port, A_neg_shifted_by2_1_47_port, 
      A_neg_shifted_by2_1_46_port, A_neg_shifted_by2_1_45_port, 
      A_neg_shifted_by2_1_44_port, A_neg_shifted_by2_1_43_port, 
      A_neg_shifted_by2_1_42_port, A_neg_shifted_by2_1_41_port, 
      A_neg_shifted_by2_1_40_port, A_neg_shifted_by2_1_39_port, 
      A_neg_shifted_by2_1_38_port, A_neg_shifted_by2_1_37_port, 
      A_neg_shifted_by2_1_36_port, A_neg_shifted_by2_1_35_port, 
      A_neg_shifted_by2_1_34_port, A_neg_shifted_by2_1_33_port, 
      A_neg_shifted_by2_1_32_port, A_neg_shifted_by2_1_31_port, 
      A_neg_shifted_by2_1_30_port, A_neg_shifted_by2_1_29_port, 
      A_neg_shifted_by2_1_28_port, A_neg_shifted_by2_1_27_port, 
      A_neg_shifted_by2_1_26_port, A_neg_shifted_by2_1_25_port, 
      A_neg_shifted_by2_1_24_port, A_neg_shifted_by2_1_23_port, 
      A_neg_shifted_by2_1_22_port, A_neg_shifted_by2_1_21_port, 
      A_neg_shifted_by2_1_20_port, A_neg_shifted_by2_1_19_port, 
      A_neg_shifted_by2_1_18_port, A_neg_shifted_by2_1_17_port, 
      A_neg_shifted_by2_1_16_port, A_neg_shifted_by2_1_15_port, 
      A_neg_shifted_by2_1_14_port, A_neg_shifted_by2_1_13_port, 
      A_neg_shifted_by2_1_12_port, A_neg_shifted_by2_1_11_port, 
      A_neg_shifted_by2_1_10_port, A_neg_shifted_by2_1_9_port, 
      A_neg_shifted_by2_1_8_port, A_neg_shifted_by2_1_7_port, 
      A_neg_shifted_by2_1_6_port, A_neg_shifted_by2_1_5_port, 
      A_neg_shifted_by2_1_4_port, A_neg_shifted_by2_1_3_port, 
      A_neg_shifted_by2_1_2_port, A_neg_shifted_by2_1_1_port, 
      A_neg_shifted_by2_1_0_port, A_neg_shifted_by2_2_63_port, 
      A_neg_shifted_by2_2_62_port, A_neg_shifted_by2_2_61_port, 
      A_neg_shifted_by2_2_60_port, A_neg_shifted_by2_2_59_port, 
      A_neg_shifted_by2_2_58_port, A_neg_shifted_by2_2_57_port, 
      A_neg_shifted_by2_2_56_port, A_neg_shifted_by2_2_55_port, 
      A_neg_shifted_by2_2_54_port, A_neg_shifted_by2_2_53_port, 
      A_neg_shifted_by2_2_52_port, A_neg_shifted_by2_2_51_port, 
      A_neg_shifted_by2_2_50_port, A_neg_shifted_by2_2_49_port, 
      A_neg_shifted_by2_2_48_port, A_neg_shifted_by2_2_47_port, 
      A_neg_shifted_by2_2_46_port, A_neg_shifted_by2_2_45_port, 
      A_neg_shifted_by2_2_44_port, A_neg_shifted_by2_2_43_port, 
      A_neg_shifted_by2_2_42_port, A_neg_shifted_by2_2_41_port, 
      A_neg_shifted_by2_2_40_port, A_neg_shifted_by2_2_39_port, 
      A_neg_shifted_by2_2_38_port, A_neg_shifted_by2_2_37_port, 
      A_neg_shifted_by2_2_36_port, A_neg_shifted_by2_2_35_port, 
      A_neg_shifted_by2_2_34_port, A_neg_shifted_by2_2_33_port, 
      A_neg_shifted_by2_2_32_port, A_neg_shifted_by2_2_31_port, 
      A_neg_shifted_by2_2_30_port, A_neg_shifted_by2_2_29_port, 
      A_neg_shifted_by2_2_28_port, A_neg_shifted_by2_2_27_port, 
      A_neg_shifted_by2_2_26_port, A_neg_shifted_by2_2_25_port, 
      A_neg_shifted_by2_2_24_port, A_neg_shifted_by2_2_23_port, 
      A_neg_shifted_by2_2_22_port, A_neg_shifted_by2_2_21_port, 
      A_neg_shifted_by2_2_20_port, A_neg_shifted_by2_2_19_port, 
      A_neg_shifted_by2_2_18_port, A_neg_shifted_by2_2_17_port, 
      A_neg_shifted_by2_2_16_port, A_neg_shifted_by2_2_15_port, 
      A_neg_shifted_by2_2_14_port, A_neg_shifted_by2_2_13_port, 
      A_neg_shifted_by2_2_12_port, A_neg_shifted_by2_2_11_port, 
      A_neg_shifted_by2_2_10_port, A_neg_shifted_by2_2_9_port, 
      A_neg_shifted_by2_2_8_port, A_neg_shifted_by2_2_7_port, 
      A_neg_shifted_by2_2_6_port, A_neg_shifted_by2_2_5_port, 
      A_neg_shifted_by2_2_4_port, A_neg_shifted_by2_2_3_port, 
      A_neg_shifted_by2_2_2_port, A_neg_shifted_by2_2_1_port, 
      A_neg_shifted_by2_2_0_port, A_neg_shifted_by2_3_63_port, 
      A_neg_shifted_by2_3_62_port, A_neg_shifted_by2_3_61_port, 
      A_neg_shifted_by2_3_60_port, A_neg_shifted_by2_3_59_port, 
      A_neg_shifted_by2_3_58_port, A_neg_shifted_by2_3_57_port, 
      A_neg_shifted_by2_3_56_port, A_neg_shifted_by2_3_55_port, 
      A_neg_shifted_by2_3_54_port, A_neg_shifted_by2_3_53_port, 
      A_neg_shifted_by2_3_52_port, A_neg_shifted_by2_3_51_port, 
      A_neg_shifted_by2_3_50_port, A_neg_shifted_by2_3_49_port, 
      A_neg_shifted_by2_3_48_port, A_neg_shifted_by2_3_47_port, 
      A_neg_shifted_by2_3_46_port, A_neg_shifted_by2_3_45_port, 
      A_neg_shifted_by2_3_44_port, A_neg_shifted_by2_3_43_port, 
      A_neg_shifted_by2_3_42_port, A_neg_shifted_by2_3_41_port, 
      A_neg_shifted_by2_3_40_port, A_neg_shifted_by2_3_39_port, 
      A_neg_shifted_by2_3_38_port, A_neg_shifted_by2_3_37_port, 
      A_neg_shifted_by2_3_36_port, A_neg_shifted_by2_3_35_port, 
      A_neg_shifted_by2_3_34_port, A_neg_shifted_by2_3_33_port, 
      A_neg_shifted_by2_3_32_port, A_neg_shifted_by2_3_31_port, 
      A_neg_shifted_by2_3_30_port, A_neg_shifted_by2_3_29_port, 
      A_neg_shifted_by2_3_28_port, A_neg_shifted_by2_3_27_port, 
      A_neg_shifted_by2_3_26_port, A_neg_shifted_by2_3_25_port, 
      A_neg_shifted_by2_3_24_port, A_neg_shifted_by2_3_23_port, 
      A_neg_shifted_by2_3_22_port, A_neg_shifted_by2_3_21_port, 
      A_neg_shifted_by2_3_20_port, A_neg_shifted_by2_3_19_port, 
      A_neg_shifted_by2_3_18_port, A_neg_shifted_by2_3_17_port, 
      A_neg_shifted_by2_3_16_port, A_neg_shifted_by2_3_15_port, 
      A_neg_shifted_by2_3_14_port, A_neg_shifted_by2_3_13_port, 
      A_neg_shifted_by2_3_12_port, A_neg_shifted_by2_3_11_port, 
      A_neg_shifted_by2_3_10_port, A_neg_shifted_by2_3_9_port, 
      A_neg_shifted_by2_3_8_port, A_neg_shifted_by2_3_7_port, 
      A_neg_shifted_by2_3_6_port, A_neg_shifted_by2_3_5_port, 
      A_neg_shifted_by2_3_4_port, A_neg_shifted_by2_3_3_port, 
      A_neg_shifted_by2_3_2_port, A_neg_shifted_by2_3_1_port, 
      A_neg_shifted_by2_3_0_port, A_neg_shifted_by2_4_63_port, 
      A_neg_shifted_by2_4_62_port, A_neg_shifted_by2_4_61_port, 
      A_neg_shifted_by2_4_60_port, A_neg_shifted_by2_4_59_port, 
      A_neg_shifted_by2_4_58_port, A_neg_shifted_by2_4_57_port, 
      A_neg_shifted_by2_4_56_port, A_neg_shifted_by2_4_55_port, 
      A_neg_shifted_by2_4_54_port, A_neg_shifted_by2_4_53_port, 
      A_neg_shifted_by2_4_52_port, A_neg_shifted_by2_4_51_port, 
      A_neg_shifted_by2_4_50_port, A_neg_shifted_by2_4_49_port, 
      A_neg_shifted_by2_4_48_port, A_neg_shifted_by2_4_47_port, 
      A_neg_shifted_by2_4_46_port, A_neg_shifted_by2_4_45_port, 
      A_neg_shifted_by2_4_44_port, A_neg_shifted_by2_4_43_port, 
      A_neg_shifted_by2_4_42_port, A_neg_shifted_by2_4_41_port, 
      A_neg_shifted_by2_4_40_port, A_neg_shifted_by2_4_39_port, 
      A_neg_shifted_by2_4_38_port, A_neg_shifted_by2_4_37_port, 
      A_neg_shifted_by2_4_36_port, A_neg_shifted_by2_4_35_port, 
      A_neg_shifted_by2_4_34_port, A_neg_shifted_by2_4_33_port, 
      A_neg_shifted_by2_4_32_port, A_neg_shifted_by2_4_31_port, 
      A_neg_shifted_by2_4_30_port, A_neg_shifted_by2_4_29_port, 
      A_neg_shifted_by2_4_28_port, A_neg_shifted_by2_4_27_port, 
      A_neg_shifted_by2_4_26_port, A_neg_shifted_by2_4_25_port, 
      A_neg_shifted_by2_4_24_port, A_neg_shifted_by2_4_23_port, 
      A_neg_shifted_by2_4_22_port, A_neg_shifted_by2_4_21_port, 
      A_neg_shifted_by2_4_20_port, A_neg_shifted_by2_4_19_port, 
      A_neg_shifted_by2_4_18_port, A_neg_shifted_by2_4_17_port, 
      A_neg_shifted_by2_4_16_port, A_neg_shifted_by2_4_15_port, 
      A_neg_shifted_by2_4_14_port, A_neg_shifted_by2_4_13_port, 
      A_neg_shifted_by2_4_12_port, A_neg_shifted_by2_4_11_port, 
      A_neg_shifted_by2_4_10_port, A_neg_shifted_by2_4_9_port, 
      A_neg_shifted_by2_4_8_port, A_neg_shifted_by2_4_7_port, 
      A_neg_shifted_by2_4_6_port, A_neg_shifted_by2_4_5_port, 
      A_neg_shifted_by2_4_4_port, A_neg_shifted_by2_4_3_port, 
      A_neg_shifted_by2_4_2_port, A_neg_shifted_by2_4_1_port, 
      A_neg_shifted_by2_4_0_port, A_neg_shifted_by2_5_63_port, 
      A_neg_shifted_by2_5_62_port, A_neg_shifted_by2_5_61_port, 
      A_neg_shifted_by2_5_60_port, A_neg_shifted_by2_5_59_port, 
      A_neg_shifted_by2_5_58_port, A_neg_shifted_by2_5_57_port, 
      A_neg_shifted_by2_5_56_port, A_neg_shifted_by2_5_55_port, 
      A_neg_shifted_by2_5_54_port, A_neg_shifted_by2_5_53_port, 
      A_neg_shifted_by2_5_52_port, A_neg_shifted_by2_5_51_port, 
      A_neg_shifted_by2_5_50_port, A_neg_shifted_by2_5_49_port, 
      A_neg_shifted_by2_5_48_port, A_neg_shifted_by2_5_47_port, 
      A_neg_shifted_by2_5_46_port, A_neg_shifted_by2_5_45_port, 
      A_neg_shifted_by2_5_44_port, A_neg_shifted_by2_5_43_port, 
      A_neg_shifted_by2_5_42_port, A_neg_shifted_by2_5_41_port, 
      A_neg_shifted_by2_5_40_port, A_neg_shifted_by2_5_39_port, 
      A_neg_shifted_by2_5_38_port, A_neg_shifted_by2_5_37_port, 
      A_neg_shifted_by2_5_36_port, A_neg_shifted_by2_5_35_port, 
      A_neg_shifted_by2_5_34_port, A_neg_shifted_by2_5_33_port, 
      A_neg_shifted_by2_5_32_port, A_neg_shifted_by2_5_31_port, 
      A_neg_shifted_by2_5_30_port, A_neg_shifted_by2_5_29_port, 
      A_neg_shifted_by2_5_28_port, A_neg_shifted_by2_5_27_port, 
      A_neg_shifted_by2_5_26_port, A_neg_shifted_by2_5_25_port, 
      A_neg_shifted_by2_5_24_port, A_neg_shifted_by2_5_23_port, 
      A_neg_shifted_by2_5_22_port, A_neg_shifted_by2_5_21_port, 
      A_neg_shifted_by2_5_20_port, A_neg_shifted_by2_5_19_port, 
      A_neg_shifted_by2_5_18_port, A_neg_shifted_by2_5_17_port, 
      A_neg_shifted_by2_5_16_port, A_neg_shifted_by2_5_15_port, 
      A_neg_shifted_by2_5_14_port, A_neg_shifted_by2_5_13_port, 
      A_neg_shifted_by2_5_12_port, A_neg_shifted_by2_5_11_port, 
      A_neg_shifted_by2_5_10_port, A_neg_shifted_by2_5_9_port, 
      A_neg_shifted_by2_5_8_port, A_neg_shifted_by2_5_7_port, 
      A_neg_shifted_by2_5_6_port, A_neg_shifted_by2_5_5_port, 
      A_neg_shifted_by2_5_4_port, A_neg_shifted_by2_5_3_port, 
      A_neg_shifted_by2_5_2_port, A_neg_shifted_by2_5_1_port, 
      A_neg_shifted_by2_5_0_port, A_neg_shifted_by2_6_63_port, 
      A_neg_shifted_by2_6_62_port, A_neg_shifted_by2_6_61_port, 
      A_neg_shifted_by2_6_60_port, A_neg_shifted_by2_6_59_port, 
      A_neg_shifted_by2_6_58_port, A_neg_shifted_by2_6_57_port, 
      A_neg_shifted_by2_6_56_port, A_neg_shifted_by2_6_55_port, 
      A_neg_shifted_by2_6_54_port, A_neg_shifted_by2_6_53_port, 
      A_neg_shifted_by2_6_52_port, A_neg_shifted_by2_6_51_port, 
      A_neg_shifted_by2_6_50_port, A_neg_shifted_by2_6_49_port, 
      A_neg_shifted_by2_6_48_port, A_neg_shifted_by2_6_47_port, 
      A_neg_shifted_by2_6_46_port, A_neg_shifted_by2_6_45_port, 
      A_neg_shifted_by2_6_44_port, A_neg_shifted_by2_6_43_port, 
      A_neg_shifted_by2_6_42_port, A_neg_shifted_by2_6_41_port, 
      A_neg_shifted_by2_6_40_port, A_neg_shifted_by2_6_39_port, 
      A_neg_shifted_by2_6_38_port, A_neg_shifted_by2_6_37_port, 
      A_neg_shifted_by2_6_36_port, A_neg_shifted_by2_6_35_port, 
      A_neg_shifted_by2_6_34_port, A_neg_shifted_by2_6_33_port, 
      A_neg_shifted_by2_6_32_port, A_neg_shifted_by2_6_31_port, 
      A_neg_shifted_by2_6_30_port, A_neg_shifted_by2_6_29_port, 
      A_neg_shifted_by2_6_28_port, A_neg_shifted_by2_6_27_port, 
      A_neg_shifted_by2_6_26_port, A_neg_shifted_by2_6_25_port, 
      A_neg_shifted_by2_6_24_port, A_neg_shifted_by2_6_23_port, 
      A_neg_shifted_by2_6_22_port, A_neg_shifted_by2_6_21_port, 
      A_neg_shifted_by2_6_20_port, A_neg_shifted_by2_6_19_port, 
      A_neg_shifted_by2_6_18_port, A_neg_shifted_by2_6_17_port, 
      A_neg_shifted_by2_6_16_port, A_neg_shifted_by2_6_15_port, 
      A_neg_shifted_by2_6_14_port, A_neg_shifted_by2_6_13_port, 
      A_neg_shifted_by2_6_12_port, A_neg_shifted_by2_6_11_port, 
      A_neg_shifted_by2_6_10_port, A_neg_shifted_by2_6_9_port, 
      A_neg_shifted_by2_6_8_port, A_neg_shifted_by2_6_7_port, 
      A_neg_shifted_by2_6_6_port, A_neg_shifted_by2_6_5_port, 
      A_neg_shifted_by2_6_4_port, A_neg_shifted_by2_6_3_port, 
      A_neg_shifted_by2_6_2_port, A_neg_shifted_by2_6_1_port, 
      A_neg_shifted_by2_6_0_port, A_neg_shifted_by2_7_63_port, 
      A_neg_shifted_by2_7_62_port, A_neg_shifted_by2_7_61_port, 
      A_neg_shifted_by2_7_60_port, A_neg_shifted_by2_7_59_port, 
      A_neg_shifted_by2_7_58_port, A_neg_shifted_by2_7_57_port, 
      A_neg_shifted_by2_7_56_port, A_neg_shifted_by2_7_55_port, 
      A_neg_shifted_by2_7_54_port, A_neg_shifted_by2_7_53_port, 
      A_neg_shifted_by2_7_52_port, A_neg_shifted_by2_7_51_port, 
      A_neg_shifted_by2_7_50_port, A_neg_shifted_by2_7_49_port, 
      A_neg_shifted_by2_7_48_port, A_neg_shifted_by2_7_47_port, 
      A_neg_shifted_by2_7_46_port, A_neg_shifted_by2_7_45_port, 
      A_neg_shifted_by2_7_44_port, A_neg_shifted_by2_7_43_port, 
      A_neg_shifted_by2_7_42_port, A_neg_shifted_by2_7_41_port, 
      A_neg_shifted_by2_7_40_port, A_neg_shifted_by2_7_39_port, 
      A_neg_shifted_by2_7_38_port, A_neg_shifted_by2_7_37_port, 
      A_neg_shifted_by2_7_36_port, A_neg_shifted_by2_7_35_port, 
      A_neg_shifted_by2_7_34_port, A_neg_shifted_by2_7_33_port, 
      A_neg_shifted_by2_7_32_port, A_neg_shifted_by2_7_31_port, 
      A_neg_shifted_by2_7_30_port, A_neg_shifted_by2_7_29_port, 
      A_neg_shifted_by2_7_28_port, A_neg_shifted_by2_7_27_port, 
      A_neg_shifted_by2_7_26_port, A_neg_shifted_by2_7_25_port, 
      A_neg_shifted_by2_7_24_port, A_neg_shifted_by2_7_23_port, 
      A_neg_shifted_by2_7_22_port, A_neg_shifted_by2_7_21_port, 
      A_neg_shifted_by2_7_20_port, A_neg_shifted_by2_7_19_port, 
      A_neg_shifted_by2_7_18_port, A_neg_shifted_by2_7_17_port, 
      A_neg_shifted_by2_7_16_port, A_neg_shifted_by2_7_15_port, 
      A_neg_shifted_by2_7_14_port, A_neg_shifted_by2_7_13_port, 
      A_neg_shifted_by2_7_12_port, A_neg_shifted_by2_7_11_port, 
      A_neg_shifted_by2_7_10_port, A_neg_shifted_by2_7_9_port, 
      A_neg_shifted_by2_7_8_port, A_neg_shifted_by2_7_7_port, 
      A_neg_shifted_by2_7_6_port, A_neg_shifted_by2_7_5_port, 
      A_neg_shifted_by2_7_4_port, A_neg_shifted_by2_7_3_port, 
      A_neg_shifted_by2_7_2_port, A_neg_shifted_by2_7_1_port, 
      A_neg_shifted_by2_7_0_port, A_neg_shifted_by1_8_63_port, 
      A_neg_shifted_by1_8_62_port, A_neg_shifted_by1_8_61_port, 
      A_neg_shifted_by1_8_60_port, A_neg_shifted_by1_8_59_port, 
      A_neg_shifted_by1_8_58_port, A_neg_shifted_by1_8_57_port, 
      A_neg_shifted_by1_8_56_port, A_neg_shifted_by1_8_55_port, 
      A_neg_shifted_by1_8_54_port, A_neg_shifted_by1_8_53_port, 
      A_neg_shifted_by1_8_52_port, A_neg_shifted_by1_8_51_port, 
      A_neg_shifted_by1_8_50_port, A_neg_shifted_by1_8_49_port, 
      A_neg_shifted_by1_8_48_port, A_neg_shifted_by1_8_47_port, 
      A_neg_shifted_by1_8_46_port, A_neg_shifted_by1_8_45_port, 
      A_neg_shifted_by1_8_44_port, A_neg_shifted_by1_8_43_port, 
      A_neg_shifted_by1_8_42_port, A_neg_shifted_by1_8_41_port, 
      A_neg_shifted_by1_8_40_port, A_neg_shifted_by1_8_39_port, 
      A_neg_shifted_by1_8_38_port, A_neg_shifted_by1_8_37_port, 
      A_neg_shifted_by1_8_36_port, A_neg_shifted_by1_8_35_port, 
      A_neg_shifted_by1_8_34_port, A_neg_shifted_by1_8_33_port, 
      A_neg_shifted_by1_8_32_port, A_neg_shifted_by1_8_31_port, 
      A_neg_shifted_by1_8_30_port, A_neg_shifted_by1_8_29_port, 
      A_neg_shifted_by1_8_28_port, A_neg_shifted_by1_8_27_port, 
      A_neg_shifted_by1_8_26_port, A_neg_shifted_by1_8_25_port, 
      A_neg_shifted_by1_8_24_port, A_neg_shifted_by1_8_23_port, 
      A_neg_shifted_by1_8_22_port, A_neg_shifted_by1_8_21_port, 
      A_neg_shifted_by1_8_20_port, A_neg_shifted_by1_8_19_port, 
      A_neg_shifted_by1_8_18_port, A_neg_shifted_by1_8_17_port, 
      A_neg_shifted_by1_8_16_port, A_neg_shifted_by1_8_15_port, 
      A_neg_shifted_by1_8_14_port, A_neg_shifted_by1_8_13_port, 
      A_neg_shifted_by1_8_12_port, A_neg_shifted_by1_8_11_port, 
      A_neg_shifted_by1_8_10_port, A_neg_shifted_by1_8_9_port, 
      A_neg_shifted_by1_8_8_port, A_neg_shifted_by1_8_7_port, 
      A_neg_shifted_by1_8_6_port, A_neg_shifted_by1_8_5_port, 
      A_neg_shifted_by1_8_4_port, A_neg_shifted_by1_8_3_port, 
      A_neg_shifted_by1_8_2_port, A_neg_shifted_by1_8_1_port, 
      A_neg_shifted_by1_8_0_port, A_neg_shifted_by1_9_63_port, 
      A_neg_shifted_by1_9_62_port, A_neg_shifted_by1_9_61_port, 
      A_neg_shifted_by1_9_60_port, A_neg_shifted_by1_9_59_port, 
      A_neg_shifted_by1_9_58_port, A_neg_shifted_by1_9_57_port, 
      A_neg_shifted_by1_9_56_port, A_neg_shifted_by1_9_55_port, 
      A_neg_shifted_by1_9_54_port, A_neg_shifted_by1_9_53_port, 
      A_neg_shifted_by1_9_52_port, A_neg_shifted_by1_9_51_port, 
      A_neg_shifted_by1_9_50_port, A_neg_shifted_by1_9_49_port, 
      A_neg_shifted_by1_9_48_port, A_neg_shifted_by1_9_47_port, 
      A_neg_shifted_by1_9_46_port, A_neg_shifted_by1_9_45_port, 
      A_neg_shifted_by1_9_44_port, A_neg_shifted_by1_9_43_port, 
      A_neg_shifted_by1_9_42_port, A_neg_shifted_by1_9_41_port, 
      A_neg_shifted_by1_9_40_port, A_neg_shifted_by1_9_39_port, 
      A_neg_shifted_by1_9_38_port, A_neg_shifted_by1_9_37_port, 
      A_neg_shifted_by1_9_36_port, A_neg_shifted_by1_9_35_port, 
      A_neg_shifted_by1_9_34_port, A_neg_shifted_by1_9_33_port, 
      A_neg_shifted_by1_9_32_port, A_neg_shifted_by1_9_31_port, 
      A_neg_shifted_by1_9_30_port, A_neg_shifted_by1_9_29_port, 
      A_neg_shifted_by1_9_28_port, A_neg_shifted_by1_9_27_port, 
      A_neg_shifted_by1_9_26_port, A_neg_shifted_by1_9_25_port, 
      A_neg_shifted_by1_9_24_port, A_neg_shifted_by1_9_23_port, 
      A_neg_shifted_by1_9_22_port, A_neg_shifted_by1_9_21_port, 
      A_neg_shifted_by1_9_20_port, A_neg_shifted_by1_9_19_port, 
      A_neg_shifted_by1_9_18_port, A_neg_shifted_by1_9_17_port, 
      A_neg_shifted_by1_9_16_port, A_neg_shifted_by1_9_15_port, 
      A_neg_shifted_by1_9_14_port, A_neg_shifted_by1_9_13_port, 
      A_neg_shifted_by1_9_12_port, A_neg_shifted_by1_9_11_port, 
      A_neg_shifted_by1_9_10_port, A_neg_shifted_by1_9_9_port, 
      A_neg_shifted_by1_9_8_port, A_neg_shifted_by1_9_7_port, 
      A_neg_shifted_by1_9_6_port, A_neg_shifted_by1_9_5_port, 
      A_neg_shifted_by1_9_4_port, A_neg_shifted_by1_9_3_port, 
      A_neg_shifted_by1_9_2_port, A_neg_shifted_by1_9_1_port, 
      A_neg_shifted_by1_9_0_port, A_neg_shifted_by1_10_63_port, 
      A_neg_shifted_by1_10_62_port, A_neg_shifted_by1_10_61_port, 
      A_neg_shifted_by1_10_60_port, A_neg_shifted_by1_10_59_port, 
      A_neg_shifted_by1_10_58_port, A_neg_shifted_by1_10_57_port, 
      A_neg_shifted_by1_10_56_port, A_neg_shifted_by1_10_55_port, 
      A_neg_shifted_by1_10_54_port, A_neg_shifted_by1_10_53_port, 
      A_neg_shifted_by1_10_52_port, A_neg_shifted_by1_10_51_port, 
      A_neg_shifted_by1_10_50_port, A_neg_shifted_by1_10_49_port, 
      A_neg_shifted_by1_10_48_port, A_neg_shifted_by1_10_47_port, 
      A_neg_shifted_by1_10_46_port, A_neg_shifted_by1_10_45_port, 
      A_neg_shifted_by1_10_44_port, A_neg_shifted_by1_10_43_port, 
      A_neg_shifted_by1_10_42_port, A_neg_shifted_by1_10_41_port, 
      A_neg_shifted_by1_10_40_port, A_neg_shifted_by1_10_39_port, 
      A_neg_shifted_by1_10_38_port, A_neg_shifted_by1_10_37_port, 
      A_neg_shifted_by1_10_36_port, A_neg_shifted_by1_10_35_port, 
      A_neg_shifted_by1_10_34_port, A_neg_shifted_by1_10_33_port, 
      A_neg_shifted_by1_10_32_port, A_neg_shifted_by1_10_31_port, 
      A_neg_shifted_by1_10_30_port, A_neg_shifted_by1_10_29_port, 
      A_neg_shifted_by1_10_28_port, A_neg_shifted_by1_10_27_port, 
      A_neg_shifted_by1_10_26_port, A_neg_shifted_by1_10_25_port, 
      A_neg_shifted_by1_10_24_port, A_neg_shifted_by1_10_23_port, 
      A_neg_shifted_by1_10_22_port, A_neg_shifted_by1_10_21_port, 
      A_neg_shifted_by1_10_20_port, A_neg_shifted_by1_10_19_port, 
      A_neg_shifted_by1_10_18_port, A_neg_shifted_by1_10_17_port, 
      A_neg_shifted_by1_10_16_port, A_neg_shifted_by1_10_15_port, 
      A_neg_shifted_by1_10_14_port, A_neg_shifted_by1_10_13_port, 
      A_neg_shifted_by1_10_12_port, A_neg_shifted_by1_10_11_port, 
      A_neg_shifted_by1_10_10_port, A_neg_shifted_by1_10_9_port, 
      A_neg_shifted_by1_10_8_port, A_neg_shifted_by1_10_7_port, 
      A_neg_shifted_by1_10_6_port, A_neg_shifted_by1_10_5_port, 
      A_neg_shifted_by1_10_4_port, A_neg_shifted_by1_10_3_port, 
      A_neg_shifted_by1_10_2_port, A_neg_shifted_by1_10_1_port, 
      A_neg_shifted_by1_10_0_port, A_neg_shifted_by1_11_63_port, 
      A_neg_shifted_by1_11_62_port, A_neg_shifted_by1_11_61_port, 
      A_neg_shifted_by1_11_60_port, A_neg_shifted_by1_11_59_port, 
      A_neg_shifted_by1_11_58_port, A_neg_shifted_by1_11_57_port, 
      A_neg_shifted_by1_11_56_port, A_neg_shifted_by1_11_55_port, 
      A_neg_shifted_by1_11_54_port, A_neg_shifted_by1_11_53_port, 
      A_neg_shifted_by1_11_52_port, A_neg_shifted_by1_11_51_port, 
      A_neg_shifted_by1_11_50_port, A_neg_shifted_by1_11_49_port, 
      A_neg_shifted_by1_11_48_port, A_neg_shifted_by1_11_47_port, 
      A_neg_shifted_by1_11_46_port, A_neg_shifted_by1_11_45_port, 
      A_neg_shifted_by1_11_44_port, A_neg_shifted_by1_11_43_port, 
      A_neg_shifted_by1_11_42_port, A_neg_shifted_by1_11_41_port, 
      A_neg_shifted_by1_11_40_port, A_neg_shifted_by1_11_39_port, 
      A_neg_shifted_by1_11_38_port, A_neg_shifted_by1_11_37_port, 
      A_neg_shifted_by1_11_36_port, A_neg_shifted_by1_11_35_port, 
      A_neg_shifted_by1_11_34_port, A_neg_shifted_by1_11_33_port, 
      A_neg_shifted_by1_11_32_port, A_neg_shifted_by1_11_31_port, 
      A_neg_shifted_by1_11_30_port, A_neg_shifted_by1_11_29_port, 
      A_neg_shifted_by1_11_28_port, A_neg_shifted_by1_11_27_port, 
      A_neg_shifted_by1_11_26_port, A_neg_shifted_by1_11_25_port, 
      A_neg_shifted_by1_11_24_port, A_neg_shifted_by1_11_23_port, 
      A_neg_shifted_by1_11_22_port, A_neg_shifted_by1_11_21_port, 
      A_neg_shifted_by1_11_20_port, A_neg_shifted_by1_11_19_port, 
      A_neg_shifted_by1_11_18_port, A_neg_shifted_by1_11_17_port, 
      A_neg_shifted_by1_11_16_port, A_neg_shifted_by1_11_15_port, 
      A_neg_shifted_by1_11_14_port, A_neg_shifted_by1_11_13_port, 
      A_neg_shifted_by1_11_12_port, A_neg_shifted_by1_11_11_port, 
      A_neg_shifted_by1_11_10_port, A_neg_shifted_by1_11_9_port, 
      A_neg_shifted_by1_11_8_port, A_neg_shifted_by1_11_7_port, 
      A_neg_shifted_by1_11_6_port, A_neg_shifted_by1_11_5_port, 
      A_neg_shifted_by1_11_4_port, A_neg_shifted_by1_11_3_port, 
      A_neg_shifted_by1_11_2_port, A_neg_shifted_by1_11_1_port, 
      A_neg_shifted_by1_11_0_port, A_neg_shifted_by1_12_63_port, 
      A_neg_shifted_by1_12_62_port, A_neg_shifted_by1_12_61_port, 
      A_neg_shifted_by1_12_60_port, A_neg_shifted_by1_12_59_port, 
      A_neg_shifted_by1_12_58_port, A_neg_shifted_by1_12_57_port, 
      A_neg_shifted_by1_12_56_port, A_neg_shifted_by1_12_55_port, 
      A_neg_shifted_by1_12_54_port, A_neg_shifted_by1_12_53_port, 
      A_neg_shifted_by1_12_52_port, A_neg_shifted_by1_12_51_port, 
      A_neg_shifted_by1_12_50_port, A_neg_shifted_by1_12_49_port, 
      A_neg_shifted_by1_12_48_port, A_neg_shifted_by1_12_47_port, 
      A_neg_shifted_by1_12_46_port, A_neg_shifted_by1_12_45_port, 
      A_neg_shifted_by1_12_44_port, A_neg_shifted_by1_12_43_port, 
      A_neg_shifted_by1_12_42_port, A_neg_shifted_by1_12_41_port, 
      A_neg_shifted_by1_12_40_port, A_neg_shifted_by1_12_39_port, 
      A_neg_shifted_by1_12_38_port, A_neg_shifted_by1_12_37_port, 
      A_neg_shifted_by1_12_36_port, A_neg_shifted_by1_12_35_port, 
      A_neg_shifted_by1_12_34_port, A_neg_shifted_by1_12_33_port, 
      A_neg_shifted_by1_12_32_port, A_neg_shifted_by1_12_31_port, 
      A_neg_shifted_by1_12_30_port, A_neg_shifted_by1_12_29_port, 
      A_neg_shifted_by1_12_28_port, A_neg_shifted_by1_12_27_port, 
      A_neg_shifted_by1_12_26_port, A_neg_shifted_by1_12_25_port, 
      A_neg_shifted_by1_12_24_port, A_neg_shifted_by1_12_23_port, 
      A_neg_shifted_by1_12_22_port, A_neg_shifted_by1_12_21_port, 
      A_neg_shifted_by1_12_20_port, A_neg_shifted_by1_12_19_port, 
      A_neg_shifted_by1_12_18_port, A_neg_shifted_by1_12_17_port, 
      A_neg_shifted_by1_12_16_port, A_neg_shifted_by1_12_15_port, 
      A_neg_shifted_by1_12_14_port, A_neg_shifted_by1_12_13_port, 
      A_neg_shifted_by1_12_12_port, A_neg_shifted_by1_12_11_port, 
      A_neg_shifted_by1_12_10_port, A_neg_shifted_by1_12_9_port, 
      A_neg_shifted_by1_12_8_port, A_neg_shifted_by1_12_7_port, 
      A_neg_shifted_by1_12_6_port, A_neg_shifted_by1_12_5_port, 
      A_neg_shifted_by1_12_4_port, A_neg_shifted_by1_12_3_port, 
      A_neg_shifted_by1_12_2_port, A_neg_shifted_by1_12_1_port, 
      A_neg_shifted_by1_12_0_port, A_neg_shifted_by1_13_63_port, 
      A_neg_shifted_by1_13_62_port, A_neg_shifted_by1_13_61_port, 
      A_neg_shifted_by1_13_60_port, A_neg_shifted_by1_13_59_port, 
      A_neg_shifted_by1_13_58_port, A_neg_shifted_by1_13_57_port, 
      A_neg_shifted_by1_13_56_port, A_neg_shifted_by1_13_55_port, 
      A_neg_shifted_by1_13_54_port, A_neg_shifted_by1_13_53_port, 
      A_neg_shifted_by1_13_52_port, A_neg_shifted_by1_13_51_port, 
      A_neg_shifted_by1_13_50_port, A_neg_shifted_by1_13_49_port, 
      A_neg_shifted_by1_13_48_port, A_neg_shifted_by1_13_47_port, 
      A_neg_shifted_by1_13_46_port, A_neg_shifted_by1_13_45_port, 
      A_neg_shifted_by1_13_44_port, A_neg_shifted_by1_13_43_port, 
      A_neg_shifted_by1_13_42_port, A_neg_shifted_by1_13_41_port, 
      A_neg_shifted_by1_13_40_port, A_neg_shifted_by1_13_39_port, 
      A_neg_shifted_by1_13_38_port, A_neg_shifted_by1_13_37_port, 
      A_neg_shifted_by1_13_36_port, A_neg_shifted_by1_13_35_port, 
      A_neg_shifted_by1_13_34_port, A_neg_shifted_by1_13_33_port, 
      A_neg_shifted_by1_13_32_port, A_neg_shifted_by1_13_31_port, 
      A_neg_shifted_by1_13_30_port, A_neg_shifted_by1_13_29_port, 
      A_neg_shifted_by1_13_28_port, A_neg_shifted_by1_13_27_port, 
      A_neg_shifted_by1_13_26_port, A_neg_shifted_by1_13_25_port, 
      A_neg_shifted_by1_13_24_port, A_neg_shifted_by1_13_23_port, 
      A_neg_shifted_by1_13_22_port, A_neg_shifted_by1_13_21_port, 
      A_neg_shifted_by1_13_20_port, A_neg_shifted_by1_13_19_port, 
      A_neg_shifted_by1_13_18_port, A_neg_shifted_by1_13_17_port, 
      A_neg_shifted_by1_13_16_port, A_neg_shifted_by1_13_15_port, 
      A_neg_shifted_by1_13_14_port, A_neg_shifted_by1_13_13_port, 
      A_neg_shifted_by1_13_12_port, A_neg_shifted_by1_13_11_port, 
      A_neg_shifted_by1_13_10_port, A_neg_shifted_by1_13_9_port, 
      A_neg_shifted_by1_13_8_port, A_neg_shifted_by1_13_7_port, 
      A_neg_shifted_by1_13_6_port, A_neg_shifted_by1_13_5_port, 
      A_neg_shifted_by1_13_4_port, A_neg_shifted_by1_13_3_port, 
      A_neg_shifted_by1_13_2_port, A_neg_shifted_by1_13_1_port, 
      A_neg_shifted_by1_13_0_port, A_neg_shifted_by1_14_63_port, 
      A_neg_shifted_by1_14_62_port, A_neg_shifted_by1_14_61_port, 
      A_neg_shifted_by1_14_60_port, A_neg_shifted_by1_14_59_port, 
      A_neg_shifted_by1_14_58_port, A_neg_shifted_by1_14_57_port, 
      A_neg_shifted_by1_14_56_port, A_neg_shifted_by1_14_55_port, 
      A_neg_shifted_by1_14_54_port, A_neg_shifted_by1_14_53_port, 
      A_neg_shifted_by1_14_52_port, A_neg_shifted_by1_14_51_port, 
      A_neg_shifted_by1_14_50_port, A_neg_shifted_by1_14_49_port, 
      A_neg_shifted_by1_14_48_port, A_neg_shifted_by1_14_47_port, 
      A_neg_shifted_by1_14_46_port, A_neg_shifted_by1_14_45_port, 
      A_neg_shifted_by1_14_44_port, A_neg_shifted_by1_14_43_port, 
      A_neg_shifted_by1_14_42_port, A_neg_shifted_by1_14_41_port, 
      A_neg_shifted_by1_14_40_port, A_neg_shifted_by1_14_39_port, 
      A_neg_shifted_by1_14_38_port, A_neg_shifted_by1_14_37_port, 
      A_neg_shifted_by1_14_36_port, A_neg_shifted_by1_14_35_port, 
      A_neg_shifted_by1_14_34_port, A_neg_shifted_by1_14_33_port, 
      A_neg_shifted_by1_14_32_port, A_neg_shifted_by1_14_31_port, 
      A_neg_shifted_by1_14_30_port, A_neg_shifted_by1_14_29_port, 
      A_neg_shifted_by1_14_28_port, A_neg_shifted_by1_14_27_port, 
      A_neg_shifted_by1_14_26_port, A_neg_shifted_by1_14_25_port, 
      A_neg_shifted_by1_14_24_port, A_neg_shifted_by1_14_23_port, 
      A_neg_shifted_by1_14_22_port, A_neg_shifted_by1_14_21_port, 
      A_neg_shifted_by1_14_20_port, A_neg_shifted_by1_14_19_port, 
      A_neg_shifted_by1_14_18_port, A_neg_shifted_by1_14_17_port, 
      A_neg_shifted_by1_14_16_port, A_neg_shifted_by1_14_15_port, 
      A_neg_shifted_by1_14_14_port, A_neg_shifted_by1_14_13_port, 
      A_neg_shifted_by1_14_12_port, A_neg_shifted_by1_14_11_port, 
      A_neg_shifted_by1_14_10_port, A_neg_shifted_by1_14_9_port, 
      A_neg_shifted_by1_14_8_port, A_neg_shifted_by1_14_7_port, 
      A_neg_shifted_by1_14_6_port, A_neg_shifted_by1_14_5_port, 
      A_neg_shifted_by1_14_4_port, A_neg_shifted_by1_14_3_port, 
      A_neg_shifted_by1_14_2_port, A_neg_shifted_by1_14_1_port, 
      A_neg_shifted_by1_14_0_port, A_neg_shifted_by1_15_63_port, 
      A_neg_shifted_by1_15_62_port, A_neg_shifted_by1_15_61_port, 
      A_neg_shifted_by1_15_60_port, A_neg_shifted_by1_15_59_port, 
      A_neg_shifted_by1_15_58_port, A_neg_shifted_by1_15_57_port, 
      A_neg_shifted_by1_15_56_port, A_neg_shifted_by1_15_55_port, 
      A_neg_shifted_by1_15_54_port, A_neg_shifted_by1_15_53_port, 
      A_neg_shifted_by1_15_52_port, A_neg_shifted_by1_15_51_port, 
      A_neg_shifted_by1_15_50_port, A_neg_shifted_by1_15_49_port, 
      A_neg_shifted_by1_15_48_port, A_neg_shifted_by1_15_47_port, 
      A_neg_shifted_by1_15_46_port, A_neg_shifted_by1_15_45_port, 
      A_neg_shifted_by1_15_44_port, A_neg_shifted_by1_15_43_port, 
      A_neg_shifted_by1_15_42_port, A_neg_shifted_by1_15_41_port, 
      A_neg_shifted_by1_15_40_port, A_neg_shifted_by1_15_39_port, 
      A_neg_shifted_by1_15_38_port, A_neg_shifted_by1_15_37_port, 
      A_neg_shifted_by1_15_36_port, A_neg_shifted_by1_15_35_port, 
      A_neg_shifted_by1_15_34_port, A_neg_shifted_by1_15_33_port, 
      A_neg_shifted_by1_15_32_port, A_neg_shifted_by1_15_31_port, 
      A_neg_shifted_by1_15_30_port, A_neg_shifted_by1_15_29_port, 
      A_neg_shifted_by1_15_28_port, A_neg_shifted_by1_15_27_port, 
      A_neg_shifted_by1_15_26_port, A_neg_shifted_by1_15_25_port, 
      A_neg_shifted_by1_15_24_port, A_neg_shifted_by1_15_23_port, 
      A_neg_shifted_by1_15_22_port, A_neg_shifted_by1_15_21_port, 
      A_neg_shifted_by1_15_20_port, A_neg_shifted_by1_15_19_port, 
      A_neg_shifted_by1_15_18_port, A_neg_shifted_by1_15_17_port, 
      A_neg_shifted_by1_15_16_port, A_neg_shifted_by1_15_15_port, 
      A_neg_shifted_by1_15_14_port, A_neg_shifted_by1_15_13_port, 
      A_neg_shifted_by1_15_12_port, A_neg_shifted_by1_15_11_port, 
      A_neg_shifted_by1_15_10_port, A_neg_shifted_by1_15_9_port, 
      A_neg_shifted_by1_15_8_port, A_neg_shifted_by1_15_7_port, 
      A_neg_shifted_by1_15_6_port, A_neg_shifted_by1_15_5_port, 
      A_neg_shifted_by1_15_4_port, A_neg_shifted_by1_15_3_port, 
      A_neg_shifted_by1_15_2_port, A_neg_shifted_by1_15_1_port, 
      A_neg_shifted_by1_15_0_port, A_neg_shifted_by2_8_63_port, 
      A_neg_shifted_by2_8_62_port, A_neg_shifted_by2_8_61_port, 
      A_neg_shifted_by2_8_60_port, A_neg_shifted_by2_8_59_port, 
      A_neg_shifted_by2_8_58_port, A_neg_shifted_by2_8_57_port, 
      A_neg_shifted_by2_8_56_port, A_neg_shifted_by2_8_55_port, 
      A_neg_shifted_by2_8_54_port, A_neg_shifted_by2_8_53_port, 
      A_neg_shifted_by2_8_52_port, A_neg_shifted_by2_8_51_port, 
      A_neg_shifted_by2_8_50_port, A_neg_shifted_by2_8_49_port, 
      A_neg_shifted_by2_8_48_port, A_neg_shifted_by2_8_47_port, 
      A_neg_shifted_by2_8_46_port, A_neg_shifted_by2_8_45_port, 
      A_neg_shifted_by2_8_44_port, A_neg_shifted_by2_8_43_port, 
      A_neg_shifted_by2_8_42_port, A_neg_shifted_by2_8_41_port, 
      A_neg_shifted_by2_8_40_port, A_neg_shifted_by2_8_39_port, 
      A_neg_shifted_by2_8_38_port, A_neg_shifted_by2_8_37_port, 
      A_neg_shifted_by2_8_36_port, A_neg_shifted_by2_8_35_port, 
      A_neg_shifted_by2_8_34_port, A_neg_shifted_by2_8_33_port, 
      A_neg_shifted_by2_8_32_port, A_neg_shifted_by2_8_31_port, 
      A_neg_shifted_by2_8_30_port, A_neg_shifted_by2_8_29_port, 
      A_neg_shifted_by2_8_28_port, A_neg_shifted_by2_8_27_port, 
      A_neg_shifted_by2_8_26_port, A_neg_shifted_by2_8_25_port, 
      A_neg_shifted_by2_8_24_port, A_neg_shifted_by2_8_23_port, 
      A_neg_shifted_by2_8_22_port, A_neg_shifted_by2_8_21_port, 
      A_neg_shifted_by2_8_20_port, A_neg_shifted_by2_8_19_port, 
      A_neg_shifted_by2_8_18_port, A_neg_shifted_by2_8_17_port, 
      A_neg_shifted_by2_8_16_port, A_neg_shifted_by2_8_15_port, 
      A_neg_shifted_by2_8_14_port, A_neg_shifted_by2_8_13_port, 
      A_neg_shifted_by2_8_12_port, A_neg_shifted_by2_8_11_port, 
      A_neg_shifted_by2_8_10_port, A_neg_shifted_by2_8_9_port, 
      A_neg_shifted_by2_8_8_port, A_neg_shifted_by2_8_7_port, 
      A_neg_shifted_by2_8_6_port, A_neg_shifted_by2_8_5_port, 
      A_neg_shifted_by2_8_4_port, A_neg_shifted_by2_8_3_port, 
      A_neg_shifted_by2_8_2_port, A_neg_shifted_by2_8_1_port, 
      A_neg_shifted_by2_8_0_port, A_neg_shifted_by2_9_63_port, 
      A_neg_shifted_by2_9_62_port, A_neg_shifted_by2_9_61_port, 
      A_neg_shifted_by2_9_60_port, A_neg_shifted_by2_9_59_port, 
      A_neg_shifted_by2_9_58_port, A_neg_shifted_by2_9_57_port, 
      A_neg_shifted_by2_9_56_port, A_neg_shifted_by2_9_55_port, 
      A_neg_shifted_by2_9_54_port, A_neg_shifted_by2_9_53_port, 
      A_neg_shifted_by2_9_52_port, A_neg_shifted_by2_9_51_port, 
      A_neg_shifted_by2_9_50_port, A_neg_shifted_by2_9_49_port, 
      A_neg_shifted_by2_9_48_port, A_neg_shifted_by2_9_47_port, 
      A_neg_shifted_by2_9_46_port, A_neg_shifted_by2_9_45_port, 
      A_neg_shifted_by2_9_44_port, A_neg_shifted_by2_9_43_port, 
      A_neg_shifted_by2_9_42_port, A_neg_shifted_by2_9_41_port, 
      A_neg_shifted_by2_9_40_port, A_neg_shifted_by2_9_39_port, 
      A_neg_shifted_by2_9_38_port, A_neg_shifted_by2_9_37_port, 
      A_neg_shifted_by2_9_36_port, A_neg_shifted_by2_9_35_port, 
      A_neg_shifted_by2_9_34_port, A_neg_shifted_by2_9_33_port, 
      A_neg_shifted_by2_9_32_port, A_neg_shifted_by2_9_31_port, 
      A_neg_shifted_by2_9_30_port, A_neg_shifted_by2_9_29_port, 
      A_neg_shifted_by2_9_28_port, A_neg_shifted_by2_9_27_port, 
      A_neg_shifted_by2_9_26_port, A_neg_shifted_by2_9_25_port, 
      A_neg_shifted_by2_9_24_port, A_neg_shifted_by2_9_23_port, 
      A_neg_shifted_by2_9_22_port, A_neg_shifted_by2_9_21_port, 
      A_neg_shifted_by2_9_20_port, A_neg_shifted_by2_9_19_port, 
      A_neg_shifted_by2_9_18_port, A_neg_shifted_by2_9_17_port, 
      A_neg_shifted_by2_9_16_port, A_neg_shifted_by2_9_15_port, 
      A_neg_shifted_by2_9_14_port, A_neg_shifted_by2_9_13_port, 
      A_neg_shifted_by2_9_12_port, A_neg_shifted_by2_9_11_port, 
      A_neg_shifted_by2_9_10_port, A_neg_shifted_by2_9_9_port, 
      A_neg_shifted_by2_9_8_port, A_neg_shifted_by2_9_7_port, 
      A_neg_shifted_by2_9_6_port, A_neg_shifted_by2_9_5_port, 
      A_neg_shifted_by2_9_4_port, A_neg_shifted_by2_9_3_port, 
      A_neg_shifted_by2_9_2_port, A_neg_shifted_by2_9_1_port, 
      A_neg_shifted_by2_9_0_port, A_neg_shifted_by2_10_63_port, 
      A_neg_shifted_by2_10_62_port, A_neg_shifted_by2_10_61_port, 
      A_neg_shifted_by2_10_60_port, A_neg_shifted_by2_10_59_port, 
      A_neg_shifted_by2_10_58_port, A_neg_shifted_by2_10_57_port, 
      A_neg_shifted_by2_10_56_port, A_neg_shifted_by2_10_55_port, 
      A_neg_shifted_by2_10_54_port, A_neg_shifted_by2_10_53_port, 
      A_neg_shifted_by2_10_52_port, A_neg_shifted_by2_10_51_port, 
      A_neg_shifted_by2_10_50_port, A_neg_shifted_by2_10_49_port, 
      A_neg_shifted_by2_10_48_port, A_neg_shifted_by2_10_47_port, 
      A_neg_shifted_by2_10_46_port, A_neg_shifted_by2_10_45_port, 
      A_neg_shifted_by2_10_44_port, A_neg_shifted_by2_10_43_port, 
      A_neg_shifted_by2_10_42_port, A_neg_shifted_by2_10_41_port, 
      A_neg_shifted_by2_10_40_port, A_neg_shifted_by2_10_39_port, 
      A_neg_shifted_by2_10_38_port, A_neg_shifted_by2_10_37_port, 
      A_neg_shifted_by2_10_36_port, A_neg_shifted_by2_10_35_port, 
      A_neg_shifted_by2_10_34_port, A_neg_shifted_by2_10_33_port, 
      A_neg_shifted_by2_10_32_port, A_neg_shifted_by2_10_31_port, 
      A_neg_shifted_by2_10_30_port, A_neg_shifted_by2_10_29_port, 
      A_neg_shifted_by2_10_28_port, A_neg_shifted_by2_10_27_port, 
      A_neg_shifted_by2_10_26_port, A_neg_shifted_by2_10_25_port, 
      A_neg_shifted_by2_10_24_port, A_neg_shifted_by2_10_23_port, 
      A_neg_shifted_by2_10_22_port, A_neg_shifted_by2_10_21_port, 
      A_neg_shifted_by2_10_20_port, A_neg_shifted_by2_10_19_port, 
      A_neg_shifted_by2_10_18_port, A_neg_shifted_by2_10_17_port, 
      A_neg_shifted_by2_10_16_port, A_neg_shifted_by2_10_15_port, 
      A_neg_shifted_by2_10_14_port, A_neg_shifted_by2_10_13_port, 
      A_neg_shifted_by2_10_12_port, A_neg_shifted_by2_10_11_port, 
      A_neg_shifted_by2_10_10_port, A_neg_shifted_by2_10_9_port, 
      A_neg_shifted_by2_10_8_port, A_neg_shifted_by2_10_7_port, 
      A_neg_shifted_by2_10_6_port, A_neg_shifted_by2_10_5_port, 
      A_neg_shifted_by2_10_4_port, A_neg_shifted_by2_10_3_port, 
      A_neg_shifted_by2_10_2_port, A_neg_shifted_by2_10_1_port, 
      A_neg_shifted_by2_10_0_port, A_neg_shifted_by2_11_63_port, 
      A_neg_shifted_by2_11_62_port, A_neg_shifted_by2_11_61_port, 
      A_neg_shifted_by2_11_60_port, A_neg_shifted_by2_11_59_port, 
      A_neg_shifted_by2_11_58_port, A_neg_shifted_by2_11_57_port, 
      A_neg_shifted_by2_11_56_port, A_neg_shifted_by2_11_55_port, 
      A_neg_shifted_by2_11_54_port, A_neg_shifted_by2_11_53_port, 
      A_neg_shifted_by2_11_52_port, A_neg_shifted_by2_11_51_port, 
      A_neg_shifted_by2_11_50_port, A_neg_shifted_by2_11_49_port, 
      A_neg_shifted_by2_11_48_port, A_neg_shifted_by2_11_47_port, 
      A_neg_shifted_by2_11_46_port, A_neg_shifted_by2_11_45_port, 
      A_neg_shifted_by2_11_44_port, A_neg_shifted_by2_11_43_port, 
      A_neg_shifted_by2_11_42_port, A_neg_shifted_by2_11_41_port, 
      A_neg_shifted_by2_11_40_port, A_neg_shifted_by2_11_39_port, 
      A_neg_shifted_by2_11_38_port, A_neg_shifted_by2_11_37_port, 
      A_neg_shifted_by2_11_36_port, A_neg_shifted_by2_11_35_port, 
      A_neg_shifted_by2_11_34_port, A_neg_shifted_by2_11_33_port, 
      A_neg_shifted_by2_11_32_port, A_neg_shifted_by2_11_31_port, 
      A_neg_shifted_by2_11_30_port, A_neg_shifted_by2_11_29_port, 
      A_neg_shifted_by2_11_28_port, A_neg_shifted_by2_11_27_port, 
      A_neg_shifted_by2_11_26_port, A_neg_shifted_by2_11_25_port, 
      A_neg_shifted_by2_11_24_port, A_neg_shifted_by2_11_23_port, 
      A_neg_shifted_by2_11_22_port, A_neg_shifted_by2_11_21_port, 
      A_neg_shifted_by2_11_20_port, A_neg_shifted_by2_11_19_port, 
      A_neg_shifted_by2_11_18_port, A_neg_shifted_by2_11_17_port, 
      A_neg_shifted_by2_11_16_port, A_neg_shifted_by2_11_15_port, 
      A_neg_shifted_by2_11_14_port, A_neg_shifted_by2_11_13_port, 
      A_neg_shifted_by2_11_12_port, A_neg_shifted_by2_11_11_port, 
      A_neg_shifted_by2_11_10_port, A_neg_shifted_by2_11_9_port, 
      A_neg_shifted_by2_11_8_port, A_neg_shifted_by2_11_7_port, 
      A_neg_shifted_by2_11_6_port, A_neg_shifted_by2_11_5_port, 
      A_neg_shifted_by2_11_4_port, A_neg_shifted_by2_11_3_port, 
      A_neg_shifted_by2_11_2_port, A_neg_shifted_by2_11_1_port, 
      A_neg_shifted_by2_11_0_port, A_neg_shifted_by2_12_63_port, 
      A_neg_shifted_by2_12_62_port, A_neg_shifted_by2_12_61_port, 
      A_neg_shifted_by2_12_60_port, A_neg_shifted_by2_12_59_port, 
      A_neg_shifted_by2_12_58_port, A_neg_shifted_by2_12_57_port, 
      A_neg_shifted_by2_12_56_port, A_neg_shifted_by2_12_55_port, 
      A_neg_shifted_by2_12_54_port, A_neg_shifted_by2_12_53_port, 
      A_neg_shifted_by2_12_52_port, A_neg_shifted_by2_12_51_port, 
      A_neg_shifted_by2_12_50_port, A_neg_shifted_by2_12_49_port, 
      A_neg_shifted_by2_12_48_port, A_neg_shifted_by2_12_47_port, 
      A_neg_shifted_by2_12_46_port, A_neg_shifted_by2_12_45_port, 
      A_neg_shifted_by2_12_44_port, A_neg_shifted_by2_12_43_port, 
      A_neg_shifted_by2_12_42_port, A_neg_shifted_by2_12_41_port, 
      A_neg_shifted_by2_12_40_port, A_neg_shifted_by2_12_39_port, 
      A_neg_shifted_by2_12_38_port, A_neg_shifted_by2_12_37_port, 
      A_neg_shifted_by2_12_36_port, A_neg_shifted_by2_12_35_port, 
      A_neg_shifted_by2_12_34_port, A_neg_shifted_by2_12_33_port, 
      A_neg_shifted_by2_12_32_port, A_neg_shifted_by2_12_31_port, 
      A_neg_shifted_by2_12_30_port, A_neg_shifted_by2_12_29_port, 
      A_neg_shifted_by2_12_28_port, A_neg_shifted_by2_12_27_port, 
      A_neg_shifted_by2_12_26_port, A_neg_shifted_by2_12_25_port, 
      A_neg_shifted_by2_12_24_port, A_neg_shifted_by2_12_23_port, 
      A_neg_shifted_by2_12_22_port, A_neg_shifted_by2_12_21_port, 
      A_neg_shifted_by2_12_20_port, A_neg_shifted_by2_12_19_port, 
      A_neg_shifted_by2_12_18_port, A_neg_shifted_by2_12_17_port, 
      A_neg_shifted_by2_12_16_port, A_neg_shifted_by2_12_15_port, 
      A_neg_shifted_by2_12_14_port, A_neg_shifted_by2_12_13_port, 
      A_neg_shifted_by2_12_12_port, A_neg_shifted_by2_12_11_port, 
      A_neg_shifted_by2_12_10_port, A_neg_shifted_by2_12_9_port, 
      A_neg_shifted_by2_12_8_port, A_neg_shifted_by2_12_7_port, 
      A_neg_shifted_by2_12_6_port, A_neg_shifted_by2_12_5_port, 
      A_neg_shifted_by2_12_4_port, A_neg_shifted_by2_12_3_port, 
      A_neg_shifted_by2_12_2_port, A_neg_shifted_by2_12_1_port, 
      A_neg_shifted_by2_12_0_port, A_neg_shifted_by2_13_63_port, 
      A_neg_shifted_by2_13_62_port, A_neg_shifted_by2_13_61_port, 
      A_neg_shifted_by2_13_60_port, A_neg_shifted_by2_13_59_port, 
      A_neg_shifted_by2_13_58_port, A_neg_shifted_by2_13_57_port, 
      A_neg_shifted_by2_13_56_port, A_neg_shifted_by2_13_55_port, 
      A_neg_shifted_by2_13_54_port, A_neg_shifted_by2_13_53_port, 
      A_neg_shifted_by2_13_52_port, A_neg_shifted_by2_13_51_port, 
      A_neg_shifted_by2_13_50_port, A_neg_shifted_by2_13_49_port, 
      A_neg_shifted_by2_13_48_port, A_neg_shifted_by2_13_47_port, 
      A_neg_shifted_by2_13_46_port, A_neg_shifted_by2_13_45_port, 
      A_neg_shifted_by2_13_44_port, A_neg_shifted_by2_13_43_port, 
      A_neg_shifted_by2_13_42_port, A_neg_shifted_by2_13_41_port, 
      A_neg_shifted_by2_13_40_port, A_neg_shifted_by2_13_39_port, 
      A_neg_shifted_by2_13_38_port, A_neg_shifted_by2_13_37_port, 
      A_neg_shifted_by2_13_36_port, A_neg_shifted_by2_13_35_port, 
      A_neg_shifted_by2_13_34_port, A_neg_shifted_by2_13_33_port, 
      A_neg_shifted_by2_13_32_port, A_neg_shifted_by2_13_31_port, 
      A_neg_shifted_by2_13_30_port, A_neg_shifted_by2_13_29_port, 
      A_neg_shifted_by2_13_28_port, A_neg_shifted_by2_13_27_port, 
      A_neg_shifted_by2_13_26_port, A_neg_shifted_by2_13_25_port, 
      A_neg_shifted_by2_13_24_port, A_neg_shifted_by2_13_23_port, 
      A_neg_shifted_by2_13_22_port, A_neg_shifted_by2_13_21_port, 
      A_neg_shifted_by2_13_20_port, A_neg_shifted_by2_13_19_port, 
      A_neg_shifted_by2_13_18_port, A_neg_shifted_by2_13_17_port, 
      A_neg_shifted_by2_13_16_port, A_neg_shifted_by2_13_15_port, 
      A_neg_shifted_by2_13_14_port, A_neg_shifted_by2_13_13_port, 
      A_neg_shifted_by2_13_12_port, A_neg_shifted_by2_13_11_port, 
      A_neg_shifted_by2_13_10_port, A_neg_shifted_by2_13_9_port, 
      A_neg_shifted_by2_13_8_port, A_neg_shifted_by2_13_7_port, 
      A_neg_shifted_by2_13_6_port, A_neg_shifted_by2_13_5_port, 
      A_neg_shifted_by2_13_4_port, A_neg_shifted_by2_13_3_port, 
      A_neg_shifted_by2_13_2_port, A_neg_shifted_by2_13_1_port, 
      A_neg_shifted_by2_13_0_port, A_neg_shifted_by2_14_63_port, 
      A_neg_shifted_by2_14_62_port, A_neg_shifted_by2_14_61_port, 
      A_neg_shifted_by2_14_60_port, A_neg_shifted_by2_14_59_port, 
      A_neg_shifted_by2_14_58_port, A_neg_shifted_by2_14_57_port, 
      A_neg_shifted_by2_14_56_port, A_neg_shifted_by2_14_55_port, 
      A_neg_shifted_by2_14_54_port, A_neg_shifted_by2_14_53_port, 
      A_neg_shifted_by2_14_52_port, A_neg_shifted_by2_14_51_port, 
      A_neg_shifted_by2_14_50_port, A_neg_shifted_by2_14_49_port, 
      A_neg_shifted_by2_14_48_port, A_neg_shifted_by2_14_47_port, 
      A_neg_shifted_by2_14_46_port, A_neg_shifted_by2_14_45_port, 
      A_neg_shifted_by2_14_44_port, A_neg_shifted_by2_14_43_port, 
      A_neg_shifted_by2_14_42_port, A_neg_shifted_by2_14_41_port, 
      A_neg_shifted_by2_14_40_port, A_neg_shifted_by2_14_39_port, 
      A_neg_shifted_by2_14_38_port, A_neg_shifted_by2_14_37_port, 
      A_neg_shifted_by2_14_36_port, A_neg_shifted_by2_14_35_port, 
      A_neg_shifted_by2_14_34_port, A_neg_shifted_by2_14_33_port, 
      A_neg_shifted_by2_14_32_port, A_neg_shifted_by2_14_31_port, 
      A_neg_shifted_by2_14_30_port, A_neg_shifted_by2_14_29_port, 
      A_neg_shifted_by2_14_28_port, A_neg_shifted_by2_14_27_port, 
      A_neg_shifted_by2_14_26_port, A_neg_shifted_by2_14_25_port, 
      A_neg_shifted_by2_14_24_port, A_neg_shifted_by2_14_23_port, 
      A_neg_shifted_by2_14_22_port, A_neg_shifted_by2_14_21_port, 
      A_neg_shifted_by2_14_20_port, A_neg_shifted_by2_14_19_port, 
      A_neg_shifted_by2_14_18_port, A_neg_shifted_by2_14_17_port, 
      A_neg_shifted_by2_14_16_port, A_neg_shifted_by2_14_15_port, 
      A_neg_shifted_by2_14_14_port, A_neg_shifted_by2_14_13_port, 
      A_neg_shifted_by2_14_12_port, A_neg_shifted_by2_14_11_port, 
      A_neg_shifted_by2_14_10_port, A_neg_shifted_by2_14_9_port, 
      A_neg_shifted_by2_14_8_port, A_neg_shifted_by2_14_7_port, 
      A_neg_shifted_by2_14_6_port, A_neg_shifted_by2_14_5_port, 
      A_neg_shifted_by2_14_4_port, A_neg_shifted_by2_14_3_port, 
      A_neg_shifted_by2_14_2_port, A_neg_shifted_by2_14_1_port, 
      A_neg_shifted_by2_14_0_port, OUT_MUX_1_63_port, OUT_MUX_1_62_port, 
      OUT_MUX_1_61_port, OUT_MUX_1_60_port, OUT_MUX_1_59_port, 
      OUT_MUX_1_58_port, OUT_MUX_1_57_port, OUT_MUX_1_56_port, 
      OUT_MUX_1_55_port, OUT_MUX_1_54_port, OUT_MUX_1_53_port, 
      OUT_MUX_1_52_port, OUT_MUX_1_51_port, OUT_MUX_1_50_port, 
      OUT_MUX_1_49_port, OUT_MUX_1_48_port, OUT_MUX_1_47_port, 
      OUT_MUX_1_46_port, OUT_MUX_1_45_port, OUT_MUX_1_44_port, 
      OUT_MUX_1_43_port, OUT_MUX_1_42_port, OUT_MUX_1_41_port, 
      OUT_MUX_1_40_port, OUT_MUX_1_39_port, OUT_MUX_1_38_port, 
      OUT_MUX_1_37_port, OUT_MUX_1_36_port, OUT_MUX_1_35_port, 
      OUT_MUX_1_34_port, OUT_MUX_1_33_port, OUT_MUX_1_32_port, 
      OUT_MUX_1_31_port, OUT_MUX_1_30_port, OUT_MUX_1_29_port, 
      OUT_MUX_1_28_port, OUT_MUX_1_27_port, OUT_MUX_1_26_port, 
      OUT_MUX_1_25_port, OUT_MUX_1_24_port, OUT_MUX_1_23_port, 
      OUT_MUX_1_22_port, OUT_MUX_1_21_port, OUT_MUX_1_20_port, 
      OUT_MUX_1_19_port, OUT_MUX_1_18_port, OUT_MUX_1_17_port, 
      OUT_MUX_1_16_port, OUT_MUX_1_15_port, OUT_MUX_1_14_port, 
      OUT_MUX_1_13_port, OUT_MUX_1_12_port, OUT_MUX_1_11_port, 
      OUT_MUX_1_10_port, OUT_MUX_1_9_port, OUT_MUX_1_8_port, OUT_MUX_1_7_port, 
      OUT_MUX_1_6_port, OUT_MUX_1_5_port, OUT_MUX_1_4_port, OUT_MUX_1_3_port, 
      OUT_MUX_1_2_port, OUT_MUX_1_1_port, OUT_MUX_1_0_port, OUT_MUX_2_63_port, 
      OUT_MUX_2_62_port, OUT_MUX_2_61_port, OUT_MUX_2_60_port, 
      OUT_MUX_2_59_port, OUT_MUX_2_58_port, OUT_MUX_2_57_port, 
      OUT_MUX_2_56_port, OUT_MUX_2_55_port, OUT_MUX_2_54_port, 
      OUT_MUX_2_53_port, OUT_MUX_2_52_port, OUT_MUX_2_51_port, 
      OUT_MUX_2_50_port, OUT_MUX_2_49_port, OUT_MUX_2_48_port, 
      OUT_MUX_2_47_port, OUT_MUX_2_46_port, OUT_MUX_2_45_port, 
      OUT_MUX_2_44_port, OUT_MUX_2_43_port, OUT_MUX_2_42_port, 
      OUT_MUX_2_41_port, OUT_MUX_2_40_port, OUT_MUX_2_39_port, 
      OUT_MUX_2_38_port, OUT_MUX_2_37_port, OUT_MUX_2_36_port, 
      OUT_MUX_2_35_port, OUT_MUX_2_34_port, OUT_MUX_2_33_port, 
      OUT_MUX_2_32_port, OUT_MUX_2_31_port, OUT_MUX_2_30_port, 
      OUT_MUX_2_29_port, OUT_MUX_2_28_port, OUT_MUX_2_27_port, 
      OUT_MUX_2_26_port, OUT_MUX_2_25_port, OUT_MUX_2_24_port, 
      OUT_MUX_2_23_port, OUT_MUX_2_22_port, OUT_MUX_2_21_port, 
      OUT_MUX_2_20_port, OUT_MUX_2_19_port, OUT_MUX_2_18_port, 
      OUT_MUX_2_17_port, OUT_MUX_2_16_port, OUT_MUX_2_15_port, 
      OUT_MUX_2_14_port, OUT_MUX_2_13_port, OUT_MUX_2_12_port, 
      OUT_MUX_2_11_port, OUT_MUX_2_10_port, OUT_MUX_2_9_port, OUT_MUX_2_8_port,
      OUT_MUX_2_7_port, OUT_MUX_2_6_port, OUT_MUX_2_5_port, OUT_MUX_2_4_port, 
      OUT_MUX_2_3_port, OUT_MUX_2_2_port, OUT_MUX_2_1_port, OUT_MUX_2_0_port, 
      OUT_MUX_3_63_port, OUT_MUX_3_62_port, OUT_MUX_3_61_port, 
      OUT_MUX_3_60_port, OUT_MUX_3_59_port, OUT_MUX_3_58_port, 
      OUT_MUX_3_57_port, OUT_MUX_3_56_port, OUT_MUX_3_55_port, 
      OUT_MUX_3_54_port, OUT_MUX_3_53_port, OUT_MUX_3_52_port, 
      OUT_MUX_3_51_port, OUT_MUX_3_50_port, OUT_MUX_3_49_port, 
      OUT_MUX_3_48_port, OUT_MUX_3_47_port, OUT_MUX_3_46_port, 
      OUT_MUX_3_45_port, OUT_MUX_3_44_port, OUT_MUX_3_43_port, 
      OUT_MUX_3_42_port, OUT_MUX_3_41_port, OUT_MUX_3_40_port, 
      OUT_MUX_3_39_port, OUT_MUX_3_38_port, OUT_MUX_3_37_port, 
      OUT_MUX_3_36_port, OUT_MUX_3_35_port, OUT_MUX_3_34_port, 
      OUT_MUX_3_33_port, OUT_MUX_3_32_port, OUT_MUX_3_31_port, 
      OUT_MUX_3_30_port, OUT_MUX_3_29_port, OUT_MUX_3_28_port, 
      OUT_MUX_3_27_port, OUT_MUX_3_26_port, OUT_MUX_3_25_port, 
      OUT_MUX_3_24_port, OUT_MUX_3_23_port, OUT_MUX_3_22_port, 
      OUT_MUX_3_21_port, OUT_MUX_3_20_port, OUT_MUX_3_19_port, 
      OUT_MUX_3_18_port, OUT_MUX_3_17_port, OUT_MUX_3_16_port, 
      OUT_MUX_3_15_port, OUT_MUX_3_14_port, OUT_MUX_3_13_port, 
      OUT_MUX_3_12_port, OUT_MUX_3_11_port, OUT_MUX_3_10_port, OUT_MUX_3_9_port
      , OUT_MUX_3_8_port, OUT_MUX_3_7_port, OUT_MUX_3_6_port, OUT_MUX_3_5_port,
      OUT_MUX_3_4_port, OUT_MUX_3_3_port, OUT_MUX_3_2_port, OUT_MUX_3_1_port, 
      OUT_MUX_3_0_port, OUT_MUX_4_63_port, OUT_MUX_4_62_port, OUT_MUX_4_61_port
      , OUT_MUX_4_60_port, OUT_MUX_4_59_port, OUT_MUX_4_58_port, 
      OUT_MUX_4_57_port, OUT_MUX_4_56_port, OUT_MUX_4_55_port, 
      OUT_MUX_4_54_port, OUT_MUX_4_53_port, OUT_MUX_4_52_port, 
      OUT_MUX_4_51_port, OUT_MUX_4_50_port, OUT_MUX_4_49_port, 
      OUT_MUX_4_48_port, OUT_MUX_4_47_port, OUT_MUX_4_46_port, 
      OUT_MUX_4_45_port, OUT_MUX_4_44_port, OUT_MUX_4_43_port, 
      OUT_MUX_4_42_port, OUT_MUX_4_41_port, OUT_MUX_4_40_port, 
      OUT_MUX_4_39_port, OUT_MUX_4_38_port, OUT_MUX_4_37_port, 
      OUT_MUX_4_36_port, OUT_MUX_4_35_port, OUT_MUX_4_34_port, 
      OUT_MUX_4_33_port, OUT_MUX_4_32_port, OUT_MUX_4_31_port, 
      OUT_MUX_4_30_port, OUT_MUX_4_29_port, OUT_MUX_4_28_port, 
      OUT_MUX_4_27_port, OUT_MUX_4_26_port, OUT_MUX_4_25_port, 
      OUT_MUX_4_24_port, OUT_MUX_4_23_port, OUT_MUX_4_22_port, 
      OUT_MUX_4_21_port, OUT_MUX_4_20_port, OUT_MUX_4_19_port, 
      OUT_MUX_4_18_port, OUT_MUX_4_17_port, OUT_MUX_4_16_port, 
      OUT_MUX_4_15_port, OUT_MUX_4_14_port, OUT_MUX_4_13_port, 
      OUT_MUX_4_12_port, OUT_MUX_4_11_port, OUT_MUX_4_10_port, OUT_MUX_4_9_port
      , OUT_MUX_4_8_port, OUT_MUX_4_7_port, OUT_MUX_4_6_port, OUT_MUX_4_5_port,
      OUT_MUX_4_4_port, OUT_MUX_4_3_port, OUT_MUX_4_2_port, OUT_MUX_4_1_port, 
      OUT_MUX_4_0_port, OUT_MUX_5_63_port, OUT_MUX_5_62_port, OUT_MUX_5_61_port
      , OUT_MUX_5_60_port, OUT_MUX_5_59_port, OUT_MUX_5_58_port, 
      OUT_MUX_5_57_port, OUT_MUX_5_56_port, OUT_MUX_5_55_port, 
      OUT_MUX_5_54_port, OUT_MUX_5_53_port, OUT_MUX_5_52_port, 
      OUT_MUX_5_51_port, OUT_MUX_5_50_port, OUT_MUX_5_49_port, 
      OUT_MUX_5_48_port, OUT_MUX_5_47_port, OUT_MUX_5_46_port, 
      OUT_MUX_5_45_port, OUT_MUX_5_44_port, OUT_MUX_5_43_port, 
      OUT_MUX_5_42_port, OUT_MUX_5_41_port, OUT_MUX_5_40_port, 
      OUT_MUX_5_39_port, OUT_MUX_5_38_port, OUT_MUX_5_37_port, 
      OUT_MUX_5_36_port, OUT_MUX_5_35_port, OUT_MUX_5_34_port, 
      OUT_MUX_5_33_port, OUT_MUX_5_32_port, OUT_MUX_5_31_port, 
      OUT_MUX_5_30_port, OUT_MUX_5_29_port, OUT_MUX_5_28_port, 
      OUT_MUX_5_27_port, OUT_MUX_5_26_port, OUT_MUX_5_25_port, 
      OUT_MUX_5_24_port, OUT_MUX_5_23_port, OUT_MUX_5_22_port, 
      OUT_MUX_5_21_port, OUT_MUX_5_20_port, OUT_MUX_5_19_port, 
      OUT_MUX_5_18_port, OUT_MUX_5_17_port, OUT_MUX_5_16_port, 
      OUT_MUX_5_15_port, OUT_MUX_5_14_port, OUT_MUX_5_13_port, 
      OUT_MUX_5_12_port, OUT_MUX_5_11_port, OUT_MUX_5_10_port, OUT_MUX_5_9_port
      , OUT_MUX_5_8_port, OUT_MUX_5_7_port, OUT_MUX_5_6_port, OUT_MUX_5_5_port,
      OUT_MUX_5_4_port, OUT_MUX_5_3_port, OUT_MUX_5_2_port, OUT_MUX_5_1_port, 
      OUT_MUX_5_0_port, OUT_MUX_6_63_port, OUT_MUX_6_62_port, OUT_MUX_6_61_port
      , OUT_MUX_6_60_port, OUT_MUX_6_59_port, OUT_MUX_6_58_port, 
      OUT_MUX_6_57_port, OUT_MUX_6_56_port, OUT_MUX_6_55_port, 
      OUT_MUX_6_54_port, OUT_MUX_6_53_port, OUT_MUX_6_52_port, 
      OUT_MUX_6_51_port, OUT_MUX_6_50_port, OUT_MUX_6_49_port, 
      OUT_MUX_6_48_port, OUT_MUX_6_47_port, OUT_MUX_6_46_port, 
      OUT_MUX_6_45_port, OUT_MUX_6_44_port, OUT_MUX_6_43_port, 
      OUT_MUX_6_42_port, OUT_MUX_6_41_port, OUT_MUX_6_40_port, 
      OUT_MUX_6_39_port, OUT_MUX_6_38_port, OUT_MUX_6_37_port, 
      OUT_MUX_6_36_port, OUT_MUX_6_35_port, OUT_MUX_6_34_port, 
      OUT_MUX_6_33_port, OUT_MUX_6_32_port, OUT_MUX_6_31_port, 
      OUT_MUX_6_30_port, OUT_MUX_6_29_port, OUT_MUX_6_28_port, 
      OUT_MUX_6_27_port, OUT_MUX_6_26_port, OUT_MUX_6_25_port, 
      OUT_MUX_6_24_port, OUT_MUX_6_23_port, OUT_MUX_6_22_port, 
      OUT_MUX_6_21_port, OUT_MUX_6_20_port, OUT_MUX_6_19_port, 
      OUT_MUX_6_18_port, OUT_MUX_6_17_port, OUT_MUX_6_16_port, 
      OUT_MUX_6_15_port, OUT_MUX_6_14_port, OUT_MUX_6_13_port, 
      OUT_MUX_6_12_port, OUT_MUX_6_11_port, OUT_MUX_6_10_port, OUT_MUX_6_9_port
      , OUT_MUX_6_8_port, OUT_MUX_6_7_port, OUT_MUX_6_6_port, OUT_MUX_6_5_port,
      OUT_MUX_6_4_port, OUT_MUX_6_3_port, OUT_MUX_6_2_port, OUT_MUX_6_1_port, 
      OUT_MUX_6_0_port, OUT_MUX_7_63_port, OUT_MUX_7_62_port, OUT_MUX_7_61_port
      , OUT_MUX_7_60_port, OUT_MUX_7_59_port, OUT_MUX_7_58_port, 
      OUT_MUX_7_57_port, OUT_MUX_7_56_port, OUT_MUX_7_55_port, 
      OUT_MUX_7_54_port, OUT_MUX_7_53_port, OUT_MUX_7_52_port, 
      OUT_MUX_7_51_port, OUT_MUX_7_50_port, OUT_MUX_7_49_port, 
      OUT_MUX_7_48_port, OUT_MUX_7_47_port, OUT_MUX_7_46_port, 
      OUT_MUX_7_45_port, OUT_MUX_7_44_port, OUT_MUX_7_43_port, 
      OUT_MUX_7_42_port, OUT_MUX_7_41_port, OUT_MUX_7_40_port, 
      OUT_MUX_7_39_port, OUT_MUX_7_38_port, OUT_MUX_7_37_port, 
      OUT_MUX_7_36_port, OUT_MUX_7_35_port, OUT_MUX_7_34_port, 
      OUT_MUX_7_33_port, OUT_MUX_7_32_port, OUT_MUX_7_31_port, 
      OUT_MUX_7_30_port, OUT_MUX_7_29_port, OUT_MUX_7_28_port, 
      OUT_MUX_7_27_port, OUT_MUX_7_26_port, OUT_MUX_7_25_port, 
      OUT_MUX_7_24_port, OUT_MUX_7_23_port, OUT_MUX_7_22_port, 
      OUT_MUX_7_21_port, OUT_MUX_7_20_port, OUT_MUX_7_19_port, 
      OUT_MUX_7_18_port, OUT_MUX_7_17_port, OUT_MUX_7_16_port, 
      OUT_MUX_7_15_port, OUT_MUX_7_14_port, OUT_MUX_7_13_port, 
      OUT_MUX_7_12_port, OUT_MUX_7_11_port, OUT_MUX_7_10_port, OUT_MUX_7_9_port
      , OUT_MUX_7_8_port, OUT_MUX_7_7_port, OUT_MUX_7_6_port, OUT_MUX_7_5_port,
      OUT_MUX_7_4_port, OUT_MUX_7_3_port, OUT_MUX_7_2_port, OUT_MUX_7_1_port, 
      OUT_MUX_7_0_port, OUT_MUX_8_63_port, OUT_MUX_8_62_port, OUT_MUX_8_61_port
      , OUT_MUX_8_60_port, OUT_MUX_8_59_port, OUT_MUX_8_58_port, 
      OUT_MUX_8_57_port, OUT_MUX_8_56_port, OUT_MUX_8_55_port, 
      OUT_MUX_8_54_port, OUT_MUX_8_53_port, OUT_MUX_8_52_port, 
      OUT_MUX_8_51_port, OUT_MUX_8_50_port, OUT_MUX_8_49_port, 
      OUT_MUX_8_48_port, OUT_MUX_8_47_port, OUT_MUX_8_46_port, 
      OUT_MUX_8_45_port, OUT_MUX_8_44_port, OUT_MUX_8_43_port, 
      OUT_MUX_8_42_port, OUT_MUX_8_41_port, OUT_MUX_8_40_port, 
      OUT_MUX_8_39_port, OUT_MUX_8_38_port, OUT_MUX_8_37_port, 
      OUT_MUX_8_36_port, OUT_MUX_8_35_port, OUT_MUX_8_34_port, 
      OUT_MUX_8_33_port, OUT_MUX_8_32_port, OUT_MUX_8_31_port, 
      OUT_MUX_8_30_port, OUT_MUX_8_29_port, OUT_MUX_8_28_port, 
      OUT_MUX_8_27_port, OUT_MUX_8_26_port, OUT_MUX_8_25_port, 
      OUT_MUX_8_24_port, OUT_MUX_8_23_port, OUT_MUX_8_22_port, 
      OUT_MUX_8_21_port, OUT_MUX_8_20_port, OUT_MUX_8_19_port, 
      OUT_MUX_8_18_port, OUT_MUX_8_17_port, OUT_MUX_8_16_port, 
      OUT_MUX_8_15_port, OUT_MUX_8_14_port, OUT_MUX_8_13_port, 
      OUT_MUX_8_12_port, OUT_MUX_8_11_port, OUT_MUX_8_10_port, OUT_MUX_8_9_port
      , OUT_MUX_8_8_port, OUT_MUX_8_7_port, OUT_MUX_8_6_port, OUT_MUX_8_5_port,
      OUT_MUX_8_4_port, OUT_MUX_8_3_port, OUT_MUX_8_2_port, OUT_MUX_8_1_port, 
      OUT_MUX_8_0_port, OUT_MUX_9_63_port, OUT_MUX_9_62_port, OUT_MUX_9_61_port
      , OUT_MUX_9_60_port, OUT_MUX_9_59_port, OUT_MUX_9_58_port, 
      OUT_MUX_9_57_port, OUT_MUX_9_56_port, OUT_MUX_9_55_port, 
      OUT_MUX_9_54_port, OUT_MUX_9_53_port, OUT_MUX_9_52_port, 
      OUT_MUX_9_51_port, OUT_MUX_9_50_port, OUT_MUX_9_49_port, 
      OUT_MUX_9_48_port, OUT_MUX_9_47_port, OUT_MUX_9_46_port, 
      OUT_MUX_9_45_port, OUT_MUX_9_44_port, OUT_MUX_9_43_port, 
      OUT_MUX_9_42_port, OUT_MUX_9_41_port, OUT_MUX_9_40_port, 
      OUT_MUX_9_39_port, OUT_MUX_9_38_port, OUT_MUX_9_37_port, 
      OUT_MUX_9_36_port, OUT_MUX_9_35_port, OUT_MUX_9_34_port, 
      OUT_MUX_9_33_port, OUT_MUX_9_32_port, OUT_MUX_9_31_port, 
      OUT_MUX_9_30_port, OUT_MUX_9_29_port, OUT_MUX_9_28_port, 
      OUT_MUX_9_27_port, OUT_MUX_9_26_port, OUT_MUX_9_25_port, 
      OUT_MUX_9_24_port, OUT_MUX_9_23_port, OUT_MUX_9_22_port, 
      OUT_MUX_9_21_port, OUT_MUX_9_20_port, OUT_MUX_9_19_port, 
      OUT_MUX_9_18_port, OUT_MUX_9_17_port, OUT_MUX_9_16_port, 
      OUT_MUX_9_15_port, OUT_MUX_9_14_port, OUT_MUX_9_13_port, 
      OUT_MUX_9_12_port, OUT_MUX_9_11_port, OUT_MUX_9_10_port, OUT_MUX_9_9_port
      , OUT_MUX_9_8_port, OUT_MUX_9_7_port, OUT_MUX_9_6_port, OUT_MUX_9_5_port,
      OUT_MUX_9_4_port, OUT_MUX_9_3_port, OUT_MUX_9_2_port, OUT_MUX_9_1_port, 
      OUT_MUX_9_0_port, OUT_MUX_10_63_port, OUT_MUX_10_62_port, 
      OUT_MUX_10_61_port, OUT_MUX_10_60_port, OUT_MUX_10_59_port, 
      OUT_MUX_10_58_port, OUT_MUX_10_57_port, OUT_MUX_10_56_port, 
      OUT_MUX_10_55_port, OUT_MUX_10_54_port, OUT_MUX_10_53_port, 
      OUT_MUX_10_52_port, OUT_MUX_10_51_port, OUT_MUX_10_50_port, 
      OUT_MUX_10_49_port, OUT_MUX_10_48_port, OUT_MUX_10_47_port, 
      OUT_MUX_10_46_port, OUT_MUX_10_45_port, OUT_MUX_10_44_port, 
      OUT_MUX_10_43_port, OUT_MUX_10_42_port, OUT_MUX_10_41_port, 
      OUT_MUX_10_40_port, OUT_MUX_10_39_port, OUT_MUX_10_38_port, 
      OUT_MUX_10_37_port, OUT_MUX_10_36_port, OUT_MUX_10_35_port, 
      OUT_MUX_10_34_port, OUT_MUX_10_33_port, OUT_MUX_10_32_port, 
      OUT_MUX_10_31_port, OUT_MUX_10_30_port, OUT_MUX_10_29_port, 
      OUT_MUX_10_28_port, OUT_MUX_10_27_port, OUT_MUX_10_26_port, 
      OUT_MUX_10_25_port, OUT_MUX_10_24_port, OUT_MUX_10_23_port, 
      OUT_MUX_10_22_port, OUT_MUX_10_21_port, OUT_MUX_10_20_port, 
      OUT_MUX_10_19_port, OUT_MUX_10_18_port, OUT_MUX_10_17_port, 
      OUT_MUX_10_16_port, OUT_MUX_10_15_port, OUT_MUX_10_14_port, 
      OUT_MUX_10_13_port, OUT_MUX_10_12_port, OUT_MUX_10_11_port, 
      OUT_MUX_10_10_port, OUT_MUX_10_9_port, OUT_MUX_10_8_port, 
      OUT_MUX_10_7_port, OUT_MUX_10_6_port, OUT_MUX_10_5_port, 
      OUT_MUX_10_4_port, OUT_MUX_10_3_port, OUT_MUX_10_2_port, 
      OUT_MUX_10_1_port, OUT_MUX_10_0_port, OUT_MUX_11_63_port, 
      OUT_MUX_11_62_port, OUT_MUX_11_61_port, OUT_MUX_11_60_port, 
      OUT_MUX_11_59_port, OUT_MUX_11_58_port, OUT_MUX_11_57_port, 
      OUT_MUX_11_56_port, OUT_MUX_11_55_port, OUT_MUX_11_54_port, 
      OUT_MUX_11_53_port, OUT_MUX_11_52_port, OUT_MUX_11_51_port, 
      OUT_MUX_11_50_port, OUT_MUX_11_49_port, OUT_MUX_11_48_port, 
      OUT_MUX_11_47_port, OUT_MUX_11_46_port, OUT_MUX_11_45_port, 
      OUT_MUX_11_44_port, OUT_MUX_11_43_port, OUT_MUX_11_42_port, 
      OUT_MUX_11_41_port, OUT_MUX_11_40_port, OUT_MUX_11_39_port, 
      OUT_MUX_11_38_port, OUT_MUX_11_37_port, OUT_MUX_11_36_port, 
      OUT_MUX_11_35_port, OUT_MUX_11_34_port, OUT_MUX_11_33_port, 
      OUT_MUX_11_32_port, OUT_MUX_11_31_port, OUT_MUX_11_30_port, 
      OUT_MUX_11_29_port, OUT_MUX_11_28_port, OUT_MUX_11_27_port, 
      OUT_MUX_11_26_port, OUT_MUX_11_25_port, OUT_MUX_11_24_port, 
      OUT_MUX_11_23_port, OUT_MUX_11_22_port, OUT_MUX_11_21_port, 
      OUT_MUX_11_20_port, OUT_MUX_11_19_port, OUT_MUX_11_18_port, 
      OUT_MUX_11_17_port, OUT_MUX_11_16_port, OUT_MUX_11_15_port, 
      OUT_MUX_11_14_port, OUT_MUX_11_13_port, OUT_MUX_11_12_port, 
      OUT_MUX_11_11_port, OUT_MUX_11_10_port, OUT_MUX_11_9_port, 
      OUT_MUX_11_8_port, OUT_MUX_11_7_port, OUT_MUX_11_6_port, 
      OUT_MUX_11_5_port, OUT_MUX_11_4_port, OUT_MUX_11_3_port, 
      OUT_MUX_11_2_port, OUT_MUX_11_1_port, OUT_MUX_11_0_port, 
      OUT_MUX_12_63_port, OUT_MUX_12_62_port, OUT_MUX_12_61_port, 
      OUT_MUX_12_60_port, OUT_MUX_12_59_port, OUT_MUX_12_58_port, 
      OUT_MUX_12_57_port, OUT_MUX_12_56_port, OUT_MUX_12_55_port, 
      OUT_MUX_12_54_port, OUT_MUX_12_53_port, OUT_MUX_12_52_port, 
      OUT_MUX_12_51_port, OUT_MUX_12_50_port, OUT_MUX_12_49_port, 
      OUT_MUX_12_48_port, OUT_MUX_12_47_port, OUT_MUX_12_46_port, 
      OUT_MUX_12_45_port, OUT_MUX_12_44_port, OUT_MUX_12_43_port, 
      OUT_MUX_12_42_port, OUT_MUX_12_41_port, OUT_MUX_12_40_port, 
      OUT_MUX_12_39_port, OUT_MUX_12_38_port, OUT_MUX_12_37_port, 
      OUT_MUX_12_36_port, OUT_MUX_12_35_port, OUT_MUX_12_34_port, 
      OUT_MUX_12_33_port, OUT_MUX_12_32_port, OUT_MUX_12_31_port, 
      OUT_MUX_12_30_port, OUT_MUX_12_29_port, OUT_MUX_12_28_port, 
      OUT_MUX_12_27_port, OUT_MUX_12_26_port, OUT_MUX_12_25_port, 
      OUT_MUX_12_24_port, OUT_MUX_12_23_port, OUT_MUX_12_22_port, 
      OUT_MUX_12_21_port, OUT_MUX_12_20_port, OUT_MUX_12_19_port, 
      OUT_MUX_12_18_port, OUT_MUX_12_17_port, OUT_MUX_12_16_port, 
      OUT_MUX_12_15_port, OUT_MUX_12_14_port, OUT_MUX_12_13_port, 
      OUT_MUX_12_12_port, OUT_MUX_12_11_port, OUT_MUX_12_10_port, 
      OUT_MUX_12_9_port, OUT_MUX_12_8_port, OUT_MUX_12_7_port, 
      OUT_MUX_12_6_port, OUT_MUX_12_5_port, OUT_MUX_12_4_port, 
      OUT_MUX_12_3_port, OUT_MUX_12_2_port, OUT_MUX_12_1_port, 
      OUT_MUX_12_0_port, OUT_MUX_13_63_port, OUT_MUX_13_62_port, 
      OUT_MUX_13_61_port, OUT_MUX_13_60_port, OUT_MUX_13_59_port, 
      OUT_MUX_13_58_port, OUT_MUX_13_57_port, OUT_MUX_13_56_port, 
      OUT_MUX_13_55_port, OUT_MUX_13_54_port, OUT_MUX_13_53_port, 
      OUT_MUX_13_52_port, OUT_MUX_13_51_port, OUT_MUX_13_50_port, 
      OUT_MUX_13_49_port, OUT_MUX_13_48_port, OUT_MUX_13_47_port, 
      OUT_MUX_13_46_port, OUT_MUX_13_45_port, OUT_MUX_13_44_port, 
      OUT_MUX_13_43_port, OUT_MUX_13_42_port, OUT_MUX_13_41_port, 
      OUT_MUX_13_40_port, OUT_MUX_13_39_port, OUT_MUX_13_38_port, 
      OUT_MUX_13_37_port, OUT_MUX_13_36_port, OUT_MUX_13_35_port, 
      OUT_MUX_13_34_port, OUT_MUX_13_33_port, OUT_MUX_13_32_port, 
      OUT_MUX_13_31_port, OUT_MUX_13_30_port, OUT_MUX_13_29_port, 
      OUT_MUX_13_28_port, OUT_MUX_13_27_port, OUT_MUX_13_26_port, 
      OUT_MUX_13_25_port, OUT_MUX_13_24_port, OUT_MUX_13_23_port, 
      OUT_MUX_13_22_port, OUT_MUX_13_21_port, OUT_MUX_13_20_port, 
      OUT_MUX_13_19_port, OUT_MUX_13_18_port, OUT_MUX_13_17_port, 
      OUT_MUX_13_16_port, OUT_MUX_13_15_port, OUT_MUX_13_14_port, 
      OUT_MUX_13_13_port, OUT_MUX_13_12_port, OUT_MUX_13_11_port, 
      OUT_MUX_13_10_port, OUT_MUX_13_9_port, OUT_MUX_13_8_port, 
      OUT_MUX_13_7_port, OUT_MUX_13_6_port, OUT_MUX_13_5_port, 
      OUT_MUX_13_4_port, OUT_MUX_13_3_port, OUT_MUX_13_2_port, 
      OUT_MUX_13_1_port, OUT_MUX_13_0_port, OUT_MUX_14_63_port, 
      OUT_MUX_14_62_port, OUT_MUX_14_61_port, OUT_MUX_14_60_port, 
      OUT_MUX_14_59_port, OUT_MUX_14_58_port, OUT_MUX_14_57_port, 
      OUT_MUX_14_56_port, OUT_MUX_14_55_port, OUT_MUX_14_54_port, 
      OUT_MUX_14_53_port, OUT_MUX_14_52_port, OUT_MUX_14_51_port, 
      OUT_MUX_14_50_port, OUT_MUX_14_49_port, OUT_MUX_14_48_port, 
      OUT_MUX_14_47_port, OUT_MUX_14_46_port, OUT_MUX_14_45_port, 
      OUT_MUX_14_44_port, OUT_MUX_14_43_port, OUT_MUX_14_42_port, 
      OUT_MUX_14_41_port, OUT_MUX_14_40_port, OUT_MUX_14_39_port, 
      OUT_MUX_14_38_port, OUT_MUX_14_37_port, OUT_MUX_14_36_port, 
      OUT_MUX_14_35_port, OUT_MUX_14_34_port, OUT_MUX_14_33_port, 
      OUT_MUX_14_32_port, OUT_MUX_14_31_port, OUT_MUX_14_30_port, 
      OUT_MUX_14_29_port, OUT_MUX_14_28_port, OUT_MUX_14_27_port, 
      OUT_MUX_14_26_port, OUT_MUX_14_25_port, OUT_MUX_14_24_port, 
      OUT_MUX_14_23_port, OUT_MUX_14_22_port, OUT_MUX_14_21_port, 
      OUT_MUX_14_20_port, OUT_MUX_14_19_port, OUT_MUX_14_18_port, 
      OUT_MUX_14_17_port, OUT_MUX_14_16_port, OUT_MUX_14_15_port, 
      OUT_MUX_14_14_port, OUT_MUX_14_13_port, OUT_MUX_14_12_port, 
      OUT_MUX_14_11_port, OUT_MUX_14_10_port, OUT_MUX_14_9_port, 
      OUT_MUX_14_8_port, OUT_MUX_14_7_port, OUT_MUX_14_6_port, 
      OUT_MUX_14_5_port, OUT_MUX_14_4_port, OUT_MUX_14_3_port, 
      OUT_MUX_14_2_port, OUT_MUX_14_1_port, OUT_MUX_14_0_port, 
      OUT_MUX_15_63_port, OUT_MUX_15_62_port, OUT_MUX_15_61_port, 
      OUT_MUX_15_60_port, OUT_MUX_15_59_port, OUT_MUX_15_58_port, 
      OUT_MUX_15_57_port, OUT_MUX_15_56_port, OUT_MUX_15_55_port, 
      OUT_MUX_15_54_port, OUT_MUX_15_53_port, OUT_MUX_15_52_port, 
      OUT_MUX_15_51_port, OUT_MUX_15_50_port, OUT_MUX_15_49_port, 
      OUT_MUX_15_48_port, OUT_MUX_15_47_port, OUT_MUX_15_46_port, 
      OUT_MUX_15_45_port, OUT_MUX_15_44_port, OUT_MUX_15_43_port, 
      OUT_MUX_15_42_port, OUT_MUX_15_41_port, OUT_MUX_15_40_port, 
      OUT_MUX_15_39_port, OUT_MUX_15_38_port, OUT_MUX_15_37_port, 
      OUT_MUX_15_36_port, OUT_MUX_15_35_port, OUT_MUX_15_34_port, 
      OUT_MUX_15_33_port, OUT_MUX_15_32_port, OUT_MUX_15_31_port, 
      OUT_MUX_15_30_port, OUT_MUX_15_29_port, OUT_MUX_15_28_port, 
      OUT_MUX_15_27_port, OUT_MUX_15_26_port, OUT_MUX_15_25_port, 
      OUT_MUX_15_24_port, OUT_MUX_15_23_port, OUT_MUX_15_22_port, 
      OUT_MUX_15_21_port, OUT_MUX_15_20_port, OUT_MUX_15_19_port, 
      OUT_MUX_15_18_port, OUT_MUX_15_17_port, OUT_MUX_15_16_port, 
      OUT_MUX_15_15_port, OUT_MUX_15_14_port, OUT_MUX_15_13_port, 
      OUT_MUX_15_12_port, OUT_MUX_15_11_port, OUT_MUX_15_10_port, 
      OUT_MUX_15_9_port, OUT_MUX_15_8_port, OUT_MUX_15_7_port, 
      OUT_MUX_15_6_port, OUT_MUX_15_5_port, OUT_MUX_15_4_port, 
      OUT_MUX_15_3_port, OUT_MUX_15_2_port, OUT_MUX_15_1_port, 
      OUT_MUX_15_0_port, P_tmp_0_63_port, P_tmp_0_62_port, P_tmp_0_61_port, 
      P_tmp_0_60_port, P_tmp_0_59_port, P_tmp_0_58_port, P_tmp_0_57_port, 
      P_tmp_0_56_port, P_tmp_0_55_port, P_tmp_0_54_port, P_tmp_0_53_port, 
      P_tmp_0_52_port, P_tmp_0_51_port, P_tmp_0_50_port, P_tmp_0_49_port, 
      P_tmp_0_48_port, P_tmp_0_47_port, P_tmp_0_46_port, P_tmp_0_45_port, 
      P_tmp_0_44_port, P_tmp_0_43_port, P_tmp_0_42_port, P_tmp_0_41_port, 
      P_tmp_0_40_port, P_tmp_0_39_port, P_tmp_0_38_port, P_tmp_0_37_port, 
      P_tmp_0_36_port, P_tmp_0_35_port, P_tmp_0_34_port, P_tmp_0_33_port, 
      P_tmp_0_32_port, P_tmp_0_31_port, P_tmp_0_30_port, P_tmp_0_29_port, 
      P_tmp_0_28_port, P_tmp_0_27_port, P_tmp_0_26_port, P_tmp_0_25_port, 
      P_tmp_0_24_port, P_tmp_0_23_port, P_tmp_0_22_port, P_tmp_0_21_port, 
      P_tmp_0_20_port, P_tmp_0_19_port, P_tmp_0_18_port, P_tmp_0_17_port, 
      P_tmp_0_16_port, P_tmp_0_15_port, P_tmp_0_14_port, P_tmp_0_13_port, 
      P_tmp_0_12_port, P_tmp_0_11_port, P_tmp_0_10_port, P_tmp_0_9_port, 
      P_tmp_0_8_port, P_tmp_0_7_port, P_tmp_0_6_port, P_tmp_0_5_port, 
      P_tmp_0_4_port, P_tmp_0_3_port, P_tmp_0_2_port, P_tmp_0_1_port, 
      P_tmp_0_0_port, P_tmp_1_63_port, P_tmp_1_62_port, P_tmp_1_61_port, 
      P_tmp_1_60_port, P_tmp_1_59_port, P_tmp_1_58_port, P_tmp_1_57_port, 
      P_tmp_1_56_port, P_tmp_1_55_port, P_tmp_1_54_port, P_tmp_1_53_port, 
      P_tmp_1_52_port, P_tmp_1_51_port, P_tmp_1_50_port, P_tmp_1_49_port, 
      P_tmp_1_48_port, P_tmp_1_47_port, P_tmp_1_46_port, P_tmp_1_45_port, 
      P_tmp_1_44_port, P_tmp_1_43_port, P_tmp_1_42_port, P_tmp_1_41_port, 
      P_tmp_1_40_port, P_tmp_1_39_port, P_tmp_1_38_port, P_tmp_1_37_port, 
      P_tmp_1_36_port, P_tmp_1_35_port, P_tmp_1_34_port, P_tmp_1_33_port, 
      P_tmp_1_32_port, P_tmp_1_31_port, P_tmp_1_30_port, P_tmp_1_29_port, 
      P_tmp_1_28_port, P_tmp_1_27_port, P_tmp_1_26_port, P_tmp_1_25_port, 
      P_tmp_1_24_port, P_tmp_1_23_port, P_tmp_1_22_port, P_tmp_1_21_port, 
      P_tmp_1_20_port, P_tmp_1_19_port, P_tmp_1_18_port, P_tmp_1_17_port, 
      P_tmp_1_16_port, P_tmp_1_15_port, P_tmp_1_14_port, P_tmp_1_13_port, 
      P_tmp_1_12_port, P_tmp_1_11_port, P_tmp_1_10_port, P_tmp_1_9_port, 
      P_tmp_1_8_port, P_tmp_1_7_port, P_tmp_1_6_port, P_tmp_1_5_port, 
      P_tmp_1_4_port, P_tmp_1_3_port, P_tmp_1_2_port, P_tmp_1_1_port, 
      P_tmp_1_0_port, P_tmp_2_63_port, P_tmp_2_62_port, P_tmp_2_61_port, 
      P_tmp_2_60_port, P_tmp_2_59_port, P_tmp_2_58_port, P_tmp_2_57_port, 
      P_tmp_2_56_port, P_tmp_2_55_port, P_tmp_2_54_port, P_tmp_2_53_port, 
      P_tmp_2_52_port, P_tmp_2_51_port, P_tmp_2_50_port, P_tmp_2_49_port, 
      P_tmp_2_48_port, P_tmp_2_47_port, P_tmp_2_46_port, P_tmp_2_45_port, 
      P_tmp_2_44_port, P_tmp_2_43_port, P_tmp_2_42_port, P_tmp_2_41_port, 
      P_tmp_2_40_port, P_tmp_2_39_port, P_tmp_2_38_port, P_tmp_2_37_port, 
      P_tmp_2_36_port, P_tmp_2_35_port, P_tmp_2_34_port, P_tmp_2_33_port, 
      P_tmp_2_32_port, P_tmp_2_31_port, P_tmp_2_30_port, P_tmp_2_29_port, 
      P_tmp_2_28_port, P_tmp_2_27_port, P_tmp_2_26_port, P_tmp_2_25_port, 
      P_tmp_2_24_port, P_tmp_2_23_port, P_tmp_2_22_port, P_tmp_2_21_port, 
      P_tmp_2_20_port, P_tmp_2_19_port, P_tmp_2_18_port, P_tmp_2_17_port, 
      P_tmp_2_16_port, P_tmp_2_15_port, P_tmp_2_14_port, P_tmp_2_13_port, 
      P_tmp_2_12_port, P_tmp_2_11_port, P_tmp_2_10_port, P_tmp_2_9_port, 
      P_tmp_2_8_port, P_tmp_2_7_port, P_tmp_2_6_port, P_tmp_2_5_port, 
      P_tmp_2_4_port, P_tmp_2_3_port, P_tmp_2_2_port, P_tmp_2_1_port, 
      P_tmp_2_0_port, P_tmp_3_63_port, P_tmp_3_62_port, P_tmp_3_61_port, 
      P_tmp_3_60_port, P_tmp_3_59_port, P_tmp_3_58_port, P_tmp_3_57_port, 
      P_tmp_3_56_port, P_tmp_3_55_port, P_tmp_3_54_port, P_tmp_3_53_port, 
      P_tmp_3_52_port, P_tmp_3_51_port, P_tmp_3_50_port, P_tmp_3_49_port, 
      P_tmp_3_48_port, P_tmp_3_47_port, P_tmp_3_46_port, P_tmp_3_45_port, 
      P_tmp_3_44_port, P_tmp_3_43_port, P_tmp_3_42_port, P_tmp_3_41_port, 
      P_tmp_3_40_port, P_tmp_3_39_port, P_tmp_3_38_port, P_tmp_3_37_port, 
      P_tmp_3_36_port, P_tmp_3_35_port, P_tmp_3_34_port, P_tmp_3_33_port, 
      P_tmp_3_32_port, P_tmp_3_31_port, P_tmp_3_30_port, P_tmp_3_29_port, 
      P_tmp_3_28_port, P_tmp_3_27_port, P_tmp_3_26_port, P_tmp_3_25_port, 
      P_tmp_3_24_port, P_tmp_3_23_port, P_tmp_3_22_port, P_tmp_3_21_port, 
      P_tmp_3_20_port, P_tmp_3_19_port, P_tmp_3_18_port, P_tmp_3_17_port, 
      P_tmp_3_16_port, P_tmp_3_15_port, P_tmp_3_14_port, P_tmp_3_13_port, 
      P_tmp_3_12_port, P_tmp_3_11_port, P_tmp_3_10_port, P_tmp_3_9_port, 
      P_tmp_3_8_port, P_tmp_3_7_port, P_tmp_3_6_port, P_tmp_3_5_port, 
      P_tmp_3_4_port, P_tmp_3_3_port, P_tmp_3_2_port, P_tmp_3_1_port, 
      P_tmp_3_0_port, P_tmp_4_63_port, P_tmp_4_62_port, P_tmp_4_61_port, 
      P_tmp_4_60_port, P_tmp_4_59_port, P_tmp_4_58_port, P_tmp_4_57_port, 
      P_tmp_4_56_port, P_tmp_4_55_port, P_tmp_4_54_port, P_tmp_4_53_port, 
      P_tmp_4_52_port, P_tmp_4_51_port, P_tmp_4_50_port, P_tmp_4_49_port, 
      P_tmp_4_48_port, P_tmp_4_47_port, P_tmp_4_46_port, P_tmp_4_45_port, 
      P_tmp_4_44_port, P_tmp_4_43_port, P_tmp_4_42_port, P_tmp_4_41_port, 
      P_tmp_4_40_port, P_tmp_4_39_port, P_tmp_4_38_port, P_tmp_4_37_port, 
      P_tmp_4_36_port, P_tmp_4_35_port, P_tmp_4_34_port, P_tmp_4_33_port, 
      P_tmp_4_32_port, P_tmp_4_31_port, P_tmp_4_30_port, P_tmp_4_29_port, 
      P_tmp_4_28_port, P_tmp_4_27_port, P_tmp_4_26_port, P_tmp_4_25_port, 
      P_tmp_4_24_port, P_tmp_4_23_port, P_tmp_4_22_port, P_tmp_4_21_port, 
      P_tmp_4_20_port, P_tmp_4_19_port, P_tmp_4_18_port, P_tmp_4_17_port, 
      P_tmp_4_16_port, P_tmp_4_15_port, P_tmp_4_14_port, P_tmp_4_13_port, 
      P_tmp_4_12_port, P_tmp_4_11_port, P_tmp_4_10_port, P_tmp_4_9_port, 
      P_tmp_4_8_port, P_tmp_4_7_port, P_tmp_4_6_port, P_tmp_4_5_port, 
      P_tmp_4_4_port, P_tmp_4_3_port, P_tmp_4_2_port, P_tmp_4_1_port, 
      P_tmp_4_0_port, P_tmp_5_63_port, P_tmp_5_62_port, P_tmp_5_61_port, 
      P_tmp_5_60_port, P_tmp_5_59_port, P_tmp_5_58_port, P_tmp_5_57_port, 
      P_tmp_5_56_port, P_tmp_5_55_port, P_tmp_5_54_port, P_tmp_5_53_port, 
      P_tmp_5_52_port, P_tmp_5_51_port, P_tmp_5_50_port, P_tmp_5_49_port, 
      P_tmp_5_48_port, P_tmp_5_47_port, P_tmp_5_46_port, P_tmp_5_45_port, 
      P_tmp_5_44_port, P_tmp_5_43_port, P_tmp_5_42_port, P_tmp_5_41_port, 
      P_tmp_5_40_port, P_tmp_5_39_port, P_tmp_5_38_port, P_tmp_5_37_port, 
      P_tmp_5_36_port, P_tmp_5_35_port, P_tmp_5_34_port, P_tmp_5_33_port, 
      P_tmp_5_32_port, P_tmp_5_31_port, P_tmp_5_30_port, P_tmp_5_29_port, 
      P_tmp_5_28_port, P_tmp_5_27_port, P_tmp_5_26_port, P_tmp_5_25_port, 
      P_tmp_5_24_port, P_tmp_5_23_port, P_tmp_5_22_port, P_tmp_5_21_port, 
      P_tmp_5_20_port, P_tmp_5_19_port, P_tmp_5_18_port, P_tmp_5_17_port, 
      P_tmp_5_16_port, P_tmp_5_15_port, P_tmp_5_14_port, P_tmp_5_13_port, 
      P_tmp_5_12_port, P_tmp_5_11_port, P_tmp_5_10_port, P_tmp_5_9_port, 
      P_tmp_5_8_port, P_tmp_5_7_port, P_tmp_5_6_port, P_tmp_5_5_port, 
      P_tmp_5_4_port, P_tmp_5_3_port, P_tmp_5_2_port, P_tmp_5_1_port, 
      P_tmp_5_0_port, P_tmp_6_63_port, P_tmp_6_62_port, P_tmp_6_61_port, 
      P_tmp_6_60_port, P_tmp_6_59_port, P_tmp_6_58_port, P_tmp_6_57_port, 
      P_tmp_6_56_port, P_tmp_6_55_port, P_tmp_6_54_port, P_tmp_6_53_port, 
      P_tmp_6_52_port, P_tmp_6_51_port, P_tmp_6_50_port, P_tmp_6_49_port, 
      P_tmp_6_48_port, P_tmp_6_47_port, P_tmp_6_46_port, P_tmp_6_45_port, 
      P_tmp_6_44_port, P_tmp_6_43_port, P_tmp_6_42_port, P_tmp_6_41_port, 
      P_tmp_6_40_port, P_tmp_6_39_port, P_tmp_6_38_port, P_tmp_6_37_port, 
      P_tmp_6_36_port, P_tmp_6_35_port, P_tmp_6_34_port, P_tmp_6_33_port, 
      P_tmp_6_32_port, P_tmp_6_31_port, P_tmp_6_30_port, P_tmp_6_29_port, 
      P_tmp_6_28_port, P_tmp_6_27_port, P_tmp_6_26_port, P_tmp_6_25_port, 
      P_tmp_6_24_port, P_tmp_6_23_port, P_tmp_6_22_port, P_tmp_6_21_port, 
      P_tmp_6_20_port, P_tmp_6_19_port, P_tmp_6_18_port, P_tmp_6_17_port, 
      P_tmp_6_16_port, P_tmp_6_15_port, P_tmp_6_14_port, P_tmp_6_13_port, 
      P_tmp_6_12_port, P_tmp_6_11_port, P_tmp_6_10_port, P_tmp_6_9_port, 
      P_tmp_6_8_port, P_tmp_6_7_port, P_tmp_6_6_port, P_tmp_6_5_port, 
      P_tmp_6_4_port, P_tmp_6_3_port, P_tmp_6_2_port, P_tmp_6_1_port, 
      P_tmp_6_0_port, P_tmp_7_63_port, P_tmp_7_62_port, P_tmp_7_61_port, 
      P_tmp_7_60_port, P_tmp_7_59_port, P_tmp_7_58_port, P_tmp_7_57_port, 
      P_tmp_7_56_port, P_tmp_7_55_port, P_tmp_7_54_port, P_tmp_7_53_port, 
      P_tmp_7_52_port, P_tmp_7_51_port, P_tmp_7_50_port, P_tmp_7_49_port, 
      P_tmp_7_48_port, P_tmp_7_47_port, P_tmp_7_46_port, P_tmp_7_45_port, 
      P_tmp_7_44_port, P_tmp_7_43_port, P_tmp_7_42_port, P_tmp_7_41_port, 
      P_tmp_7_40_port, P_tmp_7_39_port, P_tmp_7_38_port, P_tmp_7_37_port, 
      P_tmp_7_36_port, P_tmp_7_35_port, P_tmp_7_34_port, P_tmp_7_33_port, 
      P_tmp_7_32_port, P_tmp_7_31_port, P_tmp_7_30_port, P_tmp_7_29_port, 
      P_tmp_7_28_port, P_tmp_7_27_port, P_tmp_7_26_port, P_tmp_7_25_port, 
      P_tmp_7_24_port, P_tmp_7_23_port, P_tmp_7_22_port, P_tmp_7_21_port, 
      P_tmp_7_20_port, P_tmp_7_19_port, P_tmp_7_18_port, P_tmp_7_17_port, 
      P_tmp_7_16_port, P_tmp_7_15_port, P_tmp_7_14_port, P_tmp_7_13_port, 
      P_tmp_7_12_port, P_tmp_7_11_port, P_tmp_7_10_port, P_tmp_7_9_port, 
      P_tmp_7_8_port, P_tmp_7_7_port, P_tmp_7_6_port, P_tmp_7_5_port, 
      P_tmp_7_4_port, P_tmp_7_3_port, P_tmp_7_2_port, P_tmp_7_1_port, 
      P_tmp_7_0_port, P_tmp_8_63_port, P_tmp_8_62_port, P_tmp_8_61_port, 
      P_tmp_8_60_port, P_tmp_8_59_port, P_tmp_8_58_port, P_tmp_8_57_port, 
      P_tmp_8_56_port, P_tmp_8_55_port, P_tmp_8_54_port, P_tmp_8_53_port, 
      P_tmp_8_52_port, P_tmp_8_51_port, P_tmp_8_50_port, P_tmp_8_49_port, 
      P_tmp_8_48_port, P_tmp_8_47_port, P_tmp_8_46_port, P_tmp_8_45_port, 
      P_tmp_8_44_port, P_tmp_8_43_port, P_tmp_8_42_port, P_tmp_8_41_port, 
      P_tmp_8_40_port, P_tmp_8_39_port, P_tmp_8_38_port, P_tmp_8_37_port, 
      P_tmp_8_36_port, P_tmp_8_35_port, P_tmp_8_34_port, P_tmp_8_33_port, 
      P_tmp_8_32_port, P_tmp_8_31_port, P_tmp_8_30_port, P_tmp_8_29_port, 
      P_tmp_8_28_port, P_tmp_8_27_port, P_tmp_8_26_port, P_tmp_8_25_port, 
      P_tmp_8_24_port, P_tmp_8_23_port, P_tmp_8_22_port, P_tmp_8_21_port, 
      P_tmp_8_20_port, P_tmp_8_19_port, P_tmp_8_18_port, P_tmp_8_17_port, 
      P_tmp_8_16_port, P_tmp_8_15_port, P_tmp_8_14_port, P_tmp_8_13_port, 
      P_tmp_8_12_port, P_tmp_8_11_port, P_tmp_8_10_port, P_tmp_8_9_port, 
      P_tmp_8_8_port, P_tmp_8_7_port, P_tmp_8_6_port, P_tmp_8_5_port, 
      P_tmp_8_4_port, P_tmp_8_3_port, P_tmp_8_2_port, P_tmp_8_1_port, 
      P_tmp_8_0_port, P_tmp_9_63_port, P_tmp_9_62_port, P_tmp_9_61_port, 
      P_tmp_9_60_port, P_tmp_9_59_port, P_tmp_9_58_port, P_tmp_9_57_port, 
      P_tmp_9_56_port, P_tmp_9_55_port, P_tmp_9_54_port, P_tmp_9_53_port, 
      P_tmp_9_52_port, P_tmp_9_51_port, P_tmp_9_50_port, P_tmp_9_49_port, 
      P_tmp_9_48_port, P_tmp_9_47_port, P_tmp_9_46_port, P_tmp_9_45_port, 
      P_tmp_9_44_port, P_tmp_9_43_port, P_tmp_9_42_port, P_tmp_9_41_port, 
      P_tmp_9_40_port, P_tmp_9_39_port, P_tmp_9_38_port, P_tmp_9_37_port, 
      P_tmp_9_36_port, P_tmp_9_35_port, P_tmp_9_34_port, P_tmp_9_33_port, 
      P_tmp_9_32_port, P_tmp_9_31_port, P_tmp_9_30_port, P_tmp_9_29_port, 
      P_tmp_9_28_port, P_tmp_9_27_port, P_tmp_9_26_port, P_tmp_9_25_port, 
      P_tmp_9_24_port, P_tmp_9_23_port, P_tmp_9_22_port, P_tmp_9_21_port, 
      P_tmp_9_20_port, P_tmp_9_19_port, P_tmp_9_18_port, P_tmp_9_17_port, 
      P_tmp_9_16_port, P_tmp_9_15_port, P_tmp_9_14_port, P_tmp_9_13_port, 
      P_tmp_9_12_port, P_tmp_9_11_port, P_tmp_9_10_port, P_tmp_9_9_port, 
      P_tmp_9_8_port, P_tmp_9_7_port, P_tmp_9_6_port, P_tmp_9_5_port, 
      P_tmp_9_4_port, P_tmp_9_3_port, P_tmp_9_2_port, P_tmp_9_1_port, 
      P_tmp_9_0_port, P_tmp_10_63_port, P_tmp_10_62_port, P_tmp_10_61_port, 
      P_tmp_10_60_port, P_tmp_10_59_port, P_tmp_10_58_port, P_tmp_10_57_port, 
      P_tmp_10_56_port, P_tmp_10_55_port, P_tmp_10_54_port, P_tmp_10_53_port, 
      P_tmp_10_52_port, P_tmp_10_51_port, P_tmp_10_50_port, P_tmp_10_49_port, 
      P_tmp_10_48_port, P_tmp_10_47_port, P_tmp_10_46_port, P_tmp_10_45_port, 
      P_tmp_10_44_port, P_tmp_10_43_port, P_tmp_10_42_port, P_tmp_10_41_port, 
      P_tmp_10_40_port, P_tmp_10_39_port, P_tmp_10_38_port, P_tmp_10_37_port, 
      P_tmp_10_36_port, P_tmp_10_35_port, P_tmp_10_34_port, P_tmp_10_33_port, 
      P_tmp_10_32_port, P_tmp_10_31_port, P_tmp_10_30_port, P_tmp_10_29_port, 
      P_tmp_10_28_port, P_tmp_10_27_port, P_tmp_10_26_port, P_tmp_10_25_port, 
      P_tmp_10_24_port, P_tmp_10_23_port, P_tmp_10_22_port, P_tmp_10_21_port, 
      P_tmp_10_20_port, P_tmp_10_19_port, P_tmp_10_18_port, P_tmp_10_17_port, 
      P_tmp_10_16_port, P_tmp_10_15_port, P_tmp_10_14_port, P_tmp_10_13_port, 
      P_tmp_10_12_port, P_tmp_10_11_port, P_tmp_10_10_port, P_tmp_10_9_port, 
      P_tmp_10_8_port, P_tmp_10_7_port, P_tmp_10_6_port, P_tmp_10_5_port, 
      P_tmp_10_4_port, P_tmp_10_3_port, P_tmp_10_2_port, P_tmp_10_1_port, 
      P_tmp_10_0_port, P_tmp_11_63_port, P_tmp_11_62_port, P_tmp_11_61_port, 
      P_tmp_11_60_port, P_tmp_11_59_port, P_tmp_11_58_port, P_tmp_11_57_port, 
      P_tmp_11_56_port, P_tmp_11_55_port, P_tmp_11_54_port, P_tmp_11_53_port, 
      P_tmp_11_52_port, P_tmp_11_51_port, P_tmp_11_50_port, P_tmp_11_49_port, 
      P_tmp_11_48_port, P_tmp_11_47_port, P_tmp_11_46_port, P_tmp_11_45_port, 
      P_tmp_11_44_port, P_tmp_11_43_port, P_tmp_11_42_port, P_tmp_11_41_port, 
      P_tmp_11_40_port, P_tmp_11_39_port, P_tmp_11_38_port, P_tmp_11_37_port, 
      P_tmp_11_36_port, P_tmp_11_35_port, P_tmp_11_34_port, P_tmp_11_33_port, 
      P_tmp_11_32_port, P_tmp_11_31_port, P_tmp_11_30_port, P_tmp_11_29_port, 
      P_tmp_11_28_port, P_tmp_11_27_port, P_tmp_11_26_port, P_tmp_11_25_port, 
      P_tmp_11_24_port, P_tmp_11_23_port, P_tmp_11_22_port, P_tmp_11_21_port, 
      P_tmp_11_20_port, P_tmp_11_19_port, P_tmp_11_18_port, P_tmp_11_17_port, 
      P_tmp_11_16_port, P_tmp_11_15_port, P_tmp_11_14_port, P_tmp_11_13_port, 
      P_tmp_11_12_port, P_tmp_11_11_port, P_tmp_11_10_port, P_tmp_11_9_port, 
      P_tmp_11_8_port, P_tmp_11_7_port, P_tmp_11_6_port, P_tmp_11_5_port, 
      P_tmp_11_4_port, P_tmp_11_3_port, P_tmp_11_2_port, P_tmp_11_1_port, 
      P_tmp_11_0_port, P_tmp_12_63_port, P_tmp_12_62_port, P_tmp_12_61_port, 
      P_tmp_12_60_port, P_tmp_12_59_port, P_tmp_12_58_port, P_tmp_12_57_port, 
      P_tmp_12_56_port, P_tmp_12_55_port, P_tmp_12_54_port, P_tmp_12_53_port, 
      P_tmp_12_52_port, P_tmp_12_51_port, P_tmp_12_50_port, P_tmp_12_49_port, 
      P_tmp_12_48_port, P_tmp_12_47_port, P_tmp_12_46_port, P_tmp_12_45_port, 
      P_tmp_12_44_port, P_tmp_12_43_port, P_tmp_12_42_port, P_tmp_12_41_port, 
      P_tmp_12_40_port, P_tmp_12_39_port, P_tmp_12_38_port, P_tmp_12_37_port, 
      P_tmp_12_36_port, P_tmp_12_35_port, P_tmp_12_34_port, P_tmp_12_33_port, 
      P_tmp_12_32_port, P_tmp_12_31_port, P_tmp_12_30_port, P_tmp_12_29_port, 
      P_tmp_12_28_port, P_tmp_12_27_port, P_tmp_12_26_port, P_tmp_12_25_port, 
      P_tmp_12_24_port, P_tmp_12_23_port, P_tmp_12_22_port, P_tmp_12_21_port, 
      P_tmp_12_20_port, P_tmp_12_19_port, P_tmp_12_18_port, P_tmp_12_17_port, 
      P_tmp_12_16_port, P_tmp_12_15_port, P_tmp_12_14_port, P_tmp_12_13_port, 
      P_tmp_12_12_port, P_tmp_12_11_port, P_tmp_12_10_port, P_tmp_12_9_port, 
      P_tmp_12_8_port, P_tmp_12_7_port, P_tmp_12_6_port, P_tmp_12_5_port, 
      P_tmp_12_4_port, P_tmp_12_3_port, P_tmp_12_2_port, P_tmp_12_1_port, 
      P_tmp_12_0_port, P_tmp_13_63_port, P_tmp_13_62_port, P_tmp_13_61_port, 
      P_tmp_13_60_port, P_tmp_13_59_port, P_tmp_13_58_port, P_tmp_13_57_port, 
      P_tmp_13_56_port, P_tmp_13_55_port, P_tmp_13_54_port, P_tmp_13_53_port, 
      P_tmp_13_52_port, P_tmp_13_51_port, P_tmp_13_50_port, P_tmp_13_49_port, 
      P_tmp_13_48_port, P_tmp_13_47_port, P_tmp_13_46_port, P_tmp_13_45_port, 
      P_tmp_13_44_port, P_tmp_13_43_port, P_tmp_13_42_port, P_tmp_13_41_port, 
      P_tmp_13_40_port, P_tmp_13_39_port, P_tmp_13_38_port, P_tmp_13_37_port, 
      P_tmp_13_36_port, P_tmp_13_35_port, P_tmp_13_34_port, P_tmp_13_33_port, 
      P_tmp_13_32_port, P_tmp_13_31_port, P_tmp_13_30_port, P_tmp_13_29_port, 
      P_tmp_13_28_port, P_tmp_13_27_port, P_tmp_13_26_port, P_tmp_13_25_port, 
      P_tmp_13_24_port, P_tmp_13_23_port, P_tmp_13_22_port, P_tmp_13_21_port, 
      P_tmp_13_20_port, P_tmp_13_19_port, P_tmp_13_18_port, P_tmp_13_17_port, 
      P_tmp_13_16_port, P_tmp_13_15_port, P_tmp_13_14_port, P_tmp_13_13_port, 
      P_tmp_13_12_port, P_tmp_13_11_port, P_tmp_13_10_port, P_tmp_13_9_port, 
      P_tmp_13_8_port, P_tmp_13_7_port, P_tmp_13_6_port, P_tmp_13_5_port, 
      P_tmp_13_4_port, P_tmp_13_3_port, P_tmp_13_2_port, P_tmp_13_1_port, 
      P_tmp_13_0_port, P_tmp_14_63_port, P_tmp_14_62_port, P_tmp_14_61_port, 
      P_tmp_14_60_port, P_tmp_14_59_port, P_tmp_14_58_port, P_tmp_14_57_port, 
      P_tmp_14_56_port, P_tmp_14_55_port, P_tmp_14_54_port, P_tmp_14_53_port, 
      P_tmp_14_52_port, P_tmp_14_51_port, P_tmp_14_50_port, P_tmp_14_49_port, 
      P_tmp_14_48_port, P_tmp_14_47_port, P_tmp_14_46_port, P_tmp_14_45_port, 
      P_tmp_14_44_port, P_tmp_14_43_port, P_tmp_14_42_port, P_tmp_14_41_port, 
      P_tmp_14_40_port, P_tmp_14_39_port, P_tmp_14_38_port, P_tmp_14_37_port, 
      P_tmp_14_36_port, P_tmp_14_35_port, P_tmp_14_34_port, P_tmp_14_33_port, 
      P_tmp_14_32_port, P_tmp_14_31_port, P_tmp_14_30_port, P_tmp_14_29_port, 
      P_tmp_14_28_port, P_tmp_14_27_port, P_tmp_14_26_port, P_tmp_14_25_port, 
      P_tmp_14_24_port, P_tmp_14_23_port, P_tmp_14_22_port, P_tmp_14_21_port, 
      P_tmp_14_20_port, P_tmp_14_19_port, P_tmp_14_18_port, P_tmp_14_17_port, 
      P_tmp_14_16_port, P_tmp_14_15_port, P_tmp_14_14_port, P_tmp_14_13_port, 
      P_tmp_14_12_port, P_tmp_14_11_port, P_tmp_14_10_port, P_tmp_14_9_port, 
      P_tmp_14_8_port, P_tmp_14_7_port, P_tmp_14_6_port, P_tmp_14_5_port, 
      P_tmp_14_4_port, P_tmp_14_3_port, P_tmp_14_2_port, P_tmp_14_1_port, 
      P_tmp_14_0_port, n127, net15393, net15391, net15399, net15397, net15405, 
      net15403, net15411, net15409, net15417, net15415, net15423, net15421, 
      net15429, net15427, net15435, net15433, net15441, net15439, net15447, 
      net15445, net15453, net15451, net15457, net15465, net15463, net15471, 
      net15469, net15477, net15475, net15483, net15481, net15489, net15487, 
      net15495, net15493, net15525, net15523, net15535, net15533, net15837, 
      net17026, net17038, net17036, net17729, net18006, net18009, net18016, 
      net18025, net18732, net25715, net98228, net17616, net17614, net17613, 
      n129, n128, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n_1060,
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   A_pos_shifted_by1_1_0_port <= '0';
   A_pos_shifted_by2_1_0_port <= '0';
   A_pos_shifted_by2_1_1_port <= '0';
   A_pos_shifted_by1_2_0_port <= '0';
   A_pos_shifted_by2_2_0_port <= '0';
   A_pos_shifted_by2_2_1_port <= '0';
   A_pos_shifted_by1_3_0_port <= '0';
   A_pos_shifted_by2_3_0_port <= '0';
   A_pos_shifted_by2_3_1_port <= '0';
   A_pos_shifted_by1_4_0_port <= '0';
   A_pos_shifted_by2_4_0_port <= '0';
   A_pos_shifted_by2_4_1_port <= '0';
   A_pos_shifted_by1_5_0_port <= '0';
   A_pos_shifted_by2_5_0_port <= '0';
   A_pos_shifted_by2_5_1_port <= '0';
   A_pos_shifted_by1_6_0_port <= '0';
   A_pos_shifted_by2_6_0_port <= '0';
   A_pos_shifted_by2_6_1_port <= '0';
   A_pos_shifted_by1_7_0_port <= '0';
   A_pos_shifted_by2_7_0_port <= '0';
   A_pos_shifted_by2_7_1_port <= '0';
   A_pos_shifted_by1_8_0_port <= '0';
   A_pos_shifted_by2_8_0_port <= '0';
   A_pos_shifted_by2_8_1_port <= '0';
   A_pos_shifted_by1_9_0_port <= '0';
   A_pos_shifted_by2_9_0_port <= '0';
   A_pos_shifted_by2_9_1_port <= '0';
   A_pos_shifted_by1_10_0_port <= '0';
   A_pos_shifted_by2_10_0_port <= '0';
   A_pos_shifted_by2_10_1_port <= '0';
   A_pos_shifted_by1_11_0_port <= '0';
   A_pos_shifted_by2_11_0_port <= '0';
   A_pos_shifted_by2_11_1_port <= '0';
   A_pos_shifted_by1_12_0_port <= '0';
   A_pos_shifted_by2_12_0_port <= '0';
   A_pos_shifted_by2_12_1_port <= '0';
   A_pos_shifted_by1_13_0_port <= '0';
   A_pos_shifted_by2_13_0_port <= '0';
   A_pos_shifted_by2_13_1_port <= '0';
   A_pos_shifted_by1_14_0_port <= '0';
   A_pos_shifted_by2_14_0_port <= '0';
   A_pos_shifted_by2_14_1_port <= '0';
   A_pos_shifted_by1_15_0_port <= '0';
   A_neg_shifted_by1_0_0_port <= '0';
   A_neg_shifted_by2_0_0_port <= '0';
   A_neg_shifted_by2_0_1_port <= '0';
   A_neg_shifted_by1_1_0_port <= '0';
   A_neg_shifted_by2_1_0_port <= '0';
   A_neg_shifted_by2_1_1_port <= '0';
   A_neg_shifted_by1_2_0_port <= '0';
   A_neg_shifted_by2_2_0_port <= '0';
   A_neg_shifted_by2_2_1_port <= '0';
   A_neg_shifted_by1_3_0_port <= '0';
   A_neg_shifted_by2_3_0_port <= '0';
   A_neg_shifted_by2_3_1_port <= '0';
   A_neg_shifted_by1_4_0_port <= '0';
   A_neg_shifted_by2_4_0_port <= '0';
   A_neg_shifted_by2_4_1_port <= '0';
   A_neg_shifted_by1_5_0_port <= '0';
   A_neg_shifted_by2_5_0_port <= '0';
   A_neg_shifted_by2_5_1_port <= '0';
   A_neg_shifted_by1_6_0_port <= '0';
   A_neg_shifted_by2_6_0_port <= '0';
   A_neg_shifted_by2_6_1_port <= '0';
   A_neg_shifted_by1_7_0_port <= '0';
   A_neg_shifted_by2_7_0_port <= '0';
   A_neg_shifted_by2_7_1_port <= '0';
   A_neg_shifted_by1_8_0_port <= '0';
   A_neg_shifted_by2_8_0_port <= '0';
   A_neg_shifted_by2_8_1_port <= '0';
   A_neg_shifted_by1_9_0_port <= '0';
   A_neg_shifted_by2_9_0_port <= '0';
   A_neg_shifted_by2_9_1_port <= '0';
   A_neg_shifted_by1_10_0_port <= '0';
   A_neg_shifted_by2_10_0_port <= '0';
   A_neg_shifted_by2_10_1_port <= '0';
   A_neg_shifted_by1_11_0_port <= '0';
   A_neg_shifted_by2_11_0_port <= '0';
   A_neg_shifted_by2_11_1_port <= '0';
   A_neg_shifted_by1_12_0_port <= '0';
   A_neg_shifted_by2_12_0_port <= '0';
   A_neg_shifted_by2_12_1_port <= '0';
   A_neg_shifted_by1_13_0_port <= '0';
   A_neg_shifted_by2_13_0_port <= '0';
   A_neg_shifted_by2_13_1_port <= '0';
   A_neg_shifted_by1_14_0_port <= '0';
   A_neg_shifted_by2_14_0_port <= '0';
   A_neg_shifted_by2_14_1_port <= '0';
   A_neg_shifted_by1_15_0_port <= '0';
   A_pos_shifted_by1_0_0_port <= '0';
   A_pos_shifted_by2_0_0_port <= '0';
   A_pos_shifted_by2_0_1_port <= '0';
   Booth_Encoder0_0 : Booth_Encoder_0 port map( B(2) => n193, B(1) => B(0), 
                           B(0) => X_Logic0_port, OUT_TO_MUX(2) => 
                           selection_signal_0_2_port, OUT_TO_MUX(1) => 
                           selection_signal_0_1_port, OUT_TO_MUX(0) => 
                           selection_signal_0_0_port);
   Booth_Encoderi_1 : Booth_Encoder_15 port map( B(2) => B(3), B(1) => B(2), 
                           B(0) => B(1), OUT_TO_MUX(2) => 
                           selection_signal_1_2_port, OUT_TO_MUX(1) => 
                           selection_signal_1_1_port, OUT_TO_MUX(0) => 
                           selection_signal_1_0_port);
   Booth_Encoderi_2 : Booth_Encoder_14 port map( B(2) => B(5), B(1) => B(4), 
                           B(0) => B(3), OUT_TO_MUX(2) => 
                           selection_signal_2_2_port, OUT_TO_MUX(1) => 
                           selection_signal_2_1_port, OUT_TO_MUX(0) => 
                           selection_signal_2_0_port);
   Booth_Encoderi_3 : Booth_Encoder_13 port map( B(2) => B(7), B(1) => B(6), 
                           B(0) => B(5), OUT_TO_MUX(2) => 
                           selection_signal_3_2_port, OUT_TO_MUX(1) => 
                           selection_signal_3_1_port, OUT_TO_MUX(0) => 
                           selection_signal_3_0_port);
   Booth_Encoderi_4 : Booth_Encoder_12 port map( B(2) => B(9), B(1) => B(8), 
                           B(0) => B(7), OUT_TO_MUX(2) => 
                           selection_signal_4_2_port, OUT_TO_MUX(1) => 
                           selection_signal_4_1_port, OUT_TO_MUX(0) => 
                           selection_signal_4_0_port);
   Booth_Encoderi_5 : Booth_Encoder_11 port map( B(2) => B(11), B(1) => B(10), 
                           B(0) => B(9), OUT_TO_MUX(2) => 
                           selection_signal_5_2_port, OUT_TO_MUX(1) => 
                           selection_signal_5_1_port, OUT_TO_MUX(0) => 
                           selection_signal_5_0_port);
   Booth_Encoderi_6 : Booth_Encoder_10 port map( B(2) => B(13), B(1) => B(12), 
                           B(0) => B(11), OUT_TO_MUX(2) => 
                           selection_signal_6_2_port, OUT_TO_MUX(1) => 
                           selection_signal_6_1_port, OUT_TO_MUX(0) => 
                           selection_signal_6_0_port);
   Booth_Encoderi_7 : Booth_Encoder_9 port map( B(2) => B(15), B(1) => B(14), 
                           B(0) => B(13), OUT_TO_MUX(2) => 
                           selection_signal_7_2_port, OUT_TO_MUX(1) => 
                           selection_signal_7_1_port, OUT_TO_MUX(0) => 
                           selection_signal_7_0_port);
   Booth_Encoderi_8 : Booth_Encoder_8 port map( B(2) => B(17), B(1) => B(16), 
                           B(0) => B(15), OUT_TO_MUX(2) => 
                           selection_signal_8_2_port, OUT_TO_MUX(1) => 
                           selection_signal_8_1_port, OUT_TO_MUX(0) => 
                           selection_signal_8_0_port);
   Booth_Encoderi_9 : Booth_Encoder_7 port map( B(2) => B(19), B(1) => B(18), 
                           B(0) => B(17), OUT_TO_MUX(2) => 
                           selection_signal_9_2_port, OUT_TO_MUX(1) => 
                           selection_signal_9_1_port, OUT_TO_MUX(0) => 
                           selection_signal_9_0_port);
   Booth_Encoderi_10 : Booth_Encoder_6 port map( B(2) => B(21), B(1) => B(20), 
                           B(0) => B(19), OUT_TO_MUX(2) => 
                           selection_signal_10_2_port, OUT_TO_MUX(1) => 
                           selection_signal_10_1_port, OUT_TO_MUX(0) => 
                           selection_signal_10_0_port);
   Booth_Encoderi_11 : Booth_Encoder_5 port map( B(2) => B(23), B(1) => B(22), 
                           B(0) => B(21), OUT_TO_MUX(2) => 
                           selection_signal_11_2_port, OUT_TO_MUX(1) => 
                           selection_signal_11_1_port, OUT_TO_MUX(0) => 
                           selection_signal_11_0_port);
   Booth_Encoderi_12 : Booth_Encoder_4 port map( B(2) => B(25), B(1) => B(24), 
                           B(0) => B(23), OUT_TO_MUX(2) => 
                           selection_signal_12_2_port, OUT_TO_MUX(1) => 
                           selection_signal_12_1_port, OUT_TO_MUX(0) => 
                           selection_signal_12_0_port);
   Booth_Encoderi_13 : Booth_Encoder_3 port map( B(2) => B(27), B(1) => B(26), 
                           B(0) => B(25), OUT_TO_MUX(2) => 
                           selection_signal_13_2_port, OUT_TO_MUX(1) => 
                           selection_signal_13_1_port, OUT_TO_MUX(0) => 
                           selection_signal_13_0_port);
   Booth_Encoderi_14 : Booth_Encoder_2 port map( B(2) => B(29), B(1) => B(28), 
                           B(0) => B(27), OUT_TO_MUX(2) => 
                           selection_signal_14_2_port, OUT_TO_MUX(1) => 
                           selection_signal_14_1_port, OUT_TO_MUX(0) => 
                           selection_signal_14_0_port);
   Booth_Encoderi_15 : Booth_Encoder_1 port map( B(2) => B(31), B(1) => B(30), 
                           B(0) => B(29), OUT_TO_MUX(2) => 
                           selection_signal_15_2_port, OUT_TO_MUX(1) => 
                           selection_signal_15_1_port, OUT_TO_MUX(0) => 
                           selection_signal_15_0_port);
   SHIFTER0_0 : Shifter_NBIT64_0 port map( TO_SHIFT(63) => n233, TO_SHIFT(62) 
                           => n233, TO_SHIFT(61) => n233, TO_SHIFT(60) => n232,
                           TO_SHIFT(59) => n232, TO_SHIFT(58) => n233, 
                           TO_SHIFT(57) => n233, TO_SHIFT(56) => n230, 
                           TO_SHIFT(55) => n230, TO_SHIFT(54) => n230, 
                           TO_SHIFT(53) => n230, TO_SHIFT(52) => n231, 
                           TO_SHIFT(51) => n232, TO_SHIFT(50) => n232, 
                           TO_SHIFT(49) => n231, TO_SHIFT(48) => n230, 
                           TO_SHIFT(47) => n230, TO_SHIFT(46) => n233, 
                           TO_SHIFT(45) => n233, TO_SHIFT(44) => n230, 
                           TO_SHIFT(43) => n230, TO_SHIFT(42) => n230, 
                           TO_SHIFT(41) => n232, TO_SHIFT(40) => n230, 
                           TO_SHIFT(39) => n232, TO_SHIFT(38) => n232, 
                           TO_SHIFT(37) => n232, TO_SHIFT(36) => n232, 
                           TO_SHIFT(35) => n232, TO_SHIFT(34) => n232, 
                           TO_SHIFT(33) => n231, TO_SHIFT(32) => n230, 
                           TO_SHIFT(31) => n231, TO_SHIFT(30) => n228, 
                           TO_SHIFT(29) => n226, TO_SHIFT(28) => n224, 
                           TO_SHIFT(27) => n222, TO_SHIFT(26) => n220, 
                           TO_SHIFT(25) => n218, TO_SHIFT(24) => n216, 
                           TO_SHIFT(23) => net15391, TO_SHIFT(22) => net15397, 
                           TO_SHIFT(21) => net15403, TO_SHIFT(20) => net15409, 
                           TO_SHIFT(19) => net15415, TO_SHIFT(18) => net15421, 
                           TO_SHIFT(17) => net15427, TO_SHIFT(16) => net15433, 
                           TO_SHIFT(15) => net15439, TO_SHIFT(14) => net15445, 
                           TO_SHIFT(13) => net15451, TO_SHIFT(12) => net15457, 
                           TO_SHIFT(11) => net15463, TO_SHIFT(10) => net15469, 
                           TO_SHIFT(9) => net15475, TO_SHIFT(8) => net15481, 
                           TO_SHIFT(7) => net15487, TO_SHIFT(6) => net15493, 
                           TO_SHIFT(5) => n214, TO_SHIFT(4) => n212, 
                           TO_SHIFT(3) => n210, TO_SHIFT(2) => n208, 
                           TO_SHIFT(1) => net15523, TO_SHIFT(0) => net15533, 
                           RESULT(127) => A_pos_shifted_by2_0_63_port, 
                           RESULT(126) => A_pos_shifted_by2_0_62_port, 
                           RESULT(125) => A_pos_shifted_by2_0_61_port, 
                           RESULT(124) => A_pos_shifted_by2_0_60_port, 
                           RESULT(123) => A_pos_shifted_by2_0_59_port, 
                           RESULT(122) => A_pos_shifted_by2_0_58_port, 
                           RESULT(121) => A_pos_shifted_by2_0_57_port, 
                           RESULT(120) => A_pos_shifted_by2_0_56_port, 
                           RESULT(119) => A_pos_shifted_by2_0_55_port, 
                           RESULT(118) => A_pos_shifted_by2_0_54_port, 
                           RESULT(117) => A_pos_shifted_by2_0_53_port, 
                           RESULT(116) => A_pos_shifted_by2_0_52_port, 
                           RESULT(115) => A_pos_shifted_by2_0_51_port, 
                           RESULT(114) => A_pos_shifted_by2_0_50_port, 
                           RESULT(113) => A_pos_shifted_by2_0_49_port, 
                           RESULT(112) => A_pos_shifted_by2_0_48_port, 
                           RESULT(111) => A_pos_shifted_by2_0_47_port, 
                           RESULT(110) => A_pos_shifted_by2_0_46_port, 
                           RESULT(109) => A_pos_shifted_by2_0_45_port, 
                           RESULT(108) => A_pos_shifted_by2_0_44_port, 
                           RESULT(107) => A_pos_shifted_by2_0_43_port, 
                           RESULT(106) => A_pos_shifted_by2_0_42_port, 
                           RESULT(105) => A_pos_shifted_by2_0_41_port, 
                           RESULT(104) => A_pos_shifted_by2_0_40_port, 
                           RESULT(103) => A_pos_shifted_by2_0_39_port, 
                           RESULT(102) => A_pos_shifted_by2_0_38_port, 
                           RESULT(101) => A_pos_shifted_by2_0_37_port, 
                           RESULT(100) => A_pos_shifted_by2_0_36_port, 
                           RESULT(99) => A_pos_shifted_by2_0_35_port, 
                           RESULT(98) => A_pos_shifted_by2_0_34_port, 
                           RESULT(97) => A_pos_shifted_by2_0_33_port, 
                           RESULT(96) => A_pos_shifted_by2_0_32_port, 
                           RESULT(95) => A_pos_shifted_by2_0_31_port, 
                           RESULT(94) => A_pos_shifted_by2_0_30_port, 
                           RESULT(93) => A_pos_shifted_by2_0_29_port, 
                           RESULT(92) => A_pos_shifted_by2_0_28_port, 
                           RESULT(91) => A_pos_shifted_by2_0_27_port, 
                           RESULT(90) => A_pos_shifted_by2_0_26_port, 
                           RESULT(89) => A_pos_shifted_by2_0_25_port, 
                           RESULT(88) => A_pos_shifted_by2_0_24_port, 
                           RESULT(87) => A_pos_shifted_by2_0_23_port, 
                           RESULT(86) => A_pos_shifted_by2_0_22_port, 
                           RESULT(85) => A_pos_shifted_by2_0_21_port, 
                           RESULT(84) => A_pos_shifted_by2_0_20_port, 
                           RESULT(83) => A_pos_shifted_by2_0_19_port, 
                           RESULT(82) => A_pos_shifted_by2_0_18_port, 
                           RESULT(81) => A_pos_shifted_by2_0_17_port, 
                           RESULT(80) => A_pos_shifted_by2_0_16_port, 
                           RESULT(79) => A_pos_shifted_by2_0_15_port, 
                           RESULT(78) => A_pos_shifted_by2_0_14_port, 
                           RESULT(77) => A_pos_shifted_by2_0_13_port, 
                           RESULT(76) => A_pos_shifted_by2_0_12_port, 
                           RESULT(75) => A_pos_shifted_by2_0_11_port, 
                           RESULT(74) => A_pos_shifted_by2_0_10_port, 
                           RESULT(73) => A_pos_shifted_by2_0_9_port, RESULT(72)
                           => A_pos_shifted_by2_0_8_port, RESULT(71) => 
                           A_pos_shifted_by2_0_7_port, RESULT(70) => 
                           A_pos_shifted_by2_0_6_port, RESULT(69) => 
                           A_pos_shifted_by2_0_5_port, RESULT(68) => 
                           A_pos_shifted_by2_0_4_port, RESULT(67) => 
                           A_pos_shifted_by2_0_3_port, RESULT(66) => 
                           A_pos_shifted_by2_0_2_port, RESULT(65) => n_1060, 
                           RESULT(64) => n_1061, RESULT(63) => 
                           A_pos_shifted_by1_0_63_port, RESULT(62) => 
                           A_pos_shifted_by1_0_62_port, RESULT(61) => 
                           A_pos_shifted_by1_0_61_port, RESULT(60) => 
                           A_pos_shifted_by1_0_60_port, RESULT(59) => 
                           A_pos_shifted_by1_0_59_port, RESULT(58) => 
                           A_pos_shifted_by1_0_58_port, RESULT(57) => 
                           A_pos_shifted_by1_0_57_port, RESULT(56) => 
                           A_pos_shifted_by1_0_56_port, RESULT(55) => 
                           A_pos_shifted_by1_0_55_port, RESULT(54) => 
                           A_pos_shifted_by1_0_54_port, RESULT(53) => 
                           A_pos_shifted_by1_0_53_port, RESULT(52) => 
                           A_pos_shifted_by1_0_52_port, RESULT(51) => 
                           A_pos_shifted_by1_0_51_port, RESULT(50) => 
                           A_pos_shifted_by1_0_50_port, RESULT(49) => 
                           A_pos_shifted_by1_0_49_port, RESULT(48) => 
                           A_pos_shifted_by1_0_48_port, RESULT(47) => 
                           A_pos_shifted_by1_0_47_port, RESULT(46) => 
                           A_pos_shifted_by1_0_46_port, RESULT(45) => 
                           A_pos_shifted_by1_0_45_port, RESULT(44) => 
                           A_pos_shifted_by1_0_44_port, RESULT(43) => 
                           A_pos_shifted_by1_0_43_port, RESULT(42) => 
                           A_pos_shifted_by1_0_42_port, RESULT(41) => 
                           A_pos_shifted_by1_0_41_port, RESULT(40) => 
                           A_pos_shifted_by1_0_40_port, RESULT(39) => 
                           A_pos_shifted_by1_0_39_port, RESULT(38) => 
                           A_pos_shifted_by1_0_38_port, RESULT(37) => 
                           A_pos_shifted_by1_0_37_port, RESULT(36) => 
                           A_pos_shifted_by1_0_36_port, RESULT(35) => 
                           A_pos_shifted_by1_0_35_port, RESULT(34) => 
                           A_pos_shifted_by1_0_34_port, RESULT(33) => 
                           A_pos_shifted_by1_0_33_port, RESULT(32) => 
                           A_pos_shifted_by1_0_32_port, RESULT(31) => 
                           A_pos_shifted_by1_0_31_port, RESULT(30) => 
                           A_pos_shifted_by1_0_30_port, RESULT(29) => 
                           A_pos_shifted_by1_0_29_port, RESULT(28) => 
                           A_pos_shifted_by1_0_28_port, RESULT(27) => 
                           A_pos_shifted_by1_0_27_port, RESULT(26) => 
                           A_pos_shifted_by1_0_26_port, RESULT(25) => 
                           A_pos_shifted_by1_0_25_port, RESULT(24) => 
                           A_pos_shifted_by1_0_24_port, RESULT(23) => 
                           A_pos_shifted_by1_0_23_port, RESULT(22) => 
                           A_pos_shifted_by1_0_22_port, RESULT(21) => 
                           A_pos_shifted_by1_0_21_port, RESULT(20) => 
                           A_pos_shifted_by1_0_20_port, RESULT(19) => 
                           A_pos_shifted_by1_0_19_port, RESULT(18) => 
                           A_pos_shifted_by1_0_18_port, RESULT(17) => 
                           A_pos_shifted_by1_0_17_port, RESULT(16) => 
                           A_pos_shifted_by1_0_16_port, RESULT(15) => 
                           A_pos_shifted_by1_0_15_port, RESULT(14) => 
                           A_pos_shifted_by1_0_14_port, RESULT(13) => 
                           A_pos_shifted_by1_0_13_port, RESULT(12) => 
                           A_pos_shifted_by1_0_12_port, RESULT(11) => 
                           A_pos_shifted_by1_0_11_port, RESULT(10) => 
                           A_pos_shifted_by1_0_10_port, RESULT(9) => 
                           A_pos_shifted_by1_0_9_port, RESULT(8) => 
                           A_pos_shifted_by1_0_8_port, RESULT(7) => 
                           A_pos_shifted_by1_0_7_port, RESULT(6) => 
                           A_pos_shifted_by1_0_6_port, RESULT(5) => 
                           A_pos_shifted_by1_0_5_port, RESULT(4) => 
                           A_pos_shifted_by1_0_4_port, RESULT(3) => 
                           A_pos_shifted_by1_0_3_port, RESULT(2) => 
                           A_pos_shifted_by1_0_2_port, RESULT(1) => 
                           A_pos_shifted_by1_0_1_port, RESULT(0) => n_1062);
   SHIFTERi_1 : Shifter_NBIT64_31 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_0_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_0_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_0_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_0_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_0_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_0_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_0_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_0_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_0_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_0_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_0_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_0_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_0_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_0_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_0_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_0_48_port, TO_SHIFT(47) => n242, 
                           TO_SHIFT(46) => A_pos_shifted_by2_0_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_0_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_0_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_0_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_0_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_0_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_0_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_0_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_0_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_0_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_0_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_0_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_0_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_0_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_0_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_0_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_0_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_0_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_0_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_0_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_0_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_0_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_0_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_0_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_0_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_0_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_0_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_0_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_0_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_0_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_0_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_0_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_0_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_0_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_0_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_0_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_0_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_0_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_0_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_0_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_0_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_0_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_0_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_0_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_0_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_0_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_0_0_port, 
                           RESULT(127) => A_pos_shifted_by2_1_63_port, 
                           RESULT(126) => A_pos_shifted_by2_1_62_port, 
                           RESULT(125) => A_pos_shifted_by2_1_61_port, 
                           RESULT(124) => A_pos_shifted_by2_1_60_port, 
                           RESULT(123) => A_pos_shifted_by2_1_59_port, 
                           RESULT(122) => A_pos_shifted_by2_1_58_port, 
                           RESULT(121) => A_pos_shifted_by2_1_57_port, 
                           RESULT(120) => A_pos_shifted_by2_1_56_port, 
                           RESULT(119) => A_pos_shifted_by2_1_55_port, 
                           RESULT(118) => A_pos_shifted_by2_1_54_port, 
                           RESULT(117) => A_pos_shifted_by2_1_53_port, 
                           RESULT(116) => A_pos_shifted_by2_1_52_port, 
                           RESULT(115) => A_pos_shifted_by2_1_51_port, 
                           RESULT(114) => A_pos_shifted_by2_1_50_port, 
                           RESULT(113) => A_pos_shifted_by2_1_49_port, 
                           RESULT(112) => A_pos_shifted_by2_1_48_port, 
                           RESULT(111) => A_pos_shifted_by2_1_47_port, 
                           RESULT(110) => A_pos_shifted_by2_1_46_port, 
                           RESULT(109) => A_pos_shifted_by2_1_45_port, 
                           RESULT(108) => A_pos_shifted_by2_1_44_port, 
                           RESULT(107) => A_pos_shifted_by2_1_43_port, 
                           RESULT(106) => A_pos_shifted_by2_1_42_port, 
                           RESULT(105) => A_pos_shifted_by2_1_41_port, 
                           RESULT(104) => A_pos_shifted_by2_1_40_port, 
                           RESULT(103) => A_pos_shifted_by2_1_39_port, 
                           RESULT(102) => A_pos_shifted_by2_1_38_port, 
                           RESULT(101) => A_pos_shifted_by2_1_37_port, 
                           RESULT(100) => A_pos_shifted_by2_1_36_port, 
                           RESULT(99) => A_pos_shifted_by2_1_35_port, 
                           RESULT(98) => A_pos_shifted_by2_1_34_port, 
                           RESULT(97) => A_pos_shifted_by2_1_33_port, 
                           RESULT(96) => A_pos_shifted_by2_1_32_port, 
                           RESULT(95) => A_pos_shifted_by2_1_31_port, 
                           RESULT(94) => A_pos_shifted_by2_1_30_port, 
                           RESULT(93) => A_pos_shifted_by2_1_29_port, 
                           RESULT(92) => A_pos_shifted_by2_1_28_port, 
                           RESULT(91) => A_pos_shifted_by2_1_27_port, 
                           RESULT(90) => A_pos_shifted_by2_1_26_port, 
                           RESULT(89) => A_pos_shifted_by2_1_25_port, 
                           RESULT(88) => A_pos_shifted_by2_1_24_port, 
                           RESULT(87) => A_pos_shifted_by2_1_23_port, 
                           RESULT(86) => A_pos_shifted_by2_1_22_port, 
                           RESULT(85) => A_pos_shifted_by2_1_21_port, 
                           RESULT(84) => A_pos_shifted_by2_1_20_port, 
                           RESULT(83) => A_pos_shifted_by2_1_19_port, 
                           RESULT(82) => A_pos_shifted_by2_1_18_port, 
                           RESULT(81) => A_pos_shifted_by2_1_17_port, 
                           RESULT(80) => A_pos_shifted_by2_1_16_port, 
                           RESULT(79) => A_pos_shifted_by2_1_15_port, 
                           RESULT(78) => A_pos_shifted_by2_1_14_port, 
                           RESULT(77) => A_pos_shifted_by2_1_13_port, 
                           RESULT(76) => A_pos_shifted_by2_1_12_port, 
                           RESULT(75) => A_pos_shifted_by2_1_11_port, 
                           RESULT(74) => A_pos_shifted_by2_1_10_port, 
                           RESULT(73) => A_pos_shifted_by2_1_9_port, RESULT(72)
                           => A_pos_shifted_by2_1_8_port, RESULT(71) => 
                           A_pos_shifted_by2_1_7_port, RESULT(70) => 
                           A_pos_shifted_by2_1_6_port, RESULT(69) => 
                           A_pos_shifted_by2_1_5_port, RESULT(68) => 
                           A_pos_shifted_by2_1_4_port, RESULT(67) => 
                           A_pos_shifted_by2_1_3_port, RESULT(66) => 
                           A_pos_shifted_by2_1_2_port, RESULT(65) => n_1063, 
                           RESULT(64) => n_1064, RESULT(63) => 
                           A_pos_shifted_by1_1_63_port, RESULT(62) => 
                           A_pos_shifted_by1_1_62_port, RESULT(61) => 
                           A_pos_shifted_by1_1_61_port, RESULT(60) => 
                           A_pos_shifted_by1_1_60_port, RESULT(59) => 
                           A_pos_shifted_by1_1_59_port, RESULT(58) => 
                           A_pos_shifted_by1_1_58_port, RESULT(57) => 
                           A_pos_shifted_by1_1_57_port, RESULT(56) => 
                           A_pos_shifted_by1_1_56_port, RESULT(55) => 
                           A_pos_shifted_by1_1_55_port, RESULT(54) => 
                           A_pos_shifted_by1_1_54_port, RESULT(53) => 
                           A_pos_shifted_by1_1_53_port, RESULT(52) => 
                           A_pos_shifted_by1_1_52_port, RESULT(51) => 
                           A_pos_shifted_by1_1_51_port, RESULT(50) => 
                           A_pos_shifted_by1_1_50_port, RESULT(49) => 
                           A_pos_shifted_by1_1_49_port, RESULT(48) => 
                           A_pos_shifted_by1_1_48_port, RESULT(47) => 
                           A_pos_shifted_by1_1_47_port, RESULT(46) => 
                           A_pos_shifted_by1_1_46_port, RESULT(45) => 
                           A_pos_shifted_by1_1_45_port, RESULT(44) => 
                           A_pos_shifted_by1_1_44_port, RESULT(43) => 
                           A_pos_shifted_by1_1_43_port, RESULT(42) => 
                           A_pos_shifted_by1_1_42_port, RESULT(41) => 
                           A_pos_shifted_by1_1_41_port, RESULT(40) => 
                           A_pos_shifted_by1_1_40_port, RESULT(39) => 
                           A_pos_shifted_by1_1_39_port, RESULT(38) => 
                           A_pos_shifted_by1_1_38_port, RESULT(37) => 
                           A_pos_shifted_by1_1_37_port, RESULT(36) => 
                           A_pos_shifted_by1_1_36_port, RESULT(35) => 
                           A_pos_shifted_by1_1_35_port, RESULT(34) => 
                           A_pos_shifted_by1_1_34_port, RESULT(33) => 
                           A_pos_shifted_by1_1_33_port, RESULT(32) => 
                           A_pos_shifted_by1_1_32_port, RESULT(31) => 
                           A_pos_shifted_by1_1_31_port, RESULT(30) => 
                           A_pos_shifted_by1_1_30_port, RESULT(29) => 
                           A_pos_shifted_by1_1_29_port, RESULT(28) => 
                           A_pos_shifted_by1_1_28_port, RESULT(27) => 
                           A_pos_shifted_by1_1_27_port, RESULT(26) => 
                           A_pos_shifted_by1_1_26_port, RESULT(25) => 
                           A_pos_shifted_by1_1_25_port, RESULT(24) => 
                           A_pos_shifted_by1_1_24_port, RESULT(23) => 
                           A_pos_shifted_by1_1_23_port, RESULT(22) => 
                           A_pos_shifted_by1_1_22_port, RESULT(21) => 
                           A_pos_shifted_by1_1_21_port, RESULT(20) => 
                           A_pos_shifted_by1_1_20_port, RESULT(19) => 
                           A_pos_shifted_by1_1_19_port, RESULT(18) => 
                           A_pos_shifted_by1_1_18_port, RESULT(17) => 
                           A_pos_shifted_by1_1_17_port, RESULT(16) => 
                           A_pos_shifted_by1_1_16_port, RESULT(15) => 
                           A_pos_shifted_by1_1_15_port, RESULT(14) => 
                           A_pos_shifted_by1_1_14_port, RESULT(13) => 
                           A_pos_shifted_by1_1_13_port, RESULT(12) => 
                           A_pos_shifted_by1_1_12_port, RESULT(11) => 
                           A_pos_shifted_by1_1_11_port, RESULT(10) => 
                           A_pos_shifted_by1_1_10_port, RESULT(9) => 
                           A_pos_shifted_by1_1_9_port, RESULT(8) => 
                           A_pos_shifted_by1_1_8_port, RESULT(7) => 
                           A_pos_shifted_by1_1_7_port, RESULT(6) => 
                           A_pos_shifted_by1_1_6_port, RESULT(5) => 
                           A_pos_shifted_by1_1_5_port, RESULT(4) => 
                           A_pos_shifted_by1_1_4_port, RESULT(3) => 
                           A_pos_shifted_by1_1_3_port, RESULT(2) => 
                           A_pos_shifted_by1_1_2_port, RESULT(1) => 
                           A_pos_shifted_by1_1_1_port, RESULT(0) => n_1065);
   SHIFTERi_2 : Shifter_NBIT64_30 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_1_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_1_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_1_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_1_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_1_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_1_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_1_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_1_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_1_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_1_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_1_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_1_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_1_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_1_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_1_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_1_48_port, TO_SHIFT(47) => n241, 
                           TO_SHIFT(46) => A_pos_shifted_by2_1_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_1_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_1_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_1_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_1_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_1_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_1_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_1_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_1_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_1_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_1_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_1_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_1_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_1_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_1_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_1_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_1_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_1_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_1_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_1_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_1_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_1_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_1_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_1_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_1_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_1_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_1_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_1_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_1_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_1_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_1_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_1_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_1_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_1_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_1_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_1_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_1_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_1_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_1_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_1_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_1_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_1_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_1_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_1_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_1_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_1_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_1_0_port, 
                           RESULT(127) => A_pos_shifted_by2_2_63_port, 
                           RESULT(126) => A_pos_shifted_by2_2_62_port, 
                           RESULT(125) => A_pos_shifted_by2_2_61_port, 
                           RESULT(124) => A_pos_shifted_by2_2_60_port, 
                           RESULT(123) => A_pos_shifted_by2_2_59_port, 
                           RESULT(122) => A_pos_shifted_by2_2_58_port, 
                           RESULT(121) => A_pos_shifted_by2_2_57_port, 
                           RESULT(120) => A_pos_shifted_by2_2_56_port, 
                           RESULT(119) => A_pos_shifted_by2_2_55_port, 
                           RESULT(118) => A_pos_shifted_by2_2_54_port, 
                           RESULT(117) => A_pos_shifted_by2_2_53_port, 
                           RESULT(116) => A_pos_shifted_by2_2_52_port, 
                           RESULT(115) => A_pos_shifted_by2_2_51_port, 
                           RESULT(114) => A_pos_shifted_by2_2_50_port, 
                           RESULT(113) => A_pos_shifted_by2_2_49_port, 
                           RESULT(112) => A_pos_shifted_by2_2_48_port, 
                           RESULT(111) => A_pos_shifted_by2_2_47_port, 
                           RESULT(110) => A_pos_shifted_by2_2_46_port, 
                           RESULT(109) => A_pos_shifted_by2_2_45_port, 
                           RESULT(108) => A_pos_shifted_by2_2_44_port, 
                           RESULT(107) => A_pos_shifted_by2_2_43_port, 
                           RESULT(106) => A_pos_shifted_by2_2_42_port, 
                           RESULT(105) => A_pos_shifted_by2_2_41_port, 
                           RESULT(104) => A_pos_shifted_by2_2_40_port, 
                           RESULT(103) => A_pos_shifted_by2_2_39_port, 
                           RESULT(102) => A_pos_shifted_by2_2_38_port, 
                           RESULT(101) => A_pos_shifted_by2_2_37_port, 
                           RESULT(100) => A_pos_shifted_by2_2_36_port, 
                           RESULT(99) => A_pos_shifted_by2_2_35_port, 
                           RESULT(98) => A_pos_shifted_by2_2_34_port, 
                           RESULT(97) => A_pos_shifted_by2_2_33_port, 
                           RESULT(96) => A_pos_shifted_by2_2_32_port, 
                           RESULT(95) => A_pos_shifted_by2_2_31_port, 
                           RESULT(94) => A_pos_shifted_by2_2_30_port, 
                           RESULT(93) => A_pos_shifted_by2_2_29_port, 
                           RESULT(92) => A_pos_shifted_by2_2_28_port, 
                           RESULT(91) => A_pos_shifted_by2_2_27_port, 
                           RESULT(90) => A_pos_shifted_by2_2_26_port, 
                           RESULT(89) => A_pos_shifted_by2_2_25_port, 
                           RESULT(88) => A_pos_shifted_by2_2_24_port, 
                           RESULT(87) => A_pos_shifted_by2_2_23_port, 
                           RESULT(86) => A_pos_shifted_by2_2_22_port, 
                           RESULT(85) => A_pos_shifted_by2_2_21_port, 
                           RESULT(84) => A_pos_shifted_by2_2_20_port, 
                           RESULT(83) => A_pos_shifted_by2_2_19_port, 
                           RESULT(82) => A_pos_shifted_by2_2_18_port, 
                           RESULT(81) => A_pos_shifted_by2_2_17_port, 
                           RESULT(80) => A_pos_shifted_by2_2_16_port, 
                           RESULT(79) => A_pos_shifted_by2_2_15_port, 
                           RESULT(78) => A_pos_shifted_by2_2_14_port, 
                           RESULT(77) => A_pos_shifted_by2_2_13_port, 
                           RESULT(76) => A_pos_shifted_by2_2_12_port, 
                           RESULT(75) => A_pos_shifted_by2_2_11_port, 
                           RESULT(74) => A_pos_shifted_by2_2_10_port, 
                           RESULT(73) => A_pos_shifted_by2_2_9_port, RESULT(72)
                           => A_pos_shifted_by2_2_8_port, RESULT(71) => 
                           A_pos_shifted_by2_2_7_port, RESULT(70) => 
                           A_pos_shifted_by2_2_6_port, RESULT(69) => 
                           A_pos_shifted_by2_2_5_port, RESULT(68) => 
                           A_pos_shifted_by2_2_4_port, RESULT(67) => 
                           A_pos_shifted_by2_2_3_port, RESULT(66) => 
                           A_pos_shifted_by2_2_2_port, RESULT(65) => n_1066, 
                           RESULT(64) => n_1067, RESULT(63) => 
                           A_pos_shifted_by1_2_63_port, RESULT(62) => 
                           A_pos_shifted_by1_2_62_port, RESULT(61) => 
                           A_pos_shifted_by1_2_61_port, RESULT(60) => 
                           A_pos_shifted_by1_2_60_port, RESULT(59) => 
                           A_pos_shifted_by1_2_59_port, RESULT(58) => 
                           A_pos_shifted_by1_2_58_port, RESULT(57) => 
                           A_pos_shifted_by1_2_57_port, RESULT(56) => 
                           A_pos_shifted_by1_2_56_port, RESULT(55) => 
                           A_pos_shifted_by1_2_55_port, RESULT(54) => 
                           A_pos_shifted_by1_2_54_port, RESULT(53) => 
                           A_pos_shifted_by1_2_53_port, RESULT(52) => 
                           A_pos_shifted_by1_2_52_port, RESULT(51) => 
                           A_pos_shifted_by1_2_51_port, RESULT(50) => 
                           A_pos_shifted_by1_2_50_port, RESULT(49) => 
                           A_pos_shifted_by1_2_49_port, RESULT(48) => 
                           A_pos_shifted_by1_2_48_port, RESULT(47) => 
                           A_pos_shifted_by1_2_47_port, RESULT(46) => 
                           A_pos_shifted_by1_2_46_port, RESULT(45) => 
                           A_pos_shifted_by1_2_45_port, RESULT(44) => 
                           A_pos_shifted_by1_2_44_port, RESULT(43) => 
                           A_pos_shifted_by1_2_43_port, RESULT(42) => 
                           A_pos_shifted_by1_2_42_port, RESULT(41) => 
                           A_pos_shifted_by1_2_41_port, RESULT(40) => 
                           A_pos_shifted_by1_2_40_port, RESULT(39) => 
                           A_pos_shifted_by1_2_39_port, RESULT(38) => 
                           A_pos_shifted_by1_2_38_port, RESULT(37) => 
                           A_pos_shifted_by1_2_37_port, RESULT(36) => 
                           A_pos_shifted_by1_2_36_port, RESULT(35) => 
                           A_pos_shifted_by1_2_35_port, RESULT(34) => 
                           A_pos_shifted_by1_2_34_port, RESULT(33) => 
                           A_pos_shifted_by1_2_33_port, RESULT(32) => 
                           A_pos_shifted_by1_2_32_port, RESULT(31) => 
                           A_pos_shifted_by1_2_31_port, RESULT(30) => 
                           A_pos_shifted_by1_2_30_port, RESULT(29) => 
                           A_pos_shifted_by1_2_29_port, RESULT(28) => 
                           A_pos_shifted_by1_2_28_port, RESULT(27) => 
                           A_pos_shifted_by1_2_27_port, RESULT(26) => 
                           A_pos_shifted_by1_2_26_port, RESULT(25) => 
                           A_pos_shifted_by1_2_25_port, RESULT(24) => 
                           A_pos_shifted_by1_2_24_port, RESULT(23) => 
                           A_pos_shifted_by1_2_23_port, RESULT(22) => 
                           A_pos_shifted_by1_2_22_port, RESULT(21) => 
                           A_pos_shifted_by1_2_21_port, RESULT(20) => 
                           A_pos_shifted_by1_2_20_port, RESULT(19) => 
                           A_pos_shifted_by1_2_19_port, RESULT(18) => 
                           A_pos_shifted_by1_2_18_port, RESULT(17) => 
                           A_pos_shifted_by1_2_17_port, RESULT(16) => 
                           A_pos_shifted_by1_2_16_port, RESULT(15) => 
                           A_pos_shifted_by1_2_15_port, RESULT(14) => 
                           A_pos_shifted_by1_2_14_port, RESULT(13) => 
                           A_pos_shifted_by1_2_13_port, RESULT(12) => 
                           A_pos_shifted_by1_2_12_port, RESULT(11) => 
                           A_pos_shifted_by1_2_11_port, RESULT(10) => 
                           A_pos_shifted_by1_2_10_port, RESULT(9) => 
                           A_pos_shifted_by1_2_9_port, RESULT(8) => 
                           A_pos_shifted_by1_2_8_port, RESULT(7) => 
                           A_pos_shifted_by1_2_7_port, RESULT(6) => 
                           A_pos_shifted_by1_2_6_port, RESULT(5) => 
                           A_pos_shifted_by1_2_5_port, RESULT(4) => 
                           A_pos_shifted_by1_2_4_port, RESULT(3) => 
                           A_pos_shifted_by1_2_3_port, RESULT(2) => 
                           A_pos_shifted_by1_2_2_port, RESULT(1) => 
                           A_pos_shifted_by1_2_1_port, RESULT(0) => n_1068);
   SHIFTERi_3 : Shifter_NBIT64_29 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_2_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_2_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_2_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_2_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_2_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_2_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_2_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_2_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_2_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_2_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_2_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_2_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_2_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_2_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_2_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_2_48_port, TO_SHIFT(47) => n240, 
                           TO_SHIFT(46) => A_pos_shifted_by2_2_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_2_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_2_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_2_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_2_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_2_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_2_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_2_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_2_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_2_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_2_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_2_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_2_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_2_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_2_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_2_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_2_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_2_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_2_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_2_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_2_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_2_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_2_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_2_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_2_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_2_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_2_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_2_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_2_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_2_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_2_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_2_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_2_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_2_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_2_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_2_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_2_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_2_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_2_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_2_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_2_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_2_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_2_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_2_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_2_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_2_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_2_0_port, 
                           RESULT(127) => A_pos_shifted_by2_3_63_port, 
                           RESULT(126) => A_pos_shifted_by2_3_62_port, 
                           RESULT(125) => A_pos_shifted_by2_3_61_port, 
                           RESULT(124) => A_pos_shifted_by2_3_60_port, 
                           RESULT(123) => A_pos_shifted_by2_3_59_port, 
                           RESULT(122) => A_pos_shifted_by2_3_58_port, 
                           RESULT(121) => A_pos_shifted_by2_3_57_port, 
                           RESULT(120) => A_pos_shifted_by2_3_56_port, 
                           RESULT(119) => A_pos_shifted_by2_3_55_port, 
                           RESULT(118) => A_pos_shifted_by2_3_54_port, 
                           RESULT(117) => A_pos_shifted_by2_3_53_port, 
                           RESULT(116) => A_pos_shifted_by2_3_52_port, 
                           RESULT(115) => A_pos_shifted_by2_3_51_port, 
                           RESULT(114) => A_pos_shifted_by2_3_50_port, 
                           RESULT(113) => A_pos_shifted_by2_3_49_port, 
                           RESULT(112) => A_pos_shifted_by2_3_48_port, 
                           RESULT(111) => A_pos_shifted_by2_3_47_port, 
                           RESULT(110) => A_pos_shifted_by2_3_46_port, 
                           RESULT(109) => A_pos_shifted_by2_3_45_port, 
                           RESULT(108) => A_pos_shifted_by2_3_44_port, 
                           RESULT(107) => A_pos_shifted_by2_3_43_port, 
                           RESULT(106) => A_pos_shifted_by2_3_42_port, 
                           RESULT(105) => A_pos_shifted_by2_3_41_port, 
                           RESULT(104) => A_pos_shifted_by2_3_40_port, 
                           RESULT(103) => A_pos_shifted_by2_3_39_port, 
                           RESULT(102) => A_pos_shifted_by2_3_38_port, 
                           RESULT(101) => A_pos_shifted_by2_3_37_port, 
                           RESULT(100) => A_pos_shifted_by2_3_36_port, 
                           RESULT(99) => A_pos_shifted_by2_3_35_port, 
                           RESULT(98) => A_pos_shifted_by2_3_34_port, 
                           RESULT(97) => A_pos_shifted_by2_3_33_port, 
                           RESULT(96) => A_pos_shifted_by2_3_32_port, 
                           RESULT(95) => A_pos_shifted_by2_3_31_port, 
                           RESULT(94) => A_pos_shifted_by2_3_30_port, 
                           RESULT(93) => A_pos_shifted_by2_3_29_port, 
                           RESULT(92) => A_pos_shifted_by2_3_28_port, 
                           RESULT(91) => A_pos_shifted_by2_3_27_port, 
                           RESULT(90) => A_pos_shifted_by2_3_26_port, 
                           RESULT(89) => A_pos_shifted_by2_3_25_port, 
                           RESULT(88) => A_pos_shifted_by2_3_24_port, 
                           RESULT(87) => A_pos_shifted_by2_3_23_port, 
                           RESULT(86) => A_pos_shifted_by2_3_22_port, 
                           RESULT(85) => A_pos_shifted_by2_3_21_port, 
                           RESULT(84) => A_pos_shifted_by2_3_20_port, 
                           RESULT(83) => A_pos_shifted_by2_3_19_port, 
                           RESULT(82) => A_pos_shifted_by2_3_18_port, 
                           RESULT(81) => A_pos_shifted_by2_3_17_port, 
                           RESULT(80) => A_pos_shifted_by2_3_16_port, 
                           RESULT(79) => A_pos_shifted_by2_3_15_port, 
                           RESULT(78) => A_pos_shifted_by2_3_14_port, 
                           RESULT(77) => A_pos_shifted_by2_3_13_port, 
                           RESULT(76) => A_pos_shifted_by2_3_12_port, 
                           RESULT(75) => A_pos_shifted_by2_3_11_port, 
                           RESULT(74) => A_pos_shifted_by2_3_10_port, 
                           RESULT(73) => A_pos_shifted_by2_3_9_port, RESULT(72)
                           => A_pos_shifted_by2_3_8_port, RESULT(71) => 
                           A_pos_shifted_by2_3_7_port, RESULT(70) => 
                           A_pos_shifted_by2_3_6_port, RESULT(69) => 
                           A_pos_shifted_by2_3_5_port, RESULT(68) => 
                           A_pos_shifted_by2_3_4_port, RESULT(67) => 
                           A_pos_shifted_by2_3_3_port, RESULT(66) => 
                           A_pos_shifted_by2_3_2_port, RESULT(65) => n_1069, 
                           RESULT(64) => n_1070, RESULT(63) => 
                           A_pos_shifted_by1_3_63_port, RESULT(62) => 
                           A_pos_shifted_by1_3_62_port, RESULT(61) => 
                           A_pos_shifted_by1_3_61_port, RESULT(60) => 
                           A_pos_shifted_by1_3_60_port, RESULT(59) => 
                           A_pos_shifted_by1_3_59_port, RESULT(58) => 
                           A_pos_shifted_by1_3_58_port, RESULT(57) => 
                           A_pos_shifted_by1_3_57_port, RESULT(56) => 
                           A_pos_shifted_by1_3_56_port, RESULT(55) => 
                           A_pos_shifted_by1_3_55_port, RESULT(54) => 
                           A_pos_shifted_by1_3_54_port, RESULT(53) => 
                           A_pos_shifted_by1_3_53_port, RESULT(52) => 
                           A_pos_shifted_by1_3_52_port, RESULT(51) => 
                           A_pos_shifted_by1_3_51_port, RESULT(50) => 
                           A_pos_shifted_by1_3_50_port, RESULT(49) => 
                           A_pos_shifted_by1_3_49_port, RESULT(48) => 
                           A_pos_shifted_by1_3_48_port, RESULT(47) => 
                           A_pos_shifted_by1_3_47_port, RESULT(46) => 
                           A_pos_shifted_by1_3_46_port, RESULT(45) => 
                           A_pos_shifted_by1_3_45_port, RESULT(44) => 
                           A_pos_shifted_by1_3_44_port, RESULT(43) => 
                           A_pos_shifted_by1_3_43_port, RESULT(42) => 
                           A_pos_shifted_by1_3_42_port, RESULT(41) => 
                           A_pos_shifted_by1_3_41_port, RESULT(40) => 
                           A_pos_shifted_by1_3_40_port, RESULT(39) => 
                           A_pos_shifted_by1_3_39_port, RESULT(38) => 
                           A_pos_shifted_by1_3_38_port, RESULT(37) => 
                           A_pos_shifted_by1_3_37_port, RESULT(36) => 
                           A_pos_shifted_by1_3_36_port, RESULT(35) => 
                           A_pos_shifted_by1_3_35_port, RESULT(34) => 
                           A_pos_shifted_by1_3_34_port, RESULT(33) => 
                           A_pos_shifted_by1_3_33_port, RESULT(32) => 
                           A_pos_shifted_by1_3_32_port, RESULT(31) => 
                           A_pos_shifted_by1_3_31_port, RESULT(30) => 
                           A_pos_shifted_by1_3_30_port, RESULT(29) => 
                           A_pos_shifted_by1_3_29_port, RESULT(28) => 
                           A_pos_shifted_by1_3_28_port, RESULT(27) => 
                           A_pos_shifted_by1_3_27_port, RESULT(26) => 
                           A_pos_shifted_by1_3_26_port, RESULT(25) => 
                           A_pos_shifted_by1_3_25_port, RESULT(24) => 
                           A_pos_shifted_by1_3_24_port, RESULT(23) => 
                           A_pos_shifted_by1_3_23_port, RESULT(22) => 
                           A_pos_shifted_by1_3_22_port, RESULT(21) => 
                           A_pos_shifted_by1_3_21_port, RESULT(20) => 
                           A_pos_shifted_by1_3_20_port, RESULT(19) => 
                           A_pos_shifted_by1_3_19_port, RESULT(18) => 
                           A_pos_shifted_by1_3_18_port, RESULT(17) => 
                           A_pos_shifted_by1_3_17_port, RESULT(16) => 
                           A_pos_shifted_by1_3_16_port, RESULT(15) => 
                           A_pos_shifted_by1_3_15_port, RESULT(14) => 
                           A_pos_shifted_by1_3_14_port, RESULT(13) => 
                           A_pos_shifted_by1_3_13_port, RESULT(12) => 
                           A_pos_shifted_by1_3_12_port, RESULT(11) => 
                           A_pos_shifted_by1_3_11_port, RESULT(10) => 
                           A_pos_shifted_by1_3_10_port, RESULT(9) => 
                           A_pos_shifted_by1_3_9_port, RESULT(8) => 
                           A_pos_shifted_by1_3_8_port, RESULT(7) => 
                           A_pos_shifted_by1_3_7_port, RESULT(6) => 
                           A_pos_shifted_by1_3_6_port, RESULT(5) => 
                           A_pos_shifted_by1_3_5_port, RESULT(4) => 
                           A_pos_shifted_by1_3_4_port, RESULT(3) => 
                           A_pos_shifted_by1_3_3_port, RESULT(2) => 
                           A_pos_shifted_by1_3_2_port, RESULT(1) => 
                           A_pos_shifted_by1_3_1_port, RESULT(0) => n_1071);
   SHIFTERi_4 : Shifter_NBIT64_28 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_3_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_3_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_3_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_3_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_3_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_3_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_3_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_3_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_3_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_3_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_3_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_3_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_3_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_3_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_3_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_3_48_port, TO_SHIFT(47) => n239, 
                           TO_SHIFT(46) => A_pos_shifted_by2_3_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_3_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_3_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_3_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_3_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_3_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_3_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_3_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_3_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_3_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_3_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_3_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_3_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_3_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_3_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_3_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_3_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_3_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_3_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_3_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_3_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_3_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_3_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_3_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_3_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_3_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_3_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_3_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_3_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_3_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_3_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_3_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_3_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_3_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_3_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_3_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_3_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_3_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_3_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_3_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_3_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_3_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_3_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_3_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_3_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_3_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_3_0_port, 
                           RESULT(127) => A_pos_shifted_by2_4_63_port, 
                           RESULT(126) => A_pos_shifted_by2_4_62_port, 
                           RESULT(125) => A_pos_shifted_by2_4_61_port, 
                           RESULT(124) => A_pos_shifted_by2_4_60_port, 
                           RESULT(123) => A_pos_shifted_by2_4_59_port, 
                           RESULT(122) => A_pos_shifted_by2_4_58_port, 
                           RESULT(121) => A_pos_shifted_by2_4_57_port, 
                           RESULT(120) => A_pos_shifted_by2_4_56_port, 
                           RESULT(119) => A_pos_shifted_by2_4_55_port, 
                           RESULT(118) => A_pos_shifted_by2_4_54_port, 
                           RESULT(117) => A_pos_shifted_by2_4_53_port, 
                           RESULT(116) => A_pos_shifted_by2_4_52_port, 
                           RESULT(115) => A_pos_shifted_by2_4_51_port, 
                           RESULT(114) => A_pos_shifted_by2_4_50_port, 
                           RESULT(113) => A_pos_shifted_by2_4_49_port, 
                           RESULT(112) => A_pos_shifted_by2_4_48_port, 
                           RESULT(111) => A_pos_shifted_by2_4_47_port, 
                           RESULT(110) => A_pos_shifted_by2_4_46_port, 
                           RESULT(109) => A_pos_shifted_by2_4_45_port, 
                           RESULT(108) => A_pos_shifted_by2_4_44_port, 
                           RESULT(107) => A_pos_shifted_by2_4_43_port, 
                           RESULT(106) => A_pos_shifted_by2_4_42_port, 
                           RESULT(105) => A_pos_shifted_by2_4_41_port, 
                           RESULT(104) => A_pos_shifted_by2_4_40_port, 
                           RESULT(103) => A_pos_shifted_by2_4_39_port, 
                           RESULT(102) => A_pos_shifted_by2_4_38_port, 
                           RESULT(101) => A_pos_shifted_by2_4_37_port, 
                           RESULT(100) => A_pos_shifted_by2_4_36_port, 
                           RESULT(99) => A_pos_shifted_by2_4_35_port, 
                           RESULT(98) => A_pos_shifted_by2_4_34_port, 
                           RESULT(97) => A_pos_shifted_by2_4_33_port, 
                           RESULT(96) => A_pos_shifted_by2_4_32_port, 
                           RESULT(95) => A_pos_shifted_by2_4_31_port, 
                           RESULT(94) => A_pos_shifted_by2_4_30_port, 
                           RESULT(93) => A_pos_shifted_by2_4_29_port, 
                           RESULT(92) => A_pos_shifted_by2_4_28_port, 
                           RESULT(91) => A_pos_shifted_by2_4_27_port, 
                           RESULT(90) => A_pos_shifted_by2_4_26_port, 
                           RESULT(89) => A_pos_shifted_by2_4_25_port, 
                           RESULT(88) => A_pos_shifted_by2_4_24_port, 
                           RESULT(87) => A_pos_shifted_by2_4_23_port, 
                           RESULT(86) => A_pos_shifted_by2_4_22_port, 
                           RESULT(85) => A_pos_shifted_by2_4_21_port, 
                           RESULT(84) => A_pos_shifted_by2_4_20_port, 
                           RESULT(83) => A_pos_shifted_by2_4_19_port, 
                           RESULT(82) => A_pos_shifted_by2_4_18_port, 
                           RESULT(81) => A_pos_shifted_by2_4_17_port, 
                           RESULT(80) => A_pos_shifted_by2_4_16_port, 
                           RESULT(79) => A_pos_shifted_by2_4_15_port, 
                           RESULT(78) => A_pos_shifted_by2_4_14_port, 
                           RESULT(77) => A_pos_shifted_by2_4_13_port, 
                           RESULT(76) => A_pos_shifted_by2_4_12_port, 
                           RESULT(75) => A_pos_shifted_by2_4_11_port, 
                           RESULT(74) => A_pos_shifted_by2_4_10_port, 
                           RESULT(73) => A_pos_shifted_by2_4_9_port, RESULT(72)
                           => A_pos_shifted_by2_4_8_port, RESULT(71) => 
                           A_pos_shifted_by2_4_7_port, RESULT(70) => 
                           A_pos_shifted_by2_4_6_port, RESULT(69) => 
                           A_pos_shifted_by2_4_5_port, RESULT(68) => 
                           A_pos_shifted_by2_4_4_port, RESULT(67) => 
                           A_pos_shifted_by2_4_3_port, RESULT(66) => 
                           A_pos_shifted_by2_4_2_port, RESULT(65) => n_1072, 
                           RESULT(64) => n_1073, RESULT(63) => 
                           A_pos_shifted_by1_4_63_port, RESULT(62) => 
                           A_pos_shifted_by1_4_62_port, RESULT(61) => 
                           A_pos_shifted_by1_4_61_port, RESULT(60) => 
                           A_pos_shifted_by1_4_60_port, RESULT(59) => 
                           A_pos_shifted_by1_4_59_port, RESULT(58) => 
                           A_pos_shifted_by1_4_58_port, RESULT(57) => 
                           A_pos_shifted_by1_4_57_port, RESULT(56) => 
                           A_pos_shifted_by1_4_56_port, RESULT(55) => 
                           A_pos_shifted_by1_4_55_port, RESULT(54) => 
                           A_pos_shifted_by1_4_54_port, RESULT(53) => 
                           A_pos_shifted_by1_4_53_port, RESULT(52) => 
                           A_pos_shifted_by1_4_52_port, RESULT(51) => 
                           A_pos_shifted_by1_4_51_port, RESULT(50) => 
                           A_pos_shifted_by1_4_50_port, RESULT(49) => 
                           A_pos_shifted_by1_4_49_port, RESULT(48) => 
                           A_pos_shifted_by1_4_48_port, RESULT(47) => 
                           A_pos_shifted_by1_4_47_port, RESULT(46) => 
                           A_pos_shifted_by1_4_46_port, RESULT(45) => 
                           A_pos_shifted_by1_4_45_port, RESULT(44) => 
                           A_pos_shifted_by1_4_44_port, RESULT(43) => 
                           A_pos_shifted_by1_4_43_port, RESULT(42) => 
                           A_pos_shifted_by1_4_42_port, RESULT(41) => 
                           A_pos_shifted_by1_4_41_port, RESULT(40) => 
                           A_pos_shifted_by1_4_40_port, RESULT(39) => 
                           A_pos_shifted_by1_4_39_port, RESULT(38) => 
                           A_pos_shifted_by1_4_38_port, RESULT(37) => 
                           A_pos_shifted_by1_4_37_port, RESULT(36) => 
                           A_pos_shifted_by1_4_36_port, RESULT(35) => 
                           A_pos_shifted_by1_4_35_port, RESULT(34) => 
                           A_pos_shifted_by1_4_34_port, RESULT(33) => 
                           A_pos_shifted_by1_4_33_port, RESULT(32) => 
                           A_pos_shifted_by1_4_32_port, RESULT(31) => 
                           A_pos_shifted_by1_4_31_port, RESULT(30) => 
                           A_pos_shifted_by1_4_30_port, RESULT(29) => 
                           A_pos_shifted_by1_4_29_port, RESULT(28) => 
                           A_pos_shifted_by1_4_28_port, RESULT(27) => 
                           A_pos_shifted_by1_4_27_port, RESULT(26) => 
                           A_pos_shifted_by1_4_26_port, RESULT(25) => 
                           A_pos_shifted_by1_4_25_port, RESULT(24) => 
                           A_pos_shifted_by1_4_24_port, RESULT(23) => 
                           A_pos_shifted_by1_4_23_port, RESULT(22) => 
                           A_pos_shifted_by1_4_22_port, RESULT(21) => 
                           A_pos_shifted_by1_4_21_port, RESULT(20) => 
                           A_pos_shifted_by1_4_20_port, RESULT(19) => 
                           A_pos_shifted_by1_4_19_port, RESULT(18) => 
                           A_pos_shifted_by1_4_18_port, RESULT(17) => 
                           A_pos_shifted_by1_4_17_port, RESULT(16) => 
                           A_pos_shifted_by1_4_16_port, RESULT(15) => 
                           A_pos_shifted_by1_4_15_port, RESULT(14) => 
                           A_pos_shifted_by1_4_14_port, RESULT(13) => 
                           A_pos_shifted_by1_4_13_port, RESULT(12) => 
                           A_pos_shifted_by1_4_12_port, RESULT(11) => 
                           A_pos_shifted_by1_4_11_port, RESULT(10) => 
                           A_pos_shifted_by1_4_10_port, RESULT(9) => 
                           A_pos_shifted_by1_4_9_port, RESULT(8) => 
                           A_pos_shifted_by1_4_8_port, RESULT(7) => 
                           A_pos_shifted_by1_4_7_port, RESULT(6) => 
                           A_pos_shifted_by1_4_6_port, RESULT(5) => 
                           A_pos_shifted_by1_4_5_port, RESULT(4) => 
                           A_pos_shifted_by1_4_4_port, RESULT(3) => 
                           A_pos_shifted_by1_4_3_port, RESULT(2) => 
                           A_pos_shifted_by1_4_2_port, RESULT(1) => 
                           A_pos_shifted_by1_4_1_port, RESULT(0) => n_1074);
   SHIFTERi_5 : Shifter_NBIT64_27 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_4_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_4_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_4_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_4_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_4_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_4_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_4_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_4_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_4_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_4_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_4_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_4_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_4_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_4_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_4_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_4_48_port, TO_SHIFT(47) => n238, 
                           TO_SHIFT(46) => A_pos_shifted_by2_4_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_4_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_4_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_4_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_4_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_4_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_4_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_4_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_4_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_4_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_4_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_4_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_4_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_4_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_4_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_4_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_4_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_4_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_4_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_4_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_4_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_4_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_4_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_4_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_4_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_4_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_4_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_4_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_4_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_4_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_4_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_4_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_4_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_4_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_4_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_4_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_4_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_4_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_4_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_4_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_4_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_4_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_4_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_4_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_4_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_4_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_4_0_port, 
                           RESULT(127) => A_pos_shifted_by2_5_63_port, 
                           RESULT(126) => A_pos_shifted_by2_5_62_port, 
                           RESULT(125) => A_pos_shifted_by2_5_61_port, 
                           RESULT(124) => A_pos_shifted_by2_5_60_port, 
                           RESULT(123) => A_pos_shifted_by2_5_59_port, 
                           RESULT(122) => A_pos_shifted_by2_5_58_port, 
                           RESULT(121) => A_pos_shifted_by2_5_57_port, 
                           RESULT(120) => A_pos_shifted_by2_5_56_port, 
                           RESULT(119) => A_pos_shifted_by2_5_55_port, 
                           RESULT(118) => A_pos_shifted_by2_5_54_port, 
                           RESULT(117) => A_pos_shifted_by2_5_53_port, 
                           RESULT(116) => A_pos_shifted_by2_5_52_port, 
                           RESULT(115) => A_pos_shifted_by2_5_51_port, 
                           RESULT(114) => A_pos_shifted_by2_5_50_port, 
                           RESULT(113) => A_pos_shifted_by2_5_49_port, 
                           RESULT(112) => A_pos_shifted_by2_5_48_port, 
                           RESULT(111) => A_pos_shifted_by2_5_47_port, 
                           RESULT(110) => A_pos_shifted_by2_5_46_port, 
                           RESULT(109) => A_pos_shifted_by2_5_45_port, 
                           RESULT(108) => A_pos_shifted_by2_5_44_port, 
                           RESULT(107) => A_pos_shifted_by2_5_43_port, 
                           RESULT(106) => A_pos_shifted_by2_5_42_port, 
                           RESULT(105) => A_pos_shifted_by2_5_41_port, 
                           RESULT(104) => A_pos_shifted_by2_5_40_port, 
                           RESULT(103) => A_pos_shifted_by2_5_39_port, 
                           RESULT(102) => A_pos_shifted_by2_5_38_port, 
                           RESULT(101) => A_pos_shifted_by2_5_37_port, 
                           RESULT(100) => A_pos_shifted_by2_5_36_port, 
                           RESULT(99) => A_pos_shifted_by2_5_35_port, 
                           RESULT(98) => A_pos_shifted_by2_5_34_port, 
                           RESULT(97) => A_pos_shifted_by2_5_33_port, 
                           RESULT(96) => A_pos_shifted_by2_5_32_port, 
                           RESULT(95) => A_pos_shifted_by2_5_31_port, 
                           RESULT(94) => A_pos_shifted_by2_5_30_port, 
                           RESULT(93) => A_pos_shifted_by2_5_29_port, 
                           RESULT(92) => A_pos_shifted_by2_5_28_port, 
                           RESULT(91) => A_pos_shifted_by2_5_27_port, 
                           RESULT(90) => A_pos_shifted_by2_5_26_port, 
                           RESULT(89) => A_pos_shifted_by2_5_25_port, 
                           RESULT(88) => A_pos_shifted_by2_5_24_port, 
                           RESULT(87) => A_pos_shifted_by2_5_23_port, 
                           RESULT(86) => A_pos_shifted_by2_5_22_port, 
                           RESULT(85) => A_pos_shifted_by2_5_21_port, 
                           RESULT(84) => A_pos_shifted_by2_5_20_port, 
                           RESULT(83) => A_pos_shifted_by2_5_19_port, 
                           RESULT(82) => A_pos_shifted_by2_5_18_port, 
                           RESULT(81) => A_pos_shifted_by2_5_17_port, 
                           RESULT(80) => A_pos_shifted_by2_5_16_port, 
                           RESULT(79) => A_pos_shifted_by2_5_15_port, 
                           RESULT(78) => A_pos_shifted_by2_5_14_port, 
                           RESULT(77) => A_pos_shifted_by2_5_13_port, 
                           RESULT(76) => A_pos_shifted_by2_5_12_port, 
                           RESULT(75) => A_pos_shifted_by2_5_11_port, 
                           RESULT(74) => A_pos_shifted_by2_5_10_port, 
                           RESULT(73) => A_pos_shifted_by2_5_9_port, RESULT(72)
                           => A_pos_shifted_by2_5_8_port, RESULT(71) => 
                           A_pos_shifted_by2_5_7_port, RESULT(70) => 
                           A_pos_shifted_by2_5_6_port, RESULT(69) => 
                           A_pos_shifted_by2_5_5_port, RESULT(68) => 
                           A_pos_shifted_by2_5_4_port, RESULT(67) => 
                           A_pos_shifted_by2_5_3_port, RESULT(66) => 
                           A_pos_shifted_by2_5_2_port, RESULT(65) => n_1075, 
                           RESULT(64) => n_1076, RESULT(63) => 
                           A_pos_shifted_by1_5_63_port, RESULT(62) => 
                           A_pos_shifted_by1_5_62_port, RESULT(61) => 
                           A_pos_shifted_by1_5_61_port, RESULT(60) => 
                           A_pos_shifted_by1_5_60_port, RESULT(59) => 
                           A_pos_shifted_by1_5_59_port, RESULT(58) => 
                           A_pos_shifted_by1_5_58_port, RESULT(57) => 
                           A_pos_shifted_by1_5_57_port, RESULT(56) => 
                           A_pos_shifted_by1_5_56_port, RESULT(55) => 
                           A_pos_shifted_by1_5_55_port, RESULT(54) => 
                           A_pos_shifted_by1_5_54_port, RESULT(53) => 
                           A_pos_shifted_by1_5_53_port, RESULT(52) => 
                           A_pos_shifted_by1_5_52_port, RESULT(51) => 
                           A_pos_shifted_by1_5_51_port, RESULT(50) => 
                           A_pos_shifted_by1_5_50_port, RESULT(49) => 
                           A_pos_shifted_by1_5_49_port, RESULT(48) => 
                           A_pos_shifted_by1_5_48_port, RESULT(47) => 
                           A_pos_shifted_by1_5_47_port, RESULT(46) => 
                           A_pos_shifted_by1_5_46_port, RESULT(45) => 
                           A_pos_shifted_by1_5_45_port, RESULT(44) => 
                           A_pos_shifted_by1_5_44_port, RESULT(43) => 
                           A_pos_shifted_by1_5_43_port, RESULT(42) => 
                           A_pos_shifted_by1_5_42_port, RESULT(41) => 
                           A_pos_shifted_by1_5_41_port, RESULT(40) => 
                           A_pos_shifted_by1_5_40_port, RESULT(39) => 
                           A_pos_shifted_by1_5_39_port, RESULT(38) => 
                           A_pos_shifted_by1_5_38_port, RESULT(37) => 
                           A_pos_shifted_by1_5_37_port, RESULT(36) => 
                           A_pos_shifted_by1_5_36_port, RESULT(35) => 
                           A_pos_shifted_by1_5_35_port, RESULT(34) => 
                           A_pos_shifted_by1_5_34_port, RESULT(33) => 
                           A_pos_shifted_by1_5_33_port, RESULT(32) => 
                           A_pos_shifted_by1_5_32_port, RESULT(31) => 
                           A_pos_shifted_by1_5_31_port, RESULT(30) => 
                           A_pos_shifted_by1_5_30_port, RESULT(29) => 
                           A_pos_shifted_by1_5_29_port, RESULT(28) => 
                           A_pos_shifted_by1_5_28_port, RESULT(27) => 
                           A_pos_shifted_by1_5_27_port, RESULT(26) => 
                           A_pos_shifted_by1_5_26_port, RESULT(25) => 
                           A_pos_shifted_by1_5_25_port, RESULT(24) => 
                           A_pos_shifted_by1_5_24_port, RESULT(23) => 
                           A_pos_shifted_by1_5_23_port, RESULT(22) => 
                           A_pos_shifted_by1_5_22_port, RESULT(21) => 
                           A_pos_shifted_by1_5_21_port, RESULT(20) => 
                           A_pos_shifted_by1_5_20_port, RESULT(19) => 
                           A_pos_shifted_by1_5_19_port, RESULT(18) => 
                           A_pos_shifted_by1_5_18_port, RESULT(17) => 
                           A_pos_shifted_by1_5_17_port, RESULT(16) => 
                           A_pos_shifted_by1_5_16_port, RESULT(15) => 
                           A_pos_shifted_by1_5_15_port, RESULT(14) => 
                           A_pos_shifted_by1_5_14_port, RESULT(13) => 
                           A_pos_shifted_by1_5_13_port, RESULT(12) => 
                           A_pos_shifted_by1_5_12_port, RESULT(11) => 
                           A_pos_shifted_by1_5_11_port, RESULT(10) => 
                           A_pos_shifted_by1_5_10_port, RESULT(9) => 
                           A_pos_shifted_by1_5_9_port, RESULT(8) => 
                           A_pos_shifted_by1_5_8_port, RESULT(7) => 
                           A_pos_shifted_by1_5_7_port, RESULT(6) => 
                           A_pos_shifted_by1_5_6_port, RESULT(5) => 
                           A_pos_shifted_by1_5_5_port, RESULT(4) => 
                           A_pos_shifted_by1_5_4_port, RESULT(3) => 
                           A_pos_shifted_by1_5_3_port, RESULT(2) => 
                           A_pos_shifted_by1_5_2_port, RESULT(1) => 
                           A_pos_shifted_by1_5_1_port, RESULT(0) => n_1077);
   SHIFTERi_6 : Shifter_NBIT64_26 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_5_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_5_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_5_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_5_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_5_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_5_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_5_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_5_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_5_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_5_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_5_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_5_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_5_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_5_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_5_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_5_48_port, TO_SHIFT(47) => n237, 
                           TO_SHIFT(46) => A_pos_shifted_by2_5_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_5_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_5_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_5_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_5_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_5_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_5_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_5_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_5_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_5_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_5_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_5_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_5_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_5_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_5_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_5_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_5_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_5_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_5_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_5_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_5_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_5_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_5_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_5_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_5_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_5_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_5_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_5_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_5_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_5_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_5_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_5_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_5_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_5_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_5_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_5_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_5_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_5_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_5_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_5_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_5_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_5_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_5_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_5_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_5_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_5_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_5_0_port, 
                           RESULT(127) => A_pos_shifted_by2_6_63_port, 
                           RESULT(126) => A_pos_shifted_by2_6_62_port, 
                           RESULT(125) => A_pos_shifted_by2_6_61_port, 
                           RESULT(124) => A_pos_shifted_by2_6_60_port, 
                           RESULT(123) => A_pos_shifted_by2_6_59_port, 
                           RESULT(122) => A_pos_shifted_by2_6_58_port, 
                           RESULT(121) => A_pos_shifted_by2_6_57_port, 
                           RESULT(120) => A_pos_shifted_by2_6_56_port, 
                           RESULT(119) => A_pos_shifted_by2_6_55_port, 
                           RESULT(118) => A_pos_shifted_by2_6_54_port, 
                           RESULT(117) => A_pos_shifted_by2_6_53_port, 
                           RESULT(116) => A_pos_shifted_by2_6_52_port, 
                           RESULT(115) => A_pos_shifted_by2_6_51_port, 
                           RESULT(114) => A_pos_shifted_by2_6_50_port, 
                           RESULT(113) => A_pos_shifted_by2_6_49_port, 
                           RESULT(112) => A_pos_shifted_by2_6_48_port, 
                           RESULT(111) => A_pos_shifted_by2_6_47_port, 
                           RESULT(110) => A_pos_shifted_by2_6_46_port, 
                           RESULT(109) => A_pos_shifted_by2_6_45_port, 
                           RESULT(108) => A_pos_shifted_by2_6_44_port, 
                           RESULT(107) => A_pos_shifted_by2_6_43_port, 
                           RESULT(106) => A_pos_shifted_by2_6_42_port, 
                           RESULT(105) => A_pos_shifted_by2_6_41_port, 
                           RESULT(104) => A_pos_shifted_by2_6_40_port, 
                           RESULT(103) => A_pos_shifted_by2_6_39_port, 
                           RESULT(102) => A_pos_shifted_by2_6_38_port, 
                           RESULT(101) => A_pos_shifted_by2_6_37_port, 
                           RESULT(100) => A_pos_shifted_by2_6_36_port, 
                           RESULT(99) => A_pos_shifted_by2_6_35_port, 
                           RESULT(98) => A_pos_shifted_by2_6_34_port, 
                           RESULT(97) => A_pos_shifted_by2_6_33_port, 
                           RESULT(96) => A_pos_shifted_by2_6_32_port, 
                           RESULT(95) => A_pos_shifted_by2_6_31_port, 
                           RESULT(94) => A_pos_shifted_by2_6_30_port, 
                           RESULT(93) => A_pos_shifted_by2_6_29_port, 
                           RESULT(92) => A_pos_shifted_by2_6_28_port, 
                           RESULT(91) => A_pos_shifted_by2_6_27_port, 
                           RESULT(90) => A_pos_shifted_by2_6_26_port, 
                           RESULT(89) => A_pos_shifted_by2_6_25_port, 
                           RESULT(88) => A_pos_shifted_by2_6_24_port, 
                           RESULT(87) => A_pos_shifted_by2_6_23_port, 
                           RESULT(86) => A_pos_shifted_by2_6_22_port, 
                           RESULT(85) => A_pos_shifted_by2_6_21_port, 
                           RESULT(84) => A_pos_shifted_by2_6_20_port, 
                           RESULT(83) => A_pos_shifted_by2_6_19_port, 
                           RESULT(82) => A_pos_shifted_by2_6_18_port, 
                           RESULT(81) => A_pos_shifted_by2_6_17_port, 
                           RESULT(80) => A_pos_shifted_by2_6_16_port, 
                           RESULT(79) => A_pos_shifted_by2_6_15_port, 
                           RESULT(78) => A_pos_shifted_by2_6_14_port, 
                           RESULT(77) => A_pos_shifted_by2_6_13_port, 
                           RESULT(76) => A_pos_shifted_by2_6_12_port, 
                           RESULT(75) => A_pos_shifted_by2_6_11_port, 
                           RESULT(74) => A_pos_shifted_by2_6_10_port, 
                           RESULT(73) => A_pos_shifted_by2_6_9_port, RESULT(72)
                           => A_pos_shifted_by2_6_8_port, RESULT(71) => 
                           A_pos_shifted_by2_6_7_port, RESULT(70) => 
                           A_pos_shifted_by2_6_6_port, RESULT(69) => 
                           A_pos_shifted_by2_6_5_port, RESULT(68) => 
                           A_pos_shifted_by2_6_4_port, RESULT(67) => 
                           A_pos_shifted_by2_6_3_port, RESULT(66) => 
                           A_pos_shifted_by2_6_2_port, RESULT(65) => n_1078, 
                           RESULT(64) => n_1079, RESULT(63) => 
                           A_pos_shifted_by1_6_63_port, RESULT(62) => 
                           A_pos_shifted_by1_6_62_port, RESULT(61) => 
                           A_pos_shifted_by1_6_61_port, RESULT(60) => 
                           A_pos_shifted_by1_6_60_port, RESULT(59) => 
                           A_pos_shifted_by1_6_59_port, RESULT(58) => 
                           A_pos_shifted_by1_6_58_port, RESULT(57) => 
                           A_pos_shifted_by1_6_57_port, RESULT(56) => 
                           A_pos_shifted_by1_6_56_port, RESULT(55) => 
                           A_pos_shifted_by1_6_55_port, RESULT(54) => 
                           A_pos_shifted_by1_6_54_port, RESULT(53) => 
                           A_pos_shifted_by1_6_53_port, RESULT(52) => 
                           A_pos_shifted_by1_6_52_port, RESULT(51) => 
                           A_pos_shifted_by1_6_51_port, RESULT(50) => 
                           A_pos_shifted_by1_6_50_port, RESULT(49) => 
                           A_pos_shifted_by1_6_49_port, RESULT(48) => 
                           A_pos_shifted_by1_6_48_port, RESULT(47) => 
                           A_pos_shifted_by1_6_47_port, RESULT(46) => 
                           A_pos_shifted_by1_6_46_port, RESULT(45) => 
                           A_pos_shifted_by1_6_45_port, RESULT(44) => 
                           A_pos_shifted_by1_6_44_port, RESULT(43) => 
                           A_pos_shifted_by1_6_43_port, RESULT(42) => 
                           A_pos_shifted_by1_6_42_port, RESULT(41) => 
                           A_pos_shifted_by1_6_41_port, RESULT(40) => 
                           A_pos_shifted_by1_6_40_port, RESULT(39) => 
                           A_pos_shifted_by1_6_39_port, RESULT(38) => 
                           A_pos_shifted_by1_6_38_port, RESULT(37) => 
                           A_pos_shifted_by1_6_37_port, RESULT(36) => 
                           A_pos_shifted_by1_6_36_port, RESULT(35) => 
                           A_pos_shifted_by1_6_35_port, RESULT(34) => 
                           A_pos_shifted_by1_6_34_port, RESULT(33) => 
                           A_pos_shifted_by1_6_33_port, RESULT(32) => 
                           A_pos_shifted_by1_6_32_port, RESULT(31) => 
                           A_pos_shifted_by1_6_31_port, RESULT(30) => 
                           A_pos_shifted_by1_6_30_port, RESULT(29) => 
                           A_pos_shifted_by1_6_29_port, RESULT(28) => 
                           A_pos_shifted_by1_6_28_port, RESULT(27) => 
                           A_pos_shifted_by1_6_27_port, RESULT(26) => 
                           A_pos_shifted_by1_6_26_port, RESULT(25) => 
                           A_pos_shifted_by1_6_25_port, RESULT(24) => 
                           A_pos_shifted_by1_6_24_port, RESULT(23) => 
                           A_pos_shifted_by1_6_23_port, RESULT(22) => 
                           A_pos_shifted_by1_6_22_port, RESULT(21) => 
                           A_pos_shifted_by1_6_21_port, RESULT(20) => 
                           A_pos_shifted_by1_6_20_port, RESULT(19) => 
                           A_pos_shifted_by1_6_19_port, RESULT(18) => 
                           A_pos_shifted_by1_6_18_port, RESULT(17) => 
                           A_pos_shifted_by1_6_17_port, RESULT(16) => 
                           A_pos_shifted_by1_6_16_port, RESULT(15) => 
                           A_pos_shifted_by1_6_15_port, RESULT(14) => 
                           A_pos_shifted_by1_6_14_port, RESULT(13) => 
                           A_pos_shifted_by1_6_13_port, RESULT(12) => 
                           A_pos_shifted_by1_6_12_port, RESULT(11) => 
                           A_pos_shifted_by1_6_11_port, RESULT(10) => 
                           A_pos_shifted_by1_6_10_port, RESULT(9) => 
                           A_pos_shifted_by1_6_9_port, RESULT(8) => 
                           A_pos_shifted_by1_6_8_port, RESULT(7) => 
                           A_pos_shifted_by1_6_7_port, RESULT(6) => 
                           A_pos_shifted_by1_6_6_port, RESULT(5) => 
                           A_pos_shifted_by1_6_5_port, RESULT(4) => 
                           A_pos_shifted_by1_6_4_port, RESULT(3) => 
                           A_pos_shifted_by1_6_3_port, RESULT(2) => 
                           A_pos_shifted_by1_6_2_port, RESULT(1) => 
                           A_pos_shifted_by1_6_1_port, RESULT(0) => n_1080);
   SHIFTERi_7 : Shifter_NBIT64_25 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_6_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_6_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_6_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_6_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_6_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_6_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_6_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_6_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_6_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_6_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_6_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_6_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_6_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_6_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_6_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_6_48_port, TO_SHIFT(47) => n236, 
                           TO_SHIFT(46) => A_pos_shifted_by2_6_46_port, 
                           TO_SHIFT(45) => A_pos_shifted_by2_6_45_port, 
                           TO_SHIFT(44) => A_pos_shifted_by2_6_44_port, 
                           TO_SHIFT(43) => A_pos_shifted_by2_6_43_port, 
                           TO_SHIFT(42) => A_pos_shifted_by2_6_42_port, 
                           TO_SHIFT(41) => A_pos_shifted_by2_6_41_port, 
                           TO_SHIFT(40) => A_pos_shifted_by2_6_40_port, 
                           TO_SHIFT(39) => A_pos_shifted_by2_6_39_port, 
                           TO_SHIFT(38) => A_pos_shifted_by2_6_38_port, 
                           TO_SHIFT(37) => A_pos_shifted_by2_6_37_port, 
                           TO_SHIFT(36) => A_pos_shifted_by2_6_36_port, 
                           TO_SHIFT(35) => A_pos_shifted_by2_6_35_port, 
                           TO_SHIFT(34) => A_pos_shifted_by2_6_34_port, 
                           TO_SHIFT(33) => A_pos_shifted_by2_6_33_port, 
                           TO_SHIFT(32) => A_pos_shifted_by2_6_32_port, 
                           TO_SHIFT(31) => A_pos_shifted_by2_6_31_port, 
                           TO_SHIFT(30) => A_pos_shifted_by2_6_30_port, 
                           TO_SHIFT(29) => A_pos_shifted_by2_6_29_port, 
                           TO_SHIFT(28) => A_pos_shifted_by2_6_28_port, 
                           TO_SHIFT(27) => A_pos_shifted_by2_6_27_port, 
                           TO_SHIFT(26) => A_pos_shifted_by2_6_26_port, 
                           TO_SHIFT(25) => A_pos_shifted_by2_6_25_port, 
                           TO_SHIFT(24) => A_pos_shifted_by2_6_24_port, 
                           TO_SHIFT(23) => A_pos_shifted_by2_6_23_port, 
                           TO_SHIFT(22) => A_pos_shifted_by2_6_22_port, 
                           TO_SHIFT(21) => A_pos_shifted_by2_6_21_port, 
                           TO_SHIFT(20) => A_pos_shifted_by2_6_20_port, 
                           TO_SHIFT(19) => A_pos_shifted_by2_6_19_port, 
                           TO_SHIFT(18) => A_pos_shifted_by2_6_18_port, 
                           TO_SHIFT(17) => A_pos_shifted_by2_6_17_port, 
                           TO_SHIFT(16) => A_pos_shifted_by2_6_16_port, 
                           TO_SHIFT(15) => A_pos_shifted_by2_6_15_port, 
                           TO_SHIFT(14) => A_pos_shifted_by2_6_14_port, 
                           TO_SHIFT(13) => A_pos_shifted_by2_6_13_port, 
                           TO_SHIFT(12) => A_pos_shifted_by2_6_12_port, 
                           TO_SHIFT(11) => A_pos_shifted_by2_6_11_port, 
                           TO_SHIFT(10) => A_pos_shifted_by2_6_10_port, 
                           TO_SHIFT(9) => A_pos_shifted_by2_6_9_port, 
                           TO_SHIFT(8) => A_pos_shifted_by2_6_8_port, 
                           TO_SHIFT(7) => A_pos_shifted_by2_6_7_port, 
                           TO_SHIFT(6) => A_pos_shifted_by2_6_6_port, 
                           TO_SHIFT(5) => A_pos_shifted_by2_6_5_port, 
                           TO_SHIFT(4) => A_pos_shifted_by2_6_4_port, 
                           TO_SHIFT(3) => A_pos_shifted_by2_6_3_port, 
                           TO_SHIFT(2) => A_pos_shifted_by2_6_2_port, 
                           TO_SHIFT(1) => A_pos_shifted_by2_6_1_port, 
                           TO_SHIFT(0) => A_pos_shifted_by2_6_0_port, 
                           RESULT(127) => A_pos_shifted_by2_7_63_port, 
                           RESULT(126) => A_pos_shifted_by2_7_62_port, 
                           RESULT(125) => A_pos_shifted_by2_7_61_port, 
                           RESULT(124) => A_pos_shifted_by2_7_60_port, 
                           RESULT(123) => A_pos_shifted_by2_7_59_port, 
                           RESULT(122) => A_pos_shifted_by2_7_58_port, 
                           RESULT(121) => A_pos_shifted_by2_7_57_port, 
                           RESULT(120) => A_pos_shifted_by2_7_56_port, 
                           RESULT(119) => A_pos_shifted_by2_7_55_port, 
                           RESULT(118) => A_pos_shifted_by2_7_54_port, 
                           RESULT(117) => A_pos_shifted_by2_7_53_port, 
                           RESULT(116) => A_pos_shifted_by2_7_52_port, 
                           RESULT(115) => A_pos_shifted_by2_7_51_port, 
                           RESULT(114) => A_pos_shifted_by2_7_50_port, 
                           RESULT(113) => A_pos_shifted_by2_7_49_port, 
                           RESULT(112) => A_pos_shifted_by2_7_48_port, 
                           RESULT(111) => A_pos_shifted_by2_7_47_port, 
                           RESULT(110) => A_pos_shifted_by2_7_46_port, 
                           RESULT(109) => A_pos_shifted_by2_7_45_port, 
                           RESULT(108) => A_pos_shifted_by2_7_44_port, 
                           RESULT(107) => A_pos_shifted_by2_7_43_port, 
                           RESULT(106) => A_pos_shifted_by2_7_42_port, 
                           RESULT(105) => A_pos_shifted_by2_7_41_port, 
                           RESULT(104) => A_pos_shifted_by2_7_40_port, 
                           RESULT(103) => A_pos_shifted_by2_7_39_port, 
                           RESULT(102) => A_pos_shifted_by2_7_38_port, 
                           RESULT(101) => A_pos_shifted_by2_7_37_port, 
                           RESULT(100) => A_pos_shifted_by2_7_36_port, 
                           RESULT(99) => A_pos_shifted_by2_7_35_port, 
                           RESULT(98) => A_pos_shifted_by2_7_34_port, 
                           RESULT(97) => A_pos_shifted_by2_7_33_port, 
                           RESULT(96) => A_pos_shifted_by2_7_32_port, 
                           RESULT(95) => A_pos_shifted_by2_7_31_port, 
                           RESULT(94) => A_pos_shifted_by2_7_30_port, 
                           RESULT(93) => A_pos_shifted_by2_7_29_port, 
                           RESULT(92) => A_pos_shifted_by2_7_28_port, 
                           RESULT(91) => A_pos_shifted_by2_7_27_port, 
                           RESULT(90) => A_pos_shifted_by2_7_26_port, 
                           RESULT(89) => A_pos_shifted_by2_7_25_port, 
                           RESULT(88) => A_pos_shifted_by2_7_24_port, 
                           RESULT(87) => A_pos_shifted_by2_7_23_port, 
                           RESULT(86) => A_pos_shifted_by2_7_22_port, 
                           RESULT(85) => A_pos_shifted_by2_7_21_port, 
                           RESULT(84) => A_pos_shifted_by2_7_20_port, 
                           RESULT(83) => A_pos_shifted_by2_7_19_port, 
                           RESULT(82) => A_pos_shifted_by2_7_18_port, 
                           RESULT(81) => A_pos_shifted_by2_7_17_port, 
                           RESULT(80) => A_pos_shifted_by2_7_16_port, 
                           RESULT(79) => A_pos_shifted_by2_7_15_port, 
                           RESULT(78) => A_pos_shifted_by2_7_14_port, 
                           RESULT(77) => A_pos_shifted_by2_7_13_port, 
                           RESULT(76) => A_pos_shifted_by2_7_12_port, 
                           RESULT(75) => A_pos_shifted_by2_7_11_port, 
                           RESULT(74) => A_pos_shifted_by2_7_10_port, 
                           RESULT(73) => A_pos_shifted_by2_7_9_port, RESULT(72)
                           => A_pos_shifted_by2_7_8_port, RESULT(71) => 
                           A_pos_shifted_by2_7_7_port, RESULT(70) => 
                           A_pos_shifted_by2_7_6_port, RESULT(69) => 
                           A_pos_shifted_by2_7_5_port, RESULT(68) => 
                           A_pos_shifted_by2_7_4_port, RESULT(67) => 
                           A_pos_shifted_by2_7_3_port, RESULT(66) => 
                           A_pos_shifted_by2_7_2_port, RESULT(65) => n_1081, 
                           RESULT(64) => n_1082, RESULT(63) => 
                           A_pos_shifted_by1_7_63_port, RESULT(62) => 
                           A_pos_shifted_by1_7_62_port, RESULT(61) => 
                           A_pos_shifted_by1_7_61_port, RESULT(60) => 
                           A_pos_shifted_by1_7_60_port, RESULT(59) => 
                           A_pos_shifted_by1_7_59_port, RESULT(58) => 
                           A_pos_shifted_by1_7_58_port, RESULT(57) => 
                           A_pos_shifted_by1_7_57_port, RESULT(56) => 
                           A_pos_shifted_by1_7_56_port, RESULT(55) => 
                           A_pos_shifted_by1_7_55_port, RESULT(54) => 
                           A_pos_shifted_by1_7_54_port, RESULT(53) => 
                           A_pos_shifted_by1_7_53_port, RESULT(52) => 
                           A_pos_shifted_by1_7_52_port, RESULT(51) => 
                           A_pos_shifted_by1_7_51_port, RESULT(50) => 
                           A_pos_shifted_by1_7_50_port, RESULT(49) => 
                           A_pos_shifted_by1_7_49_port, RESULT(48) => 
                           A_pos_shifted_by1_7_48_port, RESULT(47) => 
                           A_pos_shifted_by1_7_47_port, RESULT(46) => 
                           A_pos_shifted_by1_7_46_port, RESULT(45) => 
                           A_pos_shifted_by1_7_45_port, RESULT(44) => 
                           A_pos_shifted_by1_7_44_port, RESULT(43) => 
                           A_pos_shifted_by1_7_43_port, RESULT(42) => 
                           A_pos_shifted_by1_7_42_port, RESULT(41) => 
                           A_pos_shifted_by1_7_41_port, RESULT(40) => 
                           A_pos_shifted_by1_7_40_port, RESULT(39) => 
                           A_pos_shifted_by1_7_39_port, RESULT(38) => 
                           A_pos_shifted_by1_7_38_port, RESULT(37) => 
                           A_pos_shifted_by1_7_37_port, RESULT(36) => 
                           A_pos_shifted_by1_7_36_port, RESULT(35) => 
                           A_pos_shifted_by1_7_35_port, RESULT(34) => 
                           A_pos_shifted_by1_7_34_port, RESULT(33) => 
                           A_pos_shifted_by1_7_33_port, RESULT(32) => 
                           A_pos_shifted_by1_7_32_port, RESULT(31) => 
                           A_pos_shifted_by1_7_31_port, RESULT(30) => 
                           A_pos_shifted_by1_7_30_port, RESULT(29) => 
                           A_pos_shifted_by1_7_29_port, RESULT(28) => 
                           A_pos_shifted_by1_7_28_port, RESULT(27) => 
                           A_pos_shifted_by1_7_27_port, RESULT(26) => 
                           A_pos_shifted_by1_7_26_port, RESULT(25) => 
                           A_pos_shifted_by1_7_25_port, RESULT(24) => 
                           A_pos_shifted_by1_7_24_port, RESULT(23) => 
                           A_pos_shifted_by1_7_23_port, RESULT(22) => 
                           A_pos_shifted_by1_7_22_port, RESULT(21) => 
                           A_pos_shifted_by1_7_21_port, RESULT(20) => 
                           A_pos_shifted_by1_7_20_port, RESULT(19) => 
                           A_pos_shifted_by1_7_19_port, RESULT(18) => 
                           A_pos_shifted_by1_7_18_port, RESULT(17) => 
                           A_pos_shifted_by1_7_17_port, RESULT(16) => 
                           A_pos_shifted_by1_7_16_port, RESULT(15) => 
                           A_pos_shifted_by1_7_15_port, RESULT(14) => 
                           A_pos_shifted_by1_7_14_port, RESULT(13) => 
                           A_pos_shifted_by1_7_13_port, RESULT(12) => 
                           A_pos_shifted_by1_7_12_port, RESULT(11) => 
                           A_pos_shifted_by1_7_11_port, RESULT(10) => 
                           A_pos_shifted_by1_7_10_port, RESULT(9) => 
                           A_pos_shifted_by1_7_9_port, RESULT(8) => 
                           A_pos_shifted_by1_7_8_port, RESULT(7) => 
                           A_pos_shifted_by1_7_7_port, RESULT(6) => 
                           A_pos_shifted_by1_7_6_port, RESULT(5) => 
                           A_pos_shifted_by1_7_5_port, RESULT(4) => 
                           A_pos_shifted_by1_7_4_port, RESULT(3) => 
                           A_pos_shifted_by1_7_3_port, RESULT(2) => 
                           A_pos_shifted_by1_7_2_port, RESULT(1) => 
                           A_pos_shifted_by1_7_1_port, RESULT(0) => n_1083);
   SHIFTERi_8 : Shifter_NBIT64_24 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_7_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_7_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_7_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_7_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_7_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_7_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_7_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_7_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_7_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_7_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_7_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_7_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_7_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_7_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_7_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_7_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_7_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_7_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_7_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_7_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_7_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_7_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_7_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_7_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_7_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_7_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_7_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_7_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_7_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_7_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_7_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_7_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_7_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_7_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_7_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_7_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_7_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_7_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_7_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_7_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_7_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_7_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_7_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_7_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_7_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_7_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_7_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_7_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_7_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_7_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_7_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_7_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_7_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_7_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_7_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_7_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_7_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_7_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_7_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_7_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_7_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_7_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_7_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_7_0_port, RESULT(127) => 
                           A_pos_shifted_by2_8_63_port, RESULT(126) => 
                           A_pos_shifted_by2_8_62_port, RESULT(125) => 
                           A_pos_shifted_by2_8_61_port, RESULT(124) => 
                           A_pos_shifted_by2_8_60_port, RESULT(123) => 
                           A_pos_shifted_by2_8_59_port, RESULT(122) => 
                           A_pos_shifted_by2_8_58_port, RESULT(121) => 
                           A_pos_shifted_by2_8_57_port, RESULT(120) => 
                           A_pos_shifted_by2_8_56_port, RESULT(119) => 
                           A_pos_shifted_by2_8_55_port, RESULT(118) => 
                           A_pos_shifted_by2_8_54_port, RESULT(117) => 
                           A_pos_shifted_by2_8_53_port, RESULT(116) => 
                           A_pos_shifted_by2_8_52_port, RESULT(115) => 
                           A_pos_shifted_by2_8_51_port, RESULT(114) => 
                           A_pos_shifted_by2_8_50_port, RESULT(113) => 
                           A_pos_shifted_by2_8_49_port, RESULT(112) => 
                           A_pos_shifted_by2_8_48_port, RESULT(111) => 
                           A_pos_shifted_by2_8_47_port, RESULT(110) => 
                           A_pos_shifted_by2_8_46_port, RESULT(109) => 
                           A_pos_shifted_by2_8_45_port, RESULT(108) => 
                           A_pos_shifted_by2_8_44_port, RESULT(107) => 
                           A_pos_shifted_by2_8_43_port, RESULT(106) => 
                           A_pos_shifted_by2_8_42_port, RESULT(105) => 
                           A_pos_shifted_by2_8_41_port, RESULT(104) => 
                           A_pos_shifted_by2_8_40_port, RESULT(103) => 
                           A_pos_shifted_by2_8_39_port, RESULT(102) => 
                           A_pos_shifted_by2_8_38_port, RESULT(101) => 
                           A_pos_shifted_by2_8_37_port, RESULT(100) => 
                           A_pos_shifted_by2_8_36_port, RESULT(99) => 
                           A_pos_shifted_by2_8_35_port, RESULT(98) => 
                           A_pos_shifted_by2_8_34_port, RESULT(97) => 
                           A_pos_shifted_by2_8_33_port, RESULT(96) => 
                           A_pos_shifted_by2_8_32_port, RESULT(95) => 
                           A_pos_shifted_by2_8_31_port, RESULT(94) => 
                           A_pos_shifted_by2_8_30_port, RESULT(93) => 
                           A_pos_shifted_by2_8_29_port, RESULT(92) => 
                           A_pos_shifted_by2_8_28_port, RESULT(91) => 
                           A_pos_shifted_by2_8_27_port, RESULT(90) => 
                           A_pos_shifted_by2_8_26_port, RESULT(89) => 
                           A_pos_shifted_by2_8_25_port, RESULT(88) => 
                           A_pos_shifted_by2_8_24_port, RESULT(87) => 
                           A_pos_shifted_by2_8_23_port, RESULT(86) => 
                           A_pos_shifted_by2_8_22_port, RESULT(85) => 
                           A_pos_shifted_by2_8_21_port, RESULT(84) => 
                           A_pos_shifted_by2_8_20_port, RESULT(83) => 
                           A_pos_shifted_by2_8_19_port, RESULT(82) => 
                           A_pos_shifted_by2_8_18_port, RESULT(81) => 
                           A_pos_shifted_by2_8_17_port, RESULT(80) => 
                           A_pos_shifted_by2_8_16_port, RESULT(79) => 
                           A_pos_shifted_by2_8_15_port, RESULT(78) => 
                           A_pos_shifted_by2_8_14_port, RESULT(77) => 
                           A_pos_shifted_by2_8_13_port, RESULT(76) => 
                           A_pos_shifted_by2_8_12_port, RESULT(75) => 
                           A_pos_shifted_by2_8_11_port, RESULT(74) => 
                           A_pos_shifted_by2_8_10_port, RESULT(73) => 
                           A_pos_shifted_by2_8_9_port, RESULT(72) => 
                           A_pos_shifted_by2_8_8_port, RESULT(71) => 
                           A_pos_shifted_by2_8_7_port, RESULT(70) => 
                           A_pos_shifted_by2_8_6_port, RESULT(69) => 
                           A_pos_shifted_by2_8_5_port, RESULT(68) => 
                           A_pos_shifted_by2_8_4_port, RESULT(67) => 
                           A_pos_shifted_by2_8_3_port, RESULT(66) => 
                           A_pos_shifted_by2_8_2_port, RESULT(65) => n_1084, 
                           RESULT(64) => n_1085, RESULT(63) => 
                           A_pos_shifted_by1_8_63_port, RESULT(62) => 
                           A_pos_shifted_by1_8_62_port, RESULT(61) => 
                           A_pos_shifted_by1_8_61_port, RESULT(60) => 
                           A_pos_shifted_by1_8_60_port, RESULT(59) => 
                           A_pos_shifted_by1_8_59_port, RESULT(58) => 
                           A_pos_shifted_by1_8_58_port, RESULT(57) => 
                           A_pos_shifted_by1_8_57_port, RESULT(56) => 
                           A_pos_shifted_by1_8_56_port, RESULT(55) => 
                           A_pos_shifted_by1_8_55_port, RESULT(54) => 
                           A_pos_shifted_by1_8_54_port, RESULT(53) => 
                           A_pos_shifted_by1_8_53_port, RESULT(52) => 
                           A_pos_shifted_by1_8_52_port, RESULT(51) => 
                           A_pos_shifted_by1_8_51_port, RESULT(50) => 
                           A_pos_shifted_by1_8_50_port, RESULT(49) => 
                           A_pos_shifted_by1_8_49_port, RESULT(48) => 
                           A_pos_shifted_by1_8_48_port, RESULT(47) => 
                           A_pos_shifted_by1_8_47_port, RESULT(46) => 
                           A_pos_shifted_by1_8_46_port, RESULT(45) => 
                           A_pos_shifted_by1_8_45_port, RESULT(44) => 
                           A_pos_shifted_by1_8_44_port, RESULT(43) => 
                           A_pos_shifted_by1_8_43_port, RESULT(42) => 
                           A_pos_shifted_by1_8_42_port, RESULT(41) => 
                           A_pos_shifted_by1_8_41_port, RESULT(40) => 
                           A_pos_shifted_by1_8_40_port, RESULT(39) => 
                           A_pos_shifted_by1_8_39_port, RESULT(38) => 
                           A_pos_shifted_by1_8_38_port, RESULT(37) => 
                           A_pos_shifted_by1_8_37_port, RESULT(36) => 
                           A_pos_shifted_by1_8_36_port, RESULT(35) => 
                           A_pos_shifted_by1_8_35_port, RESULT(34) => 
                           A_pos_shifted_by1_8_34_port, RESULT(33) => 
                           A_pos_shifted_by1_8_33_port, RESULT(32) => 
                           A_pos_shifted_by1_8_32_port, RESULT(31) => 
                           A_pos_shifted_by1_8_31_port, RESULT(30) => 
                           A_pos_shifted_by1_8_30_port, RESULT(29) => 
                           A_pos_shifted_by1_8_29_port, RESULT(28) => 
                           A_pos_shifted_by1_8_28_port, RESULT(27) => 
                           A_pos_shifted_by1_8_27_port, RESULT(26) => 
                           A_pos_shifted_by1_8_26_port, RESULT(25) => 
                           A_pos_shifted_by1_8_25_port, RESULT(24) => 
                           A_pos_shifted_by1_8_24_port, RESULT(23) => 
                           A_pos_shifted_by1_8_23_port, RESULT(22) => 
                           A_pos_shifted_by1_8_22_port, RESULT(21) => 
                           A_pos_shifted_by1_8_21_port, RESULT(20) => 
                           A_pos_shifted_by1_8_20_port, RESULT(19) => 
                           A_pos_shifted_by1_8_19_port, RESULT(18) => 
                           A_pos_shifted_by1_8_18_port, RESULT(17) => 
                           A_pos_shifted_by1_8_17_port, RESULT(16) => 
                           A_pos_shifted_by1_8_16_port, RESULT(15) => 
                           A_pos_shifted_by1_8_15_port, RESULT(14) => 
                           A_pos_shifted_by1_8_14_port, RESULT(13) => 
                           A_pos_shifted_by1_8_13_port, RESULT(12) => 
                           A_pos_shifted_by1_8_12_port, RESULT(11) => 
                           A_pos_shifted_by1_8_11_port, RESULT(10) => 
                           A_pos_shifted_by1_8_10_port, RESULT(9) => 
                           A_pos_shifted_by1_8_9_port, RESULT(8) => 
                           A_pos_shifted_by1_8_8_port, RESULT(7) => 
                           A_pos_shifted_by1_8_7_port, RESULT(6) => 
                           A_pos_shifted_by1_8_6_port, RESULT(5) => 
                           A_pos_shifted_by1_8_5_port, RESULT(4) => 
                           A_pos_shifted_by1_8_4_port, RESULT(3) => 
                           A_pos_shifted_by1_8_3_port, RESULT(2) => 
                           A_pos_shifted_by1_8_2_port, RESULT(1) => 
                           A_pos_shifted_by1_8_1_port, RESULT(0) => n_1086);
   SHIFTERi_9 : Shifter_NBIT64_23 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_8_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_8_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_8_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_8_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_8_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_8_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_8_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_8_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_8_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_8_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_8_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_8_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_8_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_8_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_8_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_8_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_8_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_8_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_8_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_8_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_8_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_8_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_8_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_8_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_8_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_8_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_8_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_8_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_8_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_8_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_8_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_8_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_8_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_8_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_8_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_8_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_8_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_8_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_8_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_8_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_8_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_8_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_8_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_8_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_8_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_8_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_8_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_8_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_8_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_8_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_8_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_8_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_8_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_8_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_8_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_8_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_8_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_8_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_8_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_8_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_8_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_8_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_8_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_8_0_port, RESULT(127) => 
                           A_pos_shifted_by2_9_63_port, RESULT(126) => 
                           A_pos_shifted_by2_9_62_port, RESULT(125) => 
                           A_pos_shifted_by2_9_61_port, RESULT(124) => 
                           A_pos_shifted_by2_9_60_port, RESULT(123) => 
                           A_pos_shifted_by2_9_59_port, RESULT(122) => 
                           A_pos_shifted_by2_9_58_port, RESULT(121) => 
                           A_pos_shifted_by2_9_57_port, RESULT(120) => 
                           A_pos_shifted_by2_9_56_port, RESULT(119) => 
                           A_pos_shifted_by2_9_55_port, RESULT(118) => 
                           A_pos_shifted_by2_9_54_port, RESULT(117) => 
                           A_pos_shifted_by2_9_53_port, RESULT(116) => 
                           A_pos_shifted_by2_9_52_port, RESULT(115) => 
                           A_pos_shifted_by2_9_51_port, RESULT(114) => 
                           A_pos_shifted_by2_9_50_port, RESULT(113) => 
                           A_pos_shifted_by2_9_49_port, RESULT(112) => 
                           A_pos_shifted_by2_9_48_port, RESULT(111) => 
                           A_pos_shifted_by2_9_47_port, RESULT(110) => 
                           A_pos_shifted_by2_9_46_port, RESULT(109) => 
                           A_pos_shifted_by2_9_45_port, RESULT(108) => 
                           A_pos_shifted_by2_9_44_port, RESULT(107) => 
                           A_pos_shifted_by2_9_43_port, RESULT(106) => 
                           A_pos_shifted_by2_9_42_port, RESULT(105) => 
                           A_pos_shifted_by2_9_41_port, RESULT(104) => 
                           A_pos_shifted_by2_9_40_port, RESULT(103) => 
                           A_pos_shifted_by2_9_39_port, RESULT(102) => 
                           A_pos_shifted_by2_9_38_port, RESULT(101) => 
                           A_pos_shifted_by2_9_37_port, RESULT(100) => 
                           A_pos_shifted_by2_9_36_port, RESULT(99) => 
                           A_pos_shifted_by2_9_35_port, RESULT(98) => 
                           A_pos_shifted_by2_9_34_port, RESULT(97) => 
                           A_pos_shifted_by2_9_33_port, RESULT(96) => 
                           A_pos_shifted_by2_9_32_port, RESULT(95) => 
                           A_pos_shifted_by2_9_31_port, RESULT(94) => 
                           A_pos_shifted_by2_9_30_port, RESULT(93) => 
                           A_pos_shifted_by2_9_29_port, RESULT(92) => 
                           A_pos_shifted_by2_9_28_port, RESULT(91) => 
                           A_pos_shifted_by2_9_27_port, RESULT(90) => 
                           A_pos_shifted_by2_9_26_port, RESULT(89) => 
                           A_pos_shifted_by2_9_25_port, RESULT(88) => 
                           A_pos_shifted_by2_9_24_port, RESULT(87) => 
                           A_pos_shifted_by2_9_23_port, RESULT(86) => 
                           A_pos_shifted_by2_9_22_port, RESULT(85) => 
                           A_pos_shifted_by2_9_21_port, RESULT(84) => 
                           A_pos_shifted_by2_9_20_port, RESULT(83) => 
                           A_pos_shifted_by2_9_19_port, RESULT(82) => 
                           A_pos_shifted_by2_9_18_port, RESULT(81) => 
                           A_pos_shifted_by2_9_17_port, RESULT(80) => 
                           A_pos_shifted_by2_9_16_port, RESULT(79) => 
                           A_pos_shifted_by2_9_15_port, RESULT(78) => 
                           A_pos_shifted_by2_9_14_port, RESULT(77) => 
                           A_pos_shifted_by2_9_13_port, RESULT(76) => 
                           A_pos_shifted_by2_9_12_port, RESULT(75) => 
                           A_pos_shifted_by2_9_11_port, RESULT(74) => 
                           A_pos_shifted_by2_9_10_port, RESULT(73) => 
                           A_pos_shifted_by2_9_9_port, RESULT(72) => 
                           A_pos_shifted_by2_9_8_port, RESULT(71) => 
                           A_pos_shifted_by2_9_7_port, RESULT(70) => 
                           A_pos_shifted_by2_9_6_port, RESULT(69) => 
                           A_pos_shifted_by2_9_5_port, RESULT(68) => 
                           A_pos_shifted_by2_9_4_port, RESULT(67) => 
                           A_pos_shifted_by2_9_3_port, RESULT(66) => 
                           A_pos_shifted_by2_9_2_port, RESULT(65) => n_1087, 
                           RESULT(64) => n_1088, RESULT(63) => 
                           A_pos_shifted_by1_9_63_port, RESULT(62) => 
                           A_pos_shifted_by1_9_62_port, RESULT(61) => 
                           A_pos_shifted_by1_9_61_port, RESULT(60) => 
                           A_pos_shifted_by1_9_60_port, RESULT(59) => 
                           A_pos_shifted_by1_9_59_port, RESULT(58) => 
                           A_pos_shifted_by1_9_58_port, RESULT(57) => 
                           A_pos_shifted_by1_9_57_port, RESULT(56) => 
                           A_pos_shifted_by1_9_56_port, RESULT(55) => 
                           A_pos_shifted_by1_9_55_port, RESULT(54) => 
                           A_pos_shifted_by1_9_54_port, RESULT(53) => 
                           A_pos_shifted_by1_9_53_port, RESULT(52) => 
                           A_pos_shifted_by1_9_52_port, RESULT(51) => 
                           A_pos_shifted_by1_9_51_port, RESULT(50) => 
                           A_pos_shifted_by1_9_50_port, RESULT(49) => 
                           A_pos_shifted_by1_9_49_port, RESULT(48) => 
                           A_pos_shifted_by1_9_48_port, RESULT(47) => 
                           A_pos_shifted_by1_9_47_port, RESULT(46) => 
                           A_pos_shifted_by1_9_46_port, RESULT(45) => 
                           A_pos_shifted_by1_9_45_port, RESULT(44) => 
                           A_pos_shifted_by1_9_44_port, RESULT(43) => 
                           A_pos_shifted_by1_9_43_port, RESULT(42) => 
                           A_pos_shifted_by1_9_42_port, RESULT(41) => 
                           A_pos_shifted_by1_9_41_port, RESULT(40) => 
                           A_pos_shifted_by1_9_40_port, RESULT(39) => 
                           A_pos_shifted_by1_9_39_port, RESULT(38) => 
                           A_pos_shifted_by1_9_38_port, RESULT(37) => 
                           A_pos_shifted_by1_9_37_port, RESULT(36) => 
                           A_pos_shifted_by1_9_36_port, RESULT(35) => 
                           A_pos_shifted_by1_9_35_port, RESULT(34) => 
                           A_pos_shifted_by1_9_34_port, RESULT(33) => 
                           A_pos_shifted_by1_9_33_port, RESULT(32) => 
                           A_pos_shifted_by1_9_32_port, RESULT(31) => 
                           A_pos_shifted_by1_9_31_port, RESULT(30) => 
                           A_pos_shifted_by1_9_30_port, RESULT(29) => 
                           A_pos_shifted_by1_9_29_port, RESULT(28) => 
                           A_pos_shifted_by1_9_28_port, RESULT(27) => 
                           A_pos_shifted_by1_9_27_port, RESULT(26) => 
                           A_pos_shifted_by1_9_26_port, RESULT(25) => 
                           A_pos_shifted_by1_9_25_port, RESULT(24) => 
                           A_pos_shifted_by1_9_24_port, RESULT(23) => 
                           A_pos_shifted_by1_9_23_port, RESULT(22) => 
                           A_pos_shifted_by1_9_22_port, RESULT(21) => 
                           A_pos_shifted_by1_9_21_port, RESULT(20) => 
                           A_pos_shifted_by1_9_20_port, RESULT(19) => 
                           A_pos_shifted_by1_9_19_port, RESULT(18) => 
                           A_pos_shifted_by1_9_18_port, RESULT(17) => 
                           A_pos_shifted_by1_9_17_port, RESULT(16) => 
                           A_pos_shifted_by1_9_16_port, RESULT(15) => 
                           A_pos_shifted_by1_9_15_port, RESULT(14) => 
                           A_pos_shifted_by1_9_14_port, RESULT(13) => 
                           A_pos_shifted_by1_9_13_port, RESULT(12) => 
                           A_pos_shifted_by1_9_12_port, RESULT(11) => 
                           A_pos_shifted_by1_9_11_port, RESULT(10) => 
                           A_pos_shifted_by1_9_10_port, RESULT(9) => 
                           A_pos_shifted_by1_9_9_port, RESULT(8) => 
                           A_pos_shifted_by1_9_8_port, RESULT(7) => 
                           A_pos_shifted_by1_9_7_port, RESULT(6) => 
                           A_pos_shifted_by1_9_6_port, RESULT(5) => 
                           A_pos_shifted_by1_9_5_port, RESULT(4) => 
                           A_pos_shifted_by1_9_4_port, RESULT(3) => 
                           A_pos_shifted_by1_9_3_port, RESULT(2) => 
                           A_pos_shifted_by1_9_2_port, RESULT(1) => 
                           A_pos_shifted_by1_9_1_port, RESULT(0) => n_1089);
   SHIFTERi_10 : Shifter_NBIT64_22 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_9_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_9_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_9_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_9_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_9_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_9_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_9_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_9_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_9_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_9_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_9_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_9_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_9_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_9_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_9_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_9_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_9_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_9_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_9_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_9_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_9_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_9_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_9_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_9_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_9_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_9_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_9_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_9_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_9_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_9_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_9_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_9_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_9_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_9_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_9_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_9_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_9_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_9_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_9_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_9_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_9_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_9_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_9_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_9_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_9_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_9_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_9_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_9_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_9_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_9_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_9_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_9_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_9_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_9_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_9_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_9_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_9_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_9_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_9_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_9_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_9_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_9_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_9_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_9_0_port, RESULT(127) => 
                           A_pos_shifted_by2_10_63_port, RESULT(126) => 
                           A_pos_shifted_by2_10_62_port, RESULT(125) => 
                           A_pos_shifted_by2_10_61_port, RESULT(124) => 
                           A_pos_shifted_by2_10_60_port, RESULT(123) => 
                           A_pos_shifted_by2_10_59_port, RESULT(122) => 
                           A_pos_shifted_by2_10_58_port, RESULT(121) => 
                           A_pos_shifted_by2_10_57_port, RESULT(120) => 
                           A_pos_shifted_by2_10_56_port, RESULT(119) => 
                           A_pos_shifted_by2_10_55_port, RESULT(118) => 
                           A_pos_shifted_by2_10_54_port, RESULT(117) => 
                           A_pos_shifted_by2_10_53_port, RESULT(116) => 
                           A_pos_shifted_by2_10_52_port, RESULT(115) => 
                           A_pos_shifted_by2_10_51_port, RESULT(114) => 
                           A_pos_shifted_by2_10_50_port, RESULT(113) => 
                           A_pos_shifted_by2_10_49_port, RESULT(112) => 
                           A_pos_shifted_by2_10_48_port, RESULT(111) => 
                           A_pos_shifted_by2_10_47_port, RESULT(110) => 
                           A_pos_shifted_by2_10_46_port, RESULT(109) => 
                           A_pos_shifted_by2_10_45_port, RESULT(108) => 
                           A_pos_shifted_by2_10_44_port, RESULT(107) => 
                           A_pos_shifted_by2_10_43_port, RESULT(106) => 
                           A_pos_shifted_by2_10_42_port, RESULT(105) => 
                           A_pos_shifted_by2_10_41_port, RESULT(104) => 
                           A_pos_shifted_by2_10_40_port, RESULT(103) => 
                           A_pos_shifted_by2_10_39_port, RESULT(102) => 
                           A_pos_shifted_by2_10_38_port, RESULT(101) => 
                           A_pos_shifted_by2_10_37_port, RESULT(100) => 
                           A_pos_shifted_by2_10_36_port, RESULT(99) => 
                           A_pos_shifted_by2_10_35_port, RESULT(98) => 
                           A_pos_shifted_by2_10_34_port, RESULT(97) => 
                           A_pos_shifted_by2_10_33_port, RESULT(96) => 
                           A_pos_shifted_by2_10_32_port, RESULT(95) => 
                           A_pos_shifted_by2_10_31_port, RESULT(94) => 
                           A_pos_shifted_by2_10_30_port, RESULT(93) => 
                           A_pos_shifted_by2_10_29_port, RESULT(92) => 
                           A_pos_shifted_by2_10_28_port, RESULT(91) => 
                           A_pos_shifted_by2_10_27_port, RESULT(90) => 
                           A_pos_shifted_by2_10_26_port, RESULT(89) => 
                           A_pos_shifted_by2_10_25_port, RESULT(88) => 
                           A_pos_shifted_by2_10_24_port, RESULT(87) => 
                           A_pos_shifted_by2_10_23_port, RESULT(86) => 
                           A_pos_shifted_by2_10_22_port, RESULT(85) => 
                           A_pos_shifted_by2_10_21_port, RESULT(84) => 
                           A_pos_shifted_by2_10_20_port, RESULT(83) => 
                           A_pos_shifted_by2_10_19_port, RESULT(82) => 
                           A_pos_shifted_by2_10_18_port, RESULT(81) => 
                           A_pos_shifted_by2_10_17_port, RESULT(80) => 
                           A_pos_shifted_by2_10_16_port, RESULT(79) => 
                           A_pos_shifted_by2_10_15_port, RESULT(78) => 
                           A_pos_shifted_by2_10_14_port, RESULT(77) => 
                           A_pos_shifted_by2_10_13_port, RESULT(76) => 
                           A_pos_shifted_by2_10_12_port, RESULT(75) => 
                           A_pos_shifted_by2_10_11_port, RESULT(74) => 
                           A_pos_shifted_by2_10_10_port, RESULT(73) => 
                           A_pos_shifted_by2_10_9_port, RESULT(72) => 
                           A_pos_shifted_by2_10_8_port, RESULT(71) => 
                           A_pos_shifted_by2_10_7_port, RESULT(70) => 
                           A_pos_shifted_by2_10_6_port, RESULT(69) => 
                           A_pos_shifted_by2_10_5_port, RESULT(68) => 
                           A_pos_shifted_by2_10_4_port, RESULT(67) => 
                           A_pos_shifted_by2_10_3_port, RESULT(66) => 
                           A_pos_shifted_by2_10_2_port, RESULT(65) => n_1090, 
                           RESULT(64) => n_1091, RESULT(63) => 
                           A_pos_shifted_by1_10_63_port, RESULT(62) => 
                           A_pos_shifted_by1_10_62_port, RESULT(61) => 
                           A_pos_shifted_by1_10_61_port, RESULT(60) => 
                           A_pos_shifted_by1_10_60_port, RESULT(59) => 
                           A_pos_shifted_by1_10_59_port, RESULT(58) => 
                           A_pos_shifted_by1_10_58_port, RESULT(57) => 
                           A_pos_shifted_by1_10_57_port, RESULT(56) => 
                           A_pos_shifted_by1_10_56_port, RESULT(55) => 
                           A_pos_shifted_by1_10_55_port, RESULT(54) => 
                           A_pos_shifted_by1_10_54_port, RESULT(53) => 
                           A_pos_shifted_by1_10_53_port, RESULT(52) => 
                           A_pos_shifted_by1_10_52_port, RESULT(51) => 
                           A_pos_shifted_by1_10_51_port, RESULT(50) => 
                           A_pos_shifted_by1_10_50_port, RESULT(49) => 
                           A_pos_shifted_by1_10_49_port, RESULT(48) => 
                           A_pos_shifted_by1_10_48_port, RESULT(47) => 
                           A_pos_shifted_by1_10_47_port, RESULT(46) => 
                           A_pos_shifted_by1_10_46_port, RESULT(45) => 
                           A_pos_shifted_by1_10_45_port, RESULT(44) => 
                           A_pos_shifted_by1_10_44_port, RESULT(43) => 
                           A_pos_shifted_by1_10_43_port, RESULT(42) => 
                           A_pos_shifted_by1_10_42_port, RESULT(41) => 
                           A_pos_shifted_by1_10_41_port, RESULT(40) => 
                           A_pos_shifted_by1_10_40_port, RESULT(39) => 
                           A_pos_shifted_by1_10_39_port, RESULT(38) => 
                           A_pos_shifted_by1_10_38_port, RESULT(37) => 
                           A_pos_shifted_by1_10_37_port, RESULT(36) => 
                           A_pos_shifted_by1_10_36_port, RESULT(35) => 
                           A_pos_shifted_by1_10_35_port, RESULT(34) => 
                           A_pos_shifted_by1_10_34_port, RESULT(33) => 
                           A_pos_shifted_by1_10_33_port, RESULT(32) => 
                           A_pos_shifted_by1_10_32_port, RESULT(31) => 
                           A_pos_shifted_by1_10_31_port, RESULT(30) => 
                           A_pos_shifted_by1_10_30_port, RESULT(29) => 
                           A_pos_shifted_by1_10_29_port, RESULT(28) => 
                           A_pos_shifted_by1_10_28_port, RESULT(27) => 
                           A_pos_shifted_by1_10_27_port, RESULT(26) => 
                           A_pos_shifted_by1_10_26_port, RESULT(25) => 
                           A_pos_shifted_by1_10_25_port, RESULT(24) => 
                           A_pos_shifted_by1_10_24_port, RESULT(23) => 
                           A_pos_shifted_by1_10_23_port, RESULT(22) => 
                           A_pos_shifted_by1_10_22_port, RESULT(21) => 
                           A_pos_shifted_by1_10_21_port, RESULT(20) => 
                           A_pos_shifted_by1_10_20_port, RESULT(19) => 
                           A_pos_shifted_by1_10_19_port, RESULT(18) => 
                           A_pos_shifted_by1_10_18_port, RESULT(17) => 
                           A_pos_shifted_by1_10_17_port, RESULT(16) => 
                           A_pos_shifted_by1_10_16_port, RESULT(15) => 
                           A_pos_shifted_by1_10_15_port, RESULT(14) => 
                           A_pos_shifted_by1_10_14_port, RESULT(13) => 
                           A_pos_shifted_by1_10_13_port, RESULT(12) => 
                           A_pos_shifted_by1_10_12_port, RESULT(11) => 
                           A_pos_shifted_by1_10_11_port, RESULT(10) => 
                           A_pos_shifted_by1_10_10_port, RESULT(9) => 
                           A_pos_shifted_by1_10_9_port, RESULT(8) => 
                           A_pos_shifted_by1_10_8_port, RESULT(7) => 
                           A_pos_shifted_by1_10_7_port, RESULT(6) => 
                           A_pos_shifted_by1_10_6_port, RESULT(5) => 
                           A_pos_shifted_by1_10_5_port, RESULT(4) => 
                           A_pos_shifted_by1_10_4_port, RESULT(3) => 
                           A_pos_shifted_by1_10_3_port, RESULT(2) => 
                           A_pos_shifted_by1_10_2_port, RESULT(1) => 
                           A_pos_shifted_by1_10_1_port, RESULT(0) => n_1092);
   SHIFTERi_11 : Shifter_NBIT64_21 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_10_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_10_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_10_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_10_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_10_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_10_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_10_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_10_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_10_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_10_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_10_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_10_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_10_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_10_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_10_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_10_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_10_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_10_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_10_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_10_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_10_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_10_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_10_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_10_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_10_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_10_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_10_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_10_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_10_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_10_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_10_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_10_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_10_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_10_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_10_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_10_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_10_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_10_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_10_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_10_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_10_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_10_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_10_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_10_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_10_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_10_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_10_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_10_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_10_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_10_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_10_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_10_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_10_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_10_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_10_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_10_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_10_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_10_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_10_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_10_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_10_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_10_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_10_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_10_0_port, RESULT(127) => 
                           A_pos_shifted_by2_11_63_port, RESULT(126) => 
                           A_pos_shifted_by2_11_62_port, RESULT(125) => 
                           A_pos_shifted_by2_11_61_port, RESULT(124) => 
                           A_pos_shifted_by2_11_60_port, RESULT(123) => 
                           A_pos_shifted_by2_11_59_port, RESULT(122) => 
                           A_pos_shifted_by2_11_58_port, RESULT(121) => 
                           A_pos_shifted_by2_11_57_port, RESULT(120) => 
                           A_pos_shifted_by2_11_56_port, RESULT(119) => 
                           A_pos_shifted_by2_11_55_port, RESULT(118) => 
                           A_pos_shifted_by2_11_54_port, RESULT(117) => 
                           A_pos_shifted_by2_11_53_port, RESULT(116) => 
                           A_pos_shifted_by2_11_52_port, RESULT(115) => 
                           A_pos_shifted_by2_11_51_port, RESULT(114) => 
                           A_pos_shifted_by2_11_50_port, RESULT(113) => 
                           A_pos_shifted_by2_11_49_port, RESULT(112) => 
                           A_pos_shifted_by2_11_48_port, RESULT(111) => 
                           A_pos_shifted_by2_11_47_port, RESULT(110) => 
                           A_pos_shifted_by2_11_46_port, RESULT(109) => 
                           A_pos_shifted_by2_11_45_port, RESULT(108) => 
                           A_pos_shifted_by2_11_44_port, RESULT(107) => 
                           A_pos_shifted_by2_11_43_port, RESULT(106) => 
                           A_pos_shifted_by2_11_42_port, RESULT(105) => 
                           A_pos_shifted_by2_11_41_port, RESULT(104) => 
                           A_pos_shifted_by2_11_40_port, RESULT(103) => 
                           A_pos_shifted_by2_11_39_port, RESULT(102) => 
                           A_pos_shifted_by2_11_38_port, RESULT(101) => 
                           A_pos_shifted_by2_11_37_port, RESULT(100) => 
                           A_pos_shifted_by2_11_36_port, RESULT(99) => 
                           A_pos_shifted_by2_11_35_port, RESULT(98) => 
                           A_pos_shifted_by2_11_34_port, RESULT(97) => 
                           A_pos_shifted_by2_11_33_port, RESULT(96) => 
                           A_pos_shifted_by2_11_32_port, RESULT(95) => 
                           A_pos_shifted_by2_11_31_port, RESULT(94) => 
                           A_pos_shifted_by2_11_30_port, RESULT(93) => 
                           A_pos_shifted_by2_11_29_port, RESULT(92) => 
                           A_pos_shifted_by2_11_28_port, RESULT(91) => 
                           A_pos_shifted_by2_11_27_port, RESULT(90) => 
                           A_pos_shifted_by2_11_26_port, RESULT(89) => 
                           A_pos_shifted_by2_11_25_port, RESULT(88) => 
                           A_pos_shifted_by2_11_24_port, RESULT(87) => 
                           A_pos_shifted_by2_11_23_port, RESULT(86) => 
                           A_pos_shifted_by2_11_22_port, RESULT(85) => 
                           A_pos_shifted_by2_11_21_port, RESULT(84) => 
                           A_pos_shifted_by2_11_20_port, RESULT(83) => 
                           A_pos_shifted_by2_11_19_port, RESULT(82) => 
                           A_pos_shifted_by2_11_18_port, RESULT(81) => 
                           A_pos_shifted_by2_11_17_port, RESULT(80) => 
                           A_pos_shifted_by2_11_16_port, RESULT(79) => 
                           A_pos_shifted_by2_11_15_port, RESULT(78) => 
                           A_pos_shifted_by2_11_14_port, RESULT(77) => 
                           A_pos_shifted_by2_11_13_port, RESULT(76) => 
                           A_pos_shifted_by2_11_12_port, RESULT(75) => 
                           A_pos_shifted_by2_11_11_port, RESULT(74) => 
                           A_pos_shifted_by2_11_10_port, RESULT(73) => 
                           A_pos_shifted_by2_11_9_port, RESULT(72) => 
                           A_pos_shifted_by2_11_8_port, RESULT(71) => 
                           A_pos_shifted_by2_11_7_port, RESULT(70) => 
                           A_pos_shifted_by2_11_6_port, RESULT(69) => 
                           A_pos_shifted_by2_11_5_port, RESULT(68) => 
                           A_pos_shifted_by2_11_4_port, RESULT(67) => 
                           A_pos_shifted_by2_11_3_port, RESULT(66) => 
                           A_pos_shifted_by2_11_2_port, RESULT(65) => n_1093, 
                           RESULT(64) => n_1094, RESULT(63) => 
                           A_pos_shifted_by1_11_63_port, RESULT(62) => 
                           A_pos_shifted_by1_11_62_port, RESULT(61) => 
                           A_pos_shifted_by1_11_61_port, RESULT(60) => 
                           A_pos_shifted_by1_11_60_port, RESULT(59) => 
                           A_pos_shifted_by1_11_59_port, RESULT(58) => 
                           A_pos_shifted_by1_11_58_port, RESULT(57) => 
                           A_pos_shifted_by1_11_57_port, RESULT(56) => 
                           A_pos_shifted_by1_11_56_port, RESULT(55) => 
                           A_pos_shifted_by1_11_55_port, RESULT(54) => 
                           A_pos_shifted_by1_11_54_port, RESULT(53) => 
                           A_pos_shifted_by1_11_53_port, RESULT(52) => 
                           A_pos_shifted_by1_11_52_port, RESULT(51) => 
                           A_pos_shifted_by1_11_51_port, RESULT(50) => 
                           A_pos_shifted_by1_11_50_port, RESULT(49) => 
                           A_pos_shifted_by1_11_49_port, RESULT(48) => 
                           A_pos_shifted_by1_11_48_port, RESULT(47) => 
                           A_pos_shifted_by1_11_47_port, RESULT(46) => 
                           A_pos_shifted_by1_11_46_port, RESULT(45) => 
                           A_pos_shifted_by1_11_45_port, RESULT(44) => 
                           A_pos_shifted_by1_11_44_port, RESULT(43) => 
                           A_pos_shifted_by1_11_43_port, RESULT(42) => 
                           A_pos_shifted_by1_11_42_port, RESULT(41) => 
                           A_pos_shifted_by1_11_41_port, RESULT(40) => 
                           A_pos_shifted_by1_11_40_port, RESULT(39) => 
                           A_pos_shifted_by1_11_39_port, RESULT(38) => 
                           A_pos_shifted_by1_11_38_port, RESULT(37) => 
                           A_pos_shifted_by1_11_37_port, RESULT(36) => 
                           A_pos_shifted_by1_11_36_port, RESULT(35) => 
                           A_pos_shifted_by1_11_35_port, RESULT(34) => 
                           A_pos_shifted_by1_11_34_port, RESULT(33) => 
                           A_pos_shifted_by1_11_33_port, RESULT(32) => 
                           A_pos_shifted_by1_11_32_port, RESULT(31) => 
                           A_pos_shifted_by1_11_31_port, RESULT(30) => 
                           A_pos_shifted_by1_11_30_port, RESULT(29) => 
                           A_pos_shifted_by1_11_29_port, RESULT(28) => 
                           A_pos_shifted_by1_11_28_port, RESULT(27) => 
                           A_pos_shifted_by1_11_27_port, RESULT(26) => 
                           A_pos_shifted_by1_11_26_port, RESULT(25) => 
                           A_pos_shifted_by1_11_25_port, RESULT(24) => 
                           A_pos_shifted_by1_11_24_port, RESULT(23) => 
                           A_pos_shifted_by1_11_23_port, RESULT(22) => 
                           A_pos_shifted_by1_11_22_port, RESULT(21) => 
                           A_pos_shifted_by1_11_21_port, RESULT(20) => 
                           A_pos_shifted_by1_11_20_port, RESULT(19) => 
                           A_pos_shifted_by1_11_19_port, RESULT(18) => 
                           A_pos_shifted_by1_11_18_port, RESULT(17) => 
                           A_pos_shifted_by1_11_17_port, RESULT(16) => 
                           A_pos_shifted_by1_11_16_port, RESULT(15) => 
                           A_pos_shifted_by1_11_15_port, RESULT(14) => 
                           A_pos_shifted_by1_11_14_port, RESULT(13) => 
                           A_pos_shifted_by1_11_13_port, RESULT(12) => 
                           A_pos_shifted_by1_11_12_port, RESULT(11) => 
                           A_pos_shifted_by1_11_11_port, RESULT(10) => 
                           A_pos_shifted_by1_11_10_port, RESULT(9) => 
                           A_pos_shifted_by1_11_9_port, RESULT(8) => 
                           A_pos_shifted_by1_11_8_port, RESULT(7) => 
                           A_pos_shifted_by1_11_7_port, RESULT(6) => 
                           A_pos_shifted_by1_11_6_port, RESULT(5) => 
                           A_pos_shifted_by1_11_5_port, RESULT(4) => 
                           A_pos_shifted_by1_11_4_port, RESULT(3) => 
                           A_pos_shifted_by1_11_3_port, RESULT(2) => 
                           A_pos_shifted_by1_11_2_port, RESULT(1) => 
                           A_pos_shifted_by1_11_1_port, RESULT(0) => n_1095);
   SHIFTERi_12 : Shifter_NBIT64_20 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_11_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_11_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_11_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_11_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_11_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_11_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_11_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_11_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_11_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_11_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_11_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_11_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_11_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_11_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_11_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_11_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_11_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_11_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_11_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_11_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_11_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_11_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_11_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_11_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_11_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_11_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_11_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_11_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_11_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_11_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_11_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_11_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_11_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_11_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_11_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_11_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_11_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_11_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_11_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_11_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_11_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_11_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_11_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_11_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_11_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_11_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_11_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_11_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_11_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_11_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_11_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_11_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_11_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_11_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_11_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_11_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_11_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_11_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_11_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_11_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_11_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_11_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_11_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_11_0_port, RESULT(127) => 
                           A_pos_shifted_by2_12_63_port, RESULT(126) => 
                           A_pos_shifted_by2_12_62_port, RESULT(125) => 
                           A_pos_shifted_by2_12_61_port, RESULT(124) => 
                           A_pos_shifted_by2_12_60_port, RESULT(123) => 
                           A_pos_shifted_by2_12_59_port, RESULT(122) => 
                           A_pos_shifted_by2_12_58_port, RESULT(121) => 
                           A_pos_shifted_by2_12_57_port, RESULT(120) => 
                           A_pos_shifted_by2_12_56_port, RESULT(119) => 
                           A_pos_shifted_by2_12_55_port, RESULT(118) => 
                           A_pos_shifted_by2_12_54_port, RESULT(117) => 
                           A_pos_shifted_by2_12_53_port, RESULT(116) => 
                           A_pos_shifted_by2_12_52_port, RESULT(115) => 
                           A_pos_shifted_by2_12_51_port, RESULT(114) => 
                           A_pos_shifted_by2_12_50_port, RESULT(113) => 
                           A_pos_shifted_by2_12_49_port, RESULT(112) => 
                           A_pos_shifted_by2_12_48_port, RESULT(111) => 
                           A_pos_shifted_by2_12_47_port, RESULT(110) => 
                           A_pos_shifted_by2_12_46_port, RESULT(109) => 
                           A_pos_shifted_by2_12_45_port, RESULT(108) => 
                           A_pos_shifted_by2_12_44_port, RESULT(107) => 
                           A_pos_shifted_by2_12_43_port, RESULT(106) => 
                           A_pos_shifted_by2_12_42_port, RESULT(105) => 
                           A_pos_shifted_by2_12_41_port, RESULT(104) => 
                           A_pos_shifted_by2_12_40_port, RESULT(103) => 
                           A_pos_shifted_by2_12_39_port, RESULT(102) => 
                           A_pos_shifted_by2_12_38_port, RESULT(101) => 
                           A_pos_shifted_by2_12_37_port, RESULT(100) => 
                           A_pos_shifted_by2_12_36_port, RESULT(99) => 
                           A_pos_shifted_by2_12_35_port, RESULT(98) => 
                           A_pos_shifted_by2_12_34_port, RESULT(97) => 
                           A_pos_shifted_by2_12_33_port, RESULT(96) => 
                           A_pos_shifted_by2_12_32_port, RESULT(95) => 
                           A_pos_shifted_by2_12_31_port, RESULT(94) => 
                           A_pos_shifted_by2_12_30_port, RESULT(93) => 
                           A_pos_shifted_by2_12_29_port, RESULT(92) => 
                           A_pos_shifted_by2_12_28_port, RESULT(91) => 
                           A_pos_shifted_by2_12_27_port, RESULT(90) => 
                           A_pos_shifted_by2_12_26_port, RESULT(89) => 
                           A_pos_shifted_by2_12_25_port, RESULT(88) => 
                           A_pos_shifted_by2_12_24_port, RESULT(87) => 
                           A_pos_shifted_by2_12_23_port, RESULT(86) => 
                           A_pos_shifted_by2_12_22_port, RESULT(85) => 
                           A_pos_shifted_by2_12_21_port, RESULT(84) => 
                           A_pos_shifted_by2_12_20_port, RESULT(83) => 
                           A_pos_shifted_by2_12_19_port, RESULT(82) => 
                           A_pos_shifted_by2_12_18_port, RESULT(81) => 
                           A_pos_shifted_by2_12_17_port, RESULT(80) => 
                           A_pos_shifted_by2_12_16_port, RESULT(79) => 
                           A_pos_shifted_by2_12_15_port, RESULT(78) => 
                           A_pos_shifted_by2_12_14_port, RESULT(77) => 
                           A_pos_shifted_by2_12_13_port, RESULT(76) => 
                           A_pos_shifted_by2_12_12_port, RESULT(75) => 
                           A_pos_shifted_by2_12_11_port, RESULT(74) => 
                           A_pos_shifted_by2_12_10_port, RESULT(73) => 
                           A_pos_shifted_by2_12_9_port, RESULT(72) => 
                           A_pos_shifted_by2_12_8_port, RESULT(71) => 
                           A_pos_shifted_by2_12_7_port, RESULT(70) => 
                           A_pos_shifted_by2_12_6_port, RESULT(69) => 
                           A_pos_shifted_by2_12_5_port, RESULT(68) => 
                           A_pos_shifted_by2_12_4_port, RESULT(67) => 
                           A_pos_shifted_by2_12_3_port, RESULT(66) => 
                           A_pos_shifted_by2_12_2_port, RESULT(65) => n_1096, 
                           RESULT(64) => n_1097, RESULT(63) => 
                           A_pos_shifted_by1_12_63_port, RESULT(62) => 
                           A_pos_shifted_by1_12_62_port, RESULT(61) => 
                           A_pos_shifted_by1_12_61_port, RESULT(60) => 
                           A_pos_shifted_by1_12_60_port, RESULT(59) => 
                           A_pos_shifted_by1_12_59_port, RESULT(58) => 
                           A_pos_shifted_by1_12_58_port, RESULT(57) => 
                           A_pos_shifted_by1_12_57_port, RESULT(56) => 
                           A_pos_shifted_by1_12_56_port, RESULT(55) => 
                           A_pos_shifted_by1_12_55_port, RESULT(54) => 
                           A_pos_shifted_by1_12_54_port, RESULT(53) => 
                           A_pos_shifted_by1_12_53_port, RESULT(52) => 
                           A_pos_shifted_by1_12_52_port, RESULT(51) => 
                           A_pos_shifted_by1_12_51_port, RESULT(50) => 
                           A_pos_shifted_by1_12_50_port, RESULT(49) => 
                           A_pos_shifted_by1_12_49_port, RESULT(48) => 
                           A_pos_shifted_by1_12_48_port, RESULT(47) => 
                           A_pos_shifted_by1_12_47_port, RESULT(46) => 
                           A_pos_shifted_by1_12_46_port, RESULT(45) => 
                           A_pos_shifted_by1_12_45_port, RESULT(44) => 
                           A_pos_shifted_by1_12_44_port, RESULT(43) => 
                           A_pos_shifted_by1_12_43_port, RESULT(42) => 
                           A_pos_shifted_by1_12_42_port, RESULT(41) => 
                           A_pos_shifted_by1_12_41_port, RESULT(40) => 
                           A_pos_shifted_by1_12_40_port, RESULT(39) => 
                           A_pos_shifted_by1_12_39_port, RESULT(38) => 
                           A_pos_shifted_by1_12_38_port, RESULT(37) => 
                           A_pos_shifted_by1_12_37_port, RESULT(36) => 
                           A_pos_shifted_by1_12_36_port, RESULT(35) => 
                           A_pos_shifted_by1_12_35_port, RESULT(34) => 
                           A_pos_shifted_by1_12_34_port, RESULT(33) => 
                           A_pos_shifted_by1_12_33_port, RESULT(32) => 
                           A_pos_shifted_by1_12_32_port, RESULT(31) => 
                           A_pos_shifted_by1_12_31_port, RESULT(30) => 
                           A_pos_shifted_by1_12_30_port, RESULT(29) => 
                           A_pos_shifted_by1_12_29_port, RESULT(28) => 
                           A_pos_shifted_by1_12_28_port, RESULT(27) => 
                           A_pos_shifted_by1_12_27_port, RESULT(26) => 
                           A_pos_shifted_by1_12_26_port, RESULT(25) => 
                           A_pos_shifted_by1_12_25_port, RESULT(24) => 
                           A_pos_shifted_by1_12_24_port, RESULT(23) => 
                           A_pos_shifted_by1_12_23_port, RESULT(22) => 
                           A_pos_shifted_by1_12_22_port, RESULT(21) => 
                           A_pos_shifted_by1_12_21_port, RESULT(20) => 
                           A_pos_shifted_by1_12_20_port, RESULT(19) => 
                           A_pos_shifted_by1_12_19_port, RESULT(18) => 
                           A_pos_shifted_by1_12_18_port, RESULT(17) => 
                           A_pos_shifted_by1_12_17_port, RESULT(16) => 
                           A_pos_shifted_by1_12_16_port, RESULT(15) => 
                           A_pos_shifted_by1_12_15_port, RESULT(14) => 
                           A_pos_shifted_by1_12_14_port, RESULT(13) => 
                           A_pos_shifted_by1_12_13_port, RESULT(12) => 
                           A_pos_shifted_by1_12_12_port, RESULT(11) => 
                           A_pos_shifted_by1_12_11_port, RESULT(10) => 
                           A_pos_shifted_by1_12_10_port, RESULT(9) => 
                           A_pos_shifted_by1_12_9_port, RESULT(8) => 
                           A_pos_shifted_by1_12_8_port, RESULT(7) => 
                           A_pos_shifted_by1_12_7_port, RESULT(6) => 
                           A_pos_shifted_by1_12_6_port, RESULT(5) => 
                           A_pos_shifted_by1_12_5_port, RESULT(4) => 
                           A_pos_shifted_by1_12_4_port, RESULT(3) => 
                           A_pos_shifted_by1_12_3_port, RESULT(2) => 
                           A_pos_shifted_by1_12_2_port, RESULT(1) => 
                           A_pos_shifted_by1_12_1_port, RESULT(0) => n_1098);
   SHIFTERi_13 : Shifter_NBIT64_19 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_12_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_12_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_12_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_12_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_12_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_12_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_12_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_12_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_12_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_12_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_12_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_12_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_12_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_12_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_12_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_12_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_12_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_12_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_12_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_12_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_12_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_12_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_12_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_12_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_12_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_12_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_12_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_12_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_12_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_12_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_12_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_12_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_12_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_12_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_12_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_12_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_12_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_12_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_12_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_12_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_12_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_12_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_12_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_12_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_12_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_12_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_12_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_12_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_12_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_12_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_12_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_12_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_12_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_12_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_12_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_12_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_12_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_12_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_12_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_12_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_12_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_12_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_12_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_12_0_port, RESULT(127) => 
                           A_pos_shifted_by2_13_63_port, RESULT(126) => 
                           A_pos_shifted_by2_13_62_port, RESULT(125) => 
                           A_pos_shifted_by2_13_61_port, RESULT(124) => 
                           A_pos_shifted_by2_13_60_port, RESULT(123) => 
                           A_pos_shifted_by2_13_59_port, RESULT(122) => 
                           A_pos_shifted_by2_13_58_port, RESULT(121) => 
                           A_pos_shifted_by2_13_57_port, RESULT(120) => 
                           A_pos_shifted_by2_13_56_port, RESULT(119) => 
                           A_pos_shifted_by2_13_55_port, RESULT(118) => 
                           A_pos_shifted_by2_13_54_port, RESULT(117) => 
                           A_pos_shifted_by2_13_53_port, RESULT(116) => 
                           A_pos_shifted_by2_13_52_port, RESULT(115) => 
                           A_pos_shifted_by2_13_51_port, RESULT(114) => 
                           A_pos_shifted_by2_13_50_port, RESULT(113) => 
                           A_pos_shifted_by2_13_49_port, RESULT(112) => 
                           A_pos_shifted_by2_13_48_port, RESULT(111) => 
                           A_pos_shifted_by2_13_47_port, RESULT(110) => 
                           A_pos_shifted_by2_13_46_port, RESULT(109) => 
                           A_pos_shifted_by2_13_45_port, RESULT(108) => 
                           A_pos_shifted_by2_13_44_port, RESULT(107) => 
                           A_pos_shifted_by2_13_43_port, RESULT(106) => 
                           A_pos_shifted_by2_13_42_port, RESULT(105) => 
                           A_pos_shifted_by2_13_41_port, RESULT(104) => 
                           A_pos_shifted_by2_13_40_port, RESULT(103) => 
                           A_pos_shifted_by2_13_39_port, RESULT(102) => 
                           A_pos_shifted_by2_13_38_port, RESULT(101) => 
                           A_pos_shifted_by2_13_37_port, RESULT(100) => 
                           A_pos_shifted_by2_13_36_port, RESULT(99) => 
                           A_pos_shifted_by2_13_35_port, RESULT(98) => 
                           A_pos_shifted_by2_13_34_port, RESULT(97) => 
                           A_pos_shifted_by2_13_33_port, RESULT(96) => 
                           A_pos_shifted_by2_13_32_port, RESULT(95) => 
                           A_pos_shifted_by2_13_31_port, RESULT(94) => 
                           A_pos_shifted_by2_13_30_port, RESULT(93) => 
                           A_pos_shifted_by2_13_29_port, RESULT(92) => 
                           A_pos_shifted_by2_13_28_port, RESULT(91) => 
                           A_pos_shifted_by2_13_27_port, RESULT(90) => 
                           A_pos_shifted_by2_13_26_port, RESULT(89) => 
                           A_pos_shifted_by2_13_25_port, RESULT(88) => 
                           A_pos_shifted_by2_13_24_port, RESULT(87) => 
                           A_pos_shifted_by2_13_23_port, RESULT(86) => 
                           A_pos_shifted_by2_13_22_port, RESULT(85) => 
                           A_pos_shifted_by2_13_21_port, RESULT(84) => 
                           A_pos_shifted_by2_13_20_port, RESULT(83) => 
                           A_pos_shifted_by2_13_19_port, RESULT(82) => 
                           A_pos_shifted_by2_13_18_port, RESULT(81) => 
                           A_pos_shifted_by2_13_17_port, RESULT(80) => 
                           A_pos_shifted_by2_13_16_port, RESULT(79) => 
                           A_pos_shifted_by2_13_15_port, RESULT(78) => 
                           A_pos_shifted_by2_13_14_port, RESULT(77) => 
                           A_pos_shifted_by2_13_13_port, RESULT(76) => 
                           A_pos_shifted_by2_13_12_port, RESULT(75) => 
                           A_pos_shifted_by2_13_11_port, RESULT(74) => 
                           A_pos_shifted_by2_13_10_port, RESULT(73) => 
                           A_pos_shifted_by2_13_9_port, RESULT(72) => 
                           A_pos_shifted_by2_13_8_port, RESULT(71) => 
                           A_pos_shifted_by2_13_7_port, RESULT(70) => 
                           A_pos_shifted_by2_13_6_port, RESULT(69) => 
                           A_pos_shifted_by2_13_5_port, RESULT(68) => 
                           A_pos_shifted_by2_13_4_port, RESULT(67) => 
                           A_pos_shifted_by2_13_3_port, RESULT(66) => 
                           A_pos_shifted_by2_13_2_port, RESULT(65) => n_1099, 
                           RESULT(64) => n_1100, RESULT(63) => 
                           A_pos_shifted_by1_13_63_port, RESULT(62) => 
                           A_pos_shifted_by1_13_62_port, RESULT(61) => 
                           A_pos_shifted_by1_13_61_port, RESULT(60) => 
                           A_pos_shifted_by1_13_60_port, RESULT(59) => 
                           A_pos_shifted_by1_13_59_port, RESULT(58) => 
                           A_pos_shifted_by1_13_58_port, RESULT(57) => 
                           A_pos_shifted_by1_13_57_port, RESULT(56) => 
                           A_pos_shifted_by1_13_56_port, RESULT(55) => 
                           A_pos_shifted_by1_13_55_port, RESULT(54) => 
                           A_pos_shifted_by1_13_54_port, RESULT(53) => 
                           A_pos_shifted_by1_13_53_port, RESULT(52) => 
                           A_pos_shifted_by1_13_52_port, RESULT(51) => 
                           A_pos_shifted_by1_13_51_port, RESULT(50) => 
                           A_pos_shifted_by1_13_50_port, RESULT(49) => 
                           A_pos_shifted_by1_13_49_port, RESULT(48) => 
                           A_pos_shifted_by1_13_48_port, RESULT(47) => 
                           A_pos_shifted_by1_13_47_port, RESULT(46) => 
                           A_pos_shifted_by1_13_46_port, RESULT(45) => 
                           A_pos_shifted_by1_13_45_port, RESULT(44) => 
                           A_pos_shifted_by1_13_44_port, RESULT(43) => 
                           A_pos_shifted_by1_13_43_port, RESULT(42) => 
                           A_pos_shifted_by1_13_42_port, RESULT(41) => 
                           A_pos_shifted_by1_13_41_port, RESULT(40) => 
                           A_pos_shifted_by1_13_40_port, RESULT(39) => 
                           A_pos_shifted_by1_13_39_port, RESULT(38) => 
                           A_pos_shifted_by1_13_38_port, RESULT(37) => 
                           A_pos_shifted_by1_13_37_port, RESULT(36) => 
                           A_pos_shifted_by1_13_36_port, RESULT(35) => 
                           A_pos_shifted_by1_13_35_port, RESULT(34) => 
                           A_pos_shifted_by1_13_34_port, RESULT(33) => 
                           A_pos_shifted_by1_13_33_port, RESULT(32) => 
                           A_pos_shifted_by1_13_32_port, RESULT(31) => 
                           A_pos_shifted_by1_13_31_port, RESULT(30) => 
                           A_pos_shifted_by1_13_30_port, RESULT(29) => 
                           A_pos_shifted_by1_13_29_port, RESULT(28) => 
                           A_pos_shifted_by1_13_28_port, RESULT(27) => 
                           A_pos_shifted_by1_13_27_port, RESULT(26) => 
                           A_pos_shifted_by1_13_26_port, RESULT(25) => 
                           A_pos_shifted_by1_13_25_port, RESULT(24) => 
                           A_pos_shifted_by1_13_24_port, RESULT(23) => 
                           A_pos_shifted_by1_13_23_port, RESULT(22) => 
                           A_pos_shifted_by1_13_22_port, RESULT(21) => 
                           A_pos_shifted_by1_13_21_port, RESULT(20) => 
                           A_pos_shifted_by1_13_20_port, RESULT(19) => 
                           A_pos_shifted_by1_13_19_port, RESULT(18) => 
                           A_pos_shifted_by1_13_18_port, RESULT(17) => 
                           A_pos_shifted_by1_13_17_port, RESULT(16) => 
                           A_pos_shifted_by1_13_16_port, RESULT(15) => 
                           A_pos_shifted_by1_13_15_port, RESULT(14) => 
                           A_pos_shifted_by1_13_14_port, RESULT(13) => 
                           A_pos_shifted_by1_13_13_port, RESULT(12) => 
                           A_pos_shifted_by1_13_12_port, RESULT(11) => 
                           A_pos_shifted_by1_13_11_port, RESULT(10) => 
                           A_pos_shifted_by1_13_10_port, RESULT(9) => 
                           A_pos_shifted_by1_13_9_port, RESULT(8) => 
                           A_pos_shifted_by1_13_8_port, RESULT(7) => 
                           A_pos_shifted_by1_13_7_port, RESULT(6) => 
                           A_pos_shifted_by1_13_6_port, RESULT(5) => 
                           A_pos_shifted_by1_13_5_port, RESULT(4) => 
                           A_pos_shifted_by1_13_4_port, RESULT(3) => 
                           A_pos_shifted_by1_13_3_port, RESULT(2) => 
                           A_pos_shifted_by1_13_2_port, RESULT(1) => 
                           A_pos_shifted_by1_13_1_port, RESULT(0) => n_1101);
   SHIFTERi_14 : Shifter_NBIT64_18 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_13_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_13_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_13_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_13_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_13_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_13_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_13_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_13_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_13_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_13_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_13_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_13_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_13_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_13_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_13_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_13_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_13_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_13_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_13_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_13_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_13_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_13_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_13_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_13_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_13_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_13_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_13_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_13_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_13_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_13_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_13_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_13_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_13_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_13_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_13_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_13_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_13_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_13_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_13_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_13_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_13_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_13_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_13_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_13_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_13_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_13_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_13_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_13_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_13_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_13_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_13_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_13_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_13_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_13_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_13_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_13_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_13_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_13_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_13_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_13_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_13_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_13_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_13_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_13_0_port, RESULT(127) => 
                           A_pos_shifted_by2_14_63_port, RESULT(126) => 
                           A_pos_shifted_by2_14_62_port, RESULT(125) => 
                           A_pos_shifted_by2_14_61_port, RESULT(124) => 
                           A_pos_shifted_by2_14_60_port, RESULT(123) => 
                           A_pos_shifted_by2_14_59_port, RESULT(122) => 
                           A_pos_shifted_by2_14_58_port, RESULT(121) => 
                           A_pos_shifted_by2_14_57_port, RESULT(120) => 
                           A_pos_shifted_by2_14_56_port, RESULT(119) => 
                           A_pos_shifted_by2_14_55_port, RESULT(118) => 
                           A_pos_shifted_by2_14_54_port, RESULT(117) => 
                           A_pos_shifted_by2_14_53_port, RESULT(116) => 
                           A_pos_shifted_by2_14_52_port, RESULT(115) => 
                           A_pos_shifted_by2_14_51_port, RESULT(114) => 
                           A_pos_shifted_by2_14_50_port, RESULT(113) => 
                           A_pos_shifted_by2_14_49_port, RESULT(112) => 
                           A_pos_shifted_by2_14_48_port, RESULT(111) => 
                           A_pos_shifted_by2_14_47_port, RESULT(110) => 
                           A_pos_shifted_by2_14_46_port, RESULT(109) => 
                           A_pos_shifted_by2_14_45_port, RESULT(108) => 
                           A_pos_shifted_by2_14_44_port, RESULT(107) => 
                           A_pos_shifted_by2_14_43_port, RESULT(106) => 
                           A_pos_shifted_by2_14_42_port, RESULT(105) => 
                           A_pos_shifted_by2_14_41_port, RESULT(104) => 
                           A_pos_shifted_by2_14_40_port, RESULT(103) => 
                           A_pos_shifted_by2_14_39_port, RESULT(102) => 
                           A_pos_shifted_by2_14_38_port, RESULT(101) => 
                           A_pos_shifted_by2_14_37_port, RESULT(100) => 
                           A_pos_shifted_by2_14_36_port, RESULT(99) => 
                           A_pos_shifted_by2_14_35_port, RESULT(98) => 
                           A_pos_shifted_by2_14_34_port, RESULT(97) => 
                           A_pos_shifted_by2_14_33_port, RESULT(96) => 
                           A_pos_shifted_by2_14_32_port, RESULT(95) => 
                           A_pos_shifted_by2_14_31_port, RESULT(94) => 
                           A_pos_shifted_by2_14_30_port, RESULT(93) => 
                           A_pos_shifted_by2_14_29_port, RESULT(92) => 
                           A_pos_shifted_by2_14_28_port, RESULT(91) => 
                           A_pos_shifted_by2_14_27_port, RESULT(90) => 
                           A_pos_shifted_by2_14_26_port, RESULT(89) => 
                           A_pos_shifted_by2_14_25_port, RESULT(88) => 
                           A_pos_shifted_by2_14_24_port, RESULT(87) => 
                           A_pos_shifted_by2_14_23_port, RESULT(86) => 
                           A_pos_shifted_by2_14_22_port, RESULT(85) => 
                           A_pos_shifted_by2_14_21_port, RESULT(84) => 
                           A_pos_shifted_by2_14_20_port, RESULT(83) => 
                           A_pos_shifted_by2_14_19_port, RESULT(82) => 
                           A_pos_shifted_by2_14_18_port, RESULT(81) => 
                           A_pos_shifted_by2_14_17_port, RESULT(80) => 
                           A_pos_shifted_by2_14_16_port, RESULT(79) => 
                           A_pos_shifted_by2_14_15_port, RESULT(78) => 
                           A_pos_shifted_by2_14_14_port, RESULT(77) => 
                           A_pos_shifted_by2_14_13_port, RESULT(76) => 
                           A_pos_shifted_by2_14_12_port, RESULT(75) => 
                           A_pos_shifted_by2_14_11_port, RESULT(74) => 
                           A_pos_shifted_by2_14_10_port, RESULT(73) => 
                           A_pos_shifted_by2_14_9_port, RESULT(72) => 
                           A_pos_shifted_by2_14_8_port, RESULT(71) => 
                           A_pos_shifted_by2_14_7_port, RESULT(70) => 
                           A_pos_shifted_by2_14_6_port, RESULT(69) => 
                           A_pos_shifted_by2_14_5_port, RESULT(68) => 
                           A_pos_shifted_by2_14_4_port, RESULT(67) => 
                           A_pos_shifted_by2_14_3_port, RESULT(66) => 
                           A_pos_shifted_by2_14_2_port, RESULT(65) => n_1102, 
                           RESULT(64) => n_1103, RESULT(63) => 
                           A_pos_shifted_by1_14_63_port, RESULT(62) => 
                           A_pos_shifted_by1_14_62_port, RESULT(61) => 
                           A_pos_shifted_by1_14_61_port, RESULT(60) => 
                           A_pos_shifted_by1_14_60_port, RESULT(59) => 
                           A_pos_shifted_by1_14_59_port, RESULT(58) => 
                           A_pos_shifted_by1_14_58_port, RESULT(57) => 
                           A_pos_shifted_by1_14_57_port, RESULT(56) => 
                           A_pos_shifted_by1_14_56_port, RESULT(55) => 
                           A_pos_shifted_by1_14_55_port, RESULT(54) => 
                           A_pos_shifted_by1_14_54_port, RESULT(53) => 
                           A_pos_shifted_by1_14_53_port, RESULT(52) => 
                           A_pos_shifted_by1_14_52_port, RESULT(51) => 
                           A_pos_shifted_by1_14_51_port, RESULT(50) => 
                           A_pos_shifted_by1_14_50_port, RESULT(49) => 
                           A_pos_shifted_by1_14_49_port, RESULT(48) => 
                           A_pos_shifted_by1_14_48_port, RESULT(47) => 
                           A_pos_shifted_by1_14_47_port, RESULT(46) => 
                           A_pos_shifted_by1_14_46_port, RESULT(45) => 
                           A_pos_shifted_by1_14_45_port, RESULT(44) => 
                           A_pos_shifted_by1_14_44_port, RESULT(43) => 
                           A_pos_shifted_by1_14_43_port, RESULT(42) => 
                           A_pos_shifted_by1_14_42_port, RESULT(41) => 
                           A_pos_shifted_by1_14_41_port, RESULT(40) => 
                           A_pos_shifted_by1_14_40_port, RESULT(39) => 
                           A_pos_shifted_by1_14_39_port, RESULT(38) => 
                           A_pos_shifted_by1_14_38_port, RESULT(37) => 
                           A_pos_shifted_by1_14_37_port, RESULT(36) => 
                           A_pos_shifted_by1_14_36_port, RESULT(35) => 
                           A_pos_shifted_by1_14_35_port, RESULT(34) => 
                           A_pos_shifted_by1_14_34_port, RESULT(33) => 
                           A_pos_shifted_by1_14_33_port, RESULT(32) => 
                           A_pos_shifted_by1_14_32_port, RESULT(31) => 
                           A_pos_shifted_by1_14_31_port, RESULT(30) => 
                           A_pos_shifted_by1_14_30_port, RESULT(29) => 
                           A_pos_shifted_by1_14_29_port, RESULT(28) => 
                           A_pos_shifted_by1_14_28_port, RESULT(27) => 
                           A_pos_shifted_by1_14_27_port, RESULT(26) => 
                           A_pos_shifted_by1_14_26_port, RESULT(25) => 
                           A_pos_shifted_by1_14_25_port, RESULT(24) => 
                           A_pos_shifted_by1_14_24_port, RESULT(23) => 
                           A_pos_shifted_by1_14_23_port, RESULT(22) => 
                           A_pos_shifted_by1_14_22_port, RESULT(21) => 
                           A_pos_shifted_by1_14_21_port, RESULT(20) => 
                           A_pos_shifted_by1_14_20_port, RESULT(19) => 
                           A_pos_shifted_by1_14_19_port, RESULT(18) => 
                           A_pos_shifted_by1_14_18_port, RESULT(17) => 
                           A_pos_shifted_by1_14_17_port, RESULT(16) => 
                           A_pos_shifted_by1_14_16_port, RESULT(15) => 
                           A_pos_shifted_by1_14_15_port, RESULT(14) => 
                           A_pos_shifted_by1_14_14_port, RESULT(13) => 
                           A_pos_shifted_by1_14_13_port, RESULT(12) => 
                           A_pos_shifted_by1_14_12_port, RESULT(11) => 
                           A_pos_shifted_by1_14_11_port, RESULT(10) => 
                           A_pos_shifted_by1_14_10_port, RESULT(9) => 
                           A_pos_shifted_by1_14_9_port, RESULT(8) => 
                           A_pos_shifted_by1_14_8_port, RESULT(7) => 
                           A_pos_shifted_by1_14_7_port, RESULT(6) => 
                           A_pos_shifted_by1_14_6_port, RESULT(5) => 
                           A_pos_shifted_by1_14_5_port, RESULT(4) => 
                           A_pos_shifted_by1_14_4_port, RESULT(3) => 
                           A_pos_shifted_by1_14_3_port, RESULT(2) => 
                           A_pos_shifted_by1_14_2_port, RESULT(1) => 
                           A_pos_shifted_by1_14_1_port, RESULT(0) => n_1104);
   SHIFTERi_15 : Shifter_NBIT64_17 port map( TO_SHIFT(63) => 
                           A_pos_shifted_by2_14_63_port, TO_SHIFT(62) => 
                           A_pos_shifted_by2_14_62_port, TO_SHIFT(61) => 
                           A_pos_shifted_by2_14_61_port, TO_SHIFT(60) => 
                           A_pos_shifted_by2_14_60_port, TO_SHIFT(59) => 
                           A_pos_shifted_by2_14_59_port, TO_SHIFT(58) => 
                           A_pos_shifted_by2_14_58_port, TO_SHIFT(57) => 
                           A_pos_shifted_by2_14_57_port, TO_SHIFT(56) => 
                           A_pos_shifted_by2_14_56_port, TO_SHIFT(55) => 
                           A_pos_shifted_by2_14_55_port, TO_SHIFT(54) => 
                           A_pos_shifted_by2_14_54_port, TO_SHIFT(53) => 
                           A_pos_shifted_by2_14_53_port, TO_SHIFT(52) => 
                           A_pos_shifted_by2_14_52_port, TO_SHIFT(51) => 
                           A_pos_shifted_by2_14_51_port, TO_SHIFT(50) => 
                           A_pos_shifted_by2_14_50_port, TO_SHIFT(49) => 
                           A_pos_shifted_by2_14_49_port, TO_SHIFT(48) => 
                           A_pos_shifted_by2_14_48_port, TO_SHIFT(47) => 
                           A_pos_shifted_by2_14_47_port, TO_SHIFT(46) => 
                           A_pos_shifted_by2_14_46_port, TO_SHIFT(45) => 
                           A_pos_shifted_by2_14_45_port, TO_SHIFT(44) => 
                           A_pos_shifted_by2_14_44_port, TO_SHIFT(43) => 
                           A_pos_shifted_by2_14_43_port, TO_SHIFT(42) => 
                           A_pos_shifted_by2_14_42_port, TO_SHIFT(41) => 
                           A_pos_shifted_by2_14_41_port, TO_SHIFT(40) => 
                           A_pos_shifted_by2_14_40_port, TO_SHIFT(39) => 
                           A_pos_shifted_by2_14_39_port, TO_SHIFT(38) => 
                           A_pos_shifted_by2_14_38_port, TO_SHIFT(37) => 
                           A_pos_shifted_by2_14_37_port, TO_SHIFT(36) => 
                           A_pos_shifted_by2_14_36_port, TO_SHIFT(35) => 
                           A_pos_shifted_by2_14_35_port, TO_SHIFT(34) => 
                           A_pos_shifted_by2_14_34_port, TO_SHIFT(33) => 
                           A_pos_shifted_by2_14_33_port, TO_SHIFT(32) => 
                           A_pos_shifted_by2_14_32_port, TO_SHIFT(31) => 
                           A_pos_shifted_by2_14_31_port, TO_SHIFT(30) => 
                           A_pos_shifted_by2_14_30_port, TO_SHIFT(29) => 
                           A_pos_shifted_by2_14_29_port, TO_SHIFT(28) => 
                           A_pos_shifted_by2_14_28_port, TO_SHIFT(27) => 
                           A_pos_shifted_by2_14_27_port, TO_SHIFT(26) => 
                           A_pos_shifted_by2_14_26_port, TO_SHIFT(25) => 
                           A_pos_shifted_by2_14_25_port, TO_SHIFT(24) => 
                           A_pos_shifted_by2_14_24_port, TO_SHIFT(23) => 
                           A_pos_shifted_by2_14_23_port, TO_SHIFT(22) => 
                           A_pos_shifted_by2_14_22_port, TO_SHIFT(21) => 
                           A_pos_shifted_by2_14_21_port, TO_SHIFT(20) => 
                           A_pos_shifted_by2_14_20_port, TO_SHIFT(19) => 
                           A_pos_shifted_by2_14_19_port, TO_SHIFT(18) => 
                           A_pos_shifted_by2_14_18_port, TO_SHIFT(17) => 
                           A_pos_shifted_by2_14_17_port, TO_SHIFT(16) => 
                           A_pos_shifted_by2_14_16_port, TO_SHIFT(15) => 
                           A_pos_shifted_by2_14_15_port, TO_SHIFT(14) => 
                           A_pos_shifted_by2_14_14_port, TO_SHIFT(13) => 
                           A_pos_shifted_by2_14_13_port, TO_SHIFT(12) => 
                           A_pos_shifted_by2_14_12_port, TO_SHIFT(11) => 
                           A_pos_shifted_by2_14_11_port, TO_SHIFT(10) => 
                           A_pos_shifted_by2_14_10_port, TO_SHIFT(9) => 
                           A_pos_shifted_by2_14_9_port, TO_SHIFT(8) => 
                           A_pos_shifted_by2_14_8_port, TO_SHIFT(7) => 
                           A_pos_shifted_by2_14_7_port, TO_SHIFT(6) => 
                           A_pos_shifted_by2_14_6_port, TO_SHIFT(5) => 
                           A_pos_shifted_by2_14_5_port, TO_SHIFT(4) => 
                           A_pos_shifted_by2_14_4_port, TO_SHIFT(3) => 
                           A_pos_shifted_by2_14_3_port, TO_SHIFT(2) => 
                           A_pos_shifted_by2_14_2_port, TO_SHIFT(1) => 
                           A_pos_shifted_by2_14_1_port, TO_SHIFT(0) => 
                           A_pos_shifted_by2_14_0_port, RESULT(127) => n_1105, 
                           RESULT(126) => n_1106, RESULT(125) => n_1107, 
                           RESULT(124) => n_1108, RESULT(123) => n_1109, 
                           RESULT(122) => n_1110, RESULT(121) => n_1111, 
                           RESULT(120) => n_1112, RESULT(119) => n_1113, 
                           RESULT(118) => n_1114, RESULT(117) => n_1115, 
                           RESULT(116) => n_1116, RESULT(115) => n_1117, 
                           RESULT(114) => n_1118, RESULT(113) => n_1119, 
                           RESULT(112) => n_1120, RESULT(111) => n_1121, 
                           RESULT(110) => n_1122, RESULT(109) => n_1123, 
                           RESULT(108) => n_1124, RESULT(107) => n_1125, 
                           RESULT(106) => n_1126, RESULT(105) => n_1127, 
                           RESULT(104) => n_1128, RESULT(103) => n_1129, 
                           RESULT(102) => n_1130, RESULT(101) => n_1131, 
                           RESULT(100) => n_1132, RESULT(99) => n_1133, 
                           RESULT(98) => n_1134, RESULT(97) => n_1135, 
                           RESULT(96) => n_1136, RESULT(95) => n_1137, 
                           RESULT(94) => n_1138, RESULT(93) => n_1139, 
                           RESULT(92) => n_1140, RESULT(91) => n_1141, 
                           RESULT(90) => n_1142, RESULT(89) => n_1143, 
                           RESULT(88) => n_1144, RESULT(87) => n_1145, 
                           RESULT(86) => n_1146, RESULT(85) => n_1147, 
                           RESULT(84) => n_1148, RESULT(83) => n_1149, 
                           RESULT(82) => n_1150, RESULT(81) => n_1151, 
                           RESULT(80) => n_1152, RESULT(79) => n_1153, 
                           RESULT(78) => n_1154, RESULT(77) => n_1155, 
                           RESULT(76) => n_1156, RESULT(75) => n_1157, 
                           RESULT(74) => n_1158, RESULT(73) => n_1159, 
                           RESULT(72) => n_1160, RESULT(71) => n_1161, 
                           RESULT(70) => n_1162, RESULT(69) => n_1163, 
                           RESULT(68) => n_1164, RESULT(67) => n_1165, 
                           RESULT(66) => n_1166, RESULT(65) => n_1167, 
                           RESULT(64) => n_1168, RESULT(63) => 
                           A_pos_shifted_by1_15_63_port, RESULT(62) => 
                           A_pos_shifted_by1_15_62_port, RESULT(61) => 
                           A_pos_shifted_by1_15_61_port, RESULT(60) => 
                           A_pos_shifted_by1_15_60_port, RESULT(59) => 
                           A_pos_shifted_by1_15_59_port, RESULT(58) => 
                           A_pos_shifted_by1_15_58_port, RESULT(57) => 
                           A_pos_shifted_by1_15_57_port, RESULT(56) => 
                           A_pos_shifted_by1_15_56_port, RESULT(55) => 
                           A_pos_shifted_by1_15_55_port, RESULT(54) => 
                           A_pos_shifted_by1_15_54_port, RESULT(53) => 
                           A_pos_shifted_by1_15_53_port, RESULT(52) => 
                           A_pos_shifted_by1_15_52_port, RESULT(51) => 
                           A_pos_shifted_by1_15_51_port, RESULT(50) => 
                           A_pos_shifted_by1_15_50_port, RESULT(49) => 
                           A_pos_shifted_by1_15_49_port, RESULT(48) => 
                           A_pos_shifted_by1_15_48_port, RESULT(47) => 
                           A_pos_shifted_by1_15_47_port, RESULT(46) => 
                           A_pos_shifted_by1_15_46_port, RESULT(45) => 
                           A_pos_shifted_by1_15_45_port, RESULT(44) => 
                           A_pos_shifted_by1_15_44_port, RESULT(43) => 
                           A_pos_shifted_by1_15_43_port, RESULT(42) => 
                           A_pos_shifted_by1_15_42_port, RESULT(41) => 
                           A_pos_shifted_by1_15_41_port, RESULT(40) => 
                           A_pos_shifted_by1_15_40_port, RESULT(39) => 
                           A_pos_shifted_by1_15_39_port, RESULT(38) => 
                           A_pos_shifted_by1_15_38_port, RESULT(37) => 
                           A_pos_shifted_by1_15_37_port, RESULT(36) => 
                           A_pos_shifted_by1_15_36_port, RESULT(35) => 
                           A_pos_shifted_by1_15_35_port, RESULT(34) => 
                           A_pos_shifted_by1_15_34_port, RESULT(33) => 
                           A_pos_shifted_by1_15_33_port, RESULT(32) => 
                           A_pos_shifted_by1_15_32_port, RESULT(31) => 
                           A_pos_shifted_by1_15_31_port, RESULT(30) => 
                           A_pos_shifted_by1_15_30_port, RESULT(29) => 
                           A_pos_shifted_by1_15_29_port, RESULT(28) => 
                           A_pos_shifted_by1_15_28_port, RESULT(27) => 
                           A_pos_shifted_by1_15_27_port, RESULT(26) => 
                           A_pos_shifted_by1_15_26_port, RESULT(25) => 
                           A_pos_shifted_by1_15_25_port, RESULT(24) => 
                           A_pos_shifted_by1_15_24_port, RESULT(23) => 
                           A_pos_shifted_by1_15_23_port, RESULT(22) => 
                           A_pos_shifted_by1_15_22_port, RESULT(21) => 
                           A_pos_shifted_by1_15_21_port, RESULT(20) => 
                           A_pos_shifted_by1_15_20_port, RESULT(19) => 
                           A_pos_shifted_by1_15_19_port, RESULT(18) => 
                           A_pos_shifted_by1_15_18_port, RESULT(17) => 
                           A_pos_shifted_by1_15_17_port, RESULT(16) => 
                           A_pos_shifted_by1_15_16_port, RESULT(15) => 
                           A_pos_shifted_by1_15_15_port, RESULT(14) => 
                           A_pos_shifted_by1_15_14_port, RESULT(13) => 
                           A_pos_shifted_by1_15_13_port, RESULT(12) => 
                           A_pos_shifted_by1_15_12_port, RESULT(11) => 
                           A_pos_shifted_by1_15_11_port, RESULT(10) => 
                           A_pos_shifted_by1_15_10_port, RESULT(9) => 
                           A_pos_shifted_by1_15_9_port, RESULT(8) => 
                           A_pos_shifted_by1_15_8_port, RESULT(7) => 
                           A_pos_shifted_by1_15_7_port, RESULT(6) => 
                           A_pos_shifted_by1_15_6_port, RESULT(5) => 
                           A_pos_shifted_by1_15_5_port, RESULT(4) => 
                           A_pos_shifted_by1_15_4_port, RESULT(3) => 
                           A_pos_shifted_by1_15_3_port, RESULT(2) => 
                           A_pos_shifted_by1_15_2_port, RESULT(1) => 
                           A_pos_shifted_by1_15_1_port, RESULT(0) => n_1169);
   SHIFTER0_0_0 : Shifter_NBIT64_16 port map( TO_SHIFT(63) => n196, 
                           TO_SHIFT(62) => n200, TO_SHIFT(61) => n200, 
                           TO_SHIFT(60) => n200, TO_SHIFT(59) => n200, 
                           TO_SHIFT(58) => n199, TO_SHIFT(57) => n199, 
                           TO_SHIFT(56) => n198, TO_SHIFT(55) => n199, 
                           TO_SHIFT(54) => n198, TO_SHIFT(53) => n198, 
                           TO_SHIFT(52) => n198, TO_SHIFT(51) => n197, 
                           TO_SHIFT(50) => n199, TO_SHIFT(49) => n199, 
                           TO_SHIFT(48) => n196, TO_SHIFT(47) => n196, 
                           TO_SHIFT(46) => n200, TO_SHIFT(45) => n200, 
                           TO_SHIFT(44) => n200, TO_SHIFT(43) => n200, 
                           TO_SHIFT(42) => n199, TO_SHIFT(41) => n199, 
                           TO_SHIFT(40) => n199, TO_SHIFT(39) => n199, 
                           TO_SHIFT(38) => n199, TO_SHIFT(37) => n198, 
                           TO_SHIFT(36) => n197, TO_SHIFT(35) => n197, 
                           TO_SHIFT(34) => n197, TO_SHIFT(33) => n201, 
                           TO_SHIFT(32) => n196, TO_SHIFT(31) => 
                           A_neg_tmp_31_port, TO_SHIFT(30) => A_neg_tmp_30_port
                           , TO_SHIFT(29) => A_neg_tmp_29_port, TO_SHIFT(28) =>
                           A_neg_tmp_28_port, TO_SHIFT(27) => A_neg_tmp_27_port
                           , TO_SHIFT(26) => A_neg_tmp_26_port, TO_SHIFT(25) =>
                           A_neg_tmp_25_port, TO_SHIFT(24) => A_neg_tmp_24_port
                           , TO_SHIFT(23) => A_neg_tmp_23_port, TO_SHIFT(22) =>
                           A_neg_tmp_22_port, TO_SHIFT(21) => A_neg_tmp_21_port
                           , TO_SHIFT(20) => A_neg_tmp_20_port, TO_SHIFT(19) =>
                           A_neg_tmp_19_port, TO_SHIFT(18) => A_neg_tmp_18_port
                           , TO_SHIFT(17) => A_neg_tmp_17_port, TO_SHIFT(16) =>
                           A_neg_tmp_16_port, TO_SHIFT(15) => A_neg_tmp_15_port
                           , TO_SHIFT(14) => A_neg_tmp_14_port, TO_SHIFT(13) =>
                           A_neg_tmp_13_port, TO_SHIFT(12) => A_neg_tmp_12_port
                           , TO_SHIFT(11) => A_neg_tmp_11_port, TO_SHIFT(10) =>
                           A_neg_tmp_10_port, TO_SHIFT(9) => n182, TO_SHIFT(8) 
                           => A_neg_tmp_8_port, TO_SHIFT(7) => n177, 
                           TO_SHIFT(6) => n185, TO_SHIFT(5) => n186, 
                           TO_SHIFT(4) => n194, TO_SHIFT(3) => n188, 
                           TO_SHIFT(2) => n178, TO_SHIFT(1) => A_neg_tmp_1_port
                           , TO_SHIFT(0) => A_neg_tmp_0_port, RESULT(127) => 
                           A_neg_shifted_by2_0_63_port, RESULT(126) => 
                           A_neg_shifted_by2_0_62_port, RESULT(125) => 
                           A_neg_shifted_by2_0_61_port, RESULT(124) => 
                           A_neg_shifted_by2_0_60_port, RESULT(123) => 
                           A_neg_shifted_by2_0_59_port, RESULT(122) => 
                           A_neg_shifted_by2_0_58_port, RESULT(121) => 
                           A_neg_shifted_by2_0_57_port, RESULT(120) => 
                           A_neg_shifted_by2_0_56_port, RESULT(119) => 
                           A_neg_shifted_by2_0_55_port, RESULT(118) => 
                           A_neg_shifted_by2_0_54_port, RESULT(117) => 
                           A_neg_shifted_by2_0_53_port, RESULT(116) => 
                           A_neg_shifted_by2_0_52_port, RESULT(115) => 
                           A_neg_shifted_by2_0_51_port, RESULT(114) => 
                           A_neg_shifted_by2_0_50_port, RESULT(113) => 
                           A_neg_shifted_by2_0_49_port, RESULT(112) => 
                           A_neg_shifted_by2_0_48_port, RESULT(111) => 
                           A_neg_shifted_by2_0_47_port, RESULT(110) => 
                           A_neg_shifted_by2_0_46_port, RESULT(109) => 
                           A_neg_shifted_by2_0_45_port, RESULT(108) => 
                           A_neg_shifted_by2_0_44_port, RESULT(107) => 
                           A_neg_shifted_by2_0_43_port, RESULT(106) => 
                           A_neg_shifted_by2_0_42_port, RESULT(105) => 
                           A_neg_shifted_by2_0_41_port, RESULT(104) => 
                           A_neg_shifted_by2_0_40_port, RESULT(103) => 
                           A_neg_shifted_by2_0_39_port, RESULT(102) => 
                           A_neg_shifted_by2_0_38_port, RESULT(101) => 
                           A_neg_shifted_by2_0_37_port, RESULT(100) => 
                           A_neg_shifted_by2_0_36_port, RESULT(99) => 
                           A_neg_shifted_by2_0_35_port, RESULT(98) => 
                           A_neg_shifted_by2_0_34_port, RESULT(97) => 
                           A_neg_shifted_by2_0_33_port, RESULT(96) => 
                           A_neg_shifted_by2_0_32_port, RESULT(95) => 
                           A_neg_shifted_by2_0_31_port, RESULT(94) => 
                           A_neg_shifted_by2_0_30_port, RESULT(93) => 
                           A_neg_shifted_by2_0_29_port, RESULT(92) => 
                           A_neg_shifted_by2_0_28_port, RESULT(91) => 
                           A_neg_shifted_by2_0_27_port, RESULT(90) => 
                           A_neg_shifted_by2_0_26_port, RESULT(89) => 
                           A_neg_shifted_by2_0_25_port, RESULT(88) => 
                           A_neg_shifted_by2_0_24_port, RESULT(87) => 
                           A_neg_shifted_by2_0_23_port, RESULT(86) => 
                           A_neg_shifted_by2_0_22_port, RESULT(85) => 
                           A_neg_shifted_by2_0_21_port, RESULT(84) => 
                           A_neg_shifted_by2_0_20_port, RESULT(83) => 
                           A_neg_shifted_by2_0_19_port, RESULT(82) => 
                           A_neg_shifted_by2_0_18_port, RESULT(81) => 
                           A_neg_shifted_by2_0_17_port, RESULT(80) => 
                           A_neg_shifted_by2_0_16_port, RESULT(79) => 
                           A_neg_shifted_by2_0_15_port, RESULT(78) => 
                           A_neg_shifted_by2_0_14_port, RESULT(77) => 
                           A_neg_shifted_by2_0_13_port, RESULT(76) => 
                           A_neg_shifted_by2_0_12_port, RESULT(75) => 
                           A_neg_shifted_by2_0_11_port, RESULT(74) => 
                           A_neg_shifted_by2_0_10_port, RESULT(73) => 
                           A_neg_shifted_by2_0_9_port, RESULT(72) => 
                           A_neg_shifted_by2_0_8_port, RESULT(71) => 
                           A_neg_shifted_by2_0_7_port, RESULT(70) => 
                           A_neg_shifted_by2_0_6_port, RESULT(69) => 
                           A_neg_shifted_by2_0_5_port, RESULT(68) => 
                           A_neg_shifted_by2_0_4_port, RESULT(67) => 
                           A_neg_shifted_by2_0_3_port, RESULT(66) => 
                           A_neg_shifted_by2_0_2_port, RESULT(65) => n_1170, 
                           RESULT(64) => n_1171, RESULT(63) => 
                           A_neg_shifted_by1_0_63_port, RESULT(62) => 
                           A_neg_shifted_by1_0_62_port, RESULT(61) => 
                           A_neg_shifted_by1_0_61_port, RESULT(60) => 
                           A_neg_shifted_by1_0_60_port, RESULT(59) => 
                           A_neg_shifted_by1_0_59_port, RESULT(58) => 
                           A_neg_shifted_by1_0_58_port, RESULT(57) => 
                           A_neg_shifted_by1_0_57_port, RESULT(56) => 
                           A_neg_shifted_by1_0_56_port, RESULT(55) => 
                           A_neg_shifted_by1_0_55_port, RESULT(54) => 
                           A_neg_shifted_by1_0_54_port, RESULT(53) => 
                           A_neg_shifted_by1_0_53_port, RESULT(52) => 
                           A_neg_shifted_by1_0_52_port, RESULT(51) => 
                           A_neg_shifted_by1_0_51_port, RESULT(50) => 
                           A_neg_shifted_by1_0_50_port, RESULT(49) => 
                           A_neg_shifted_by1_0_49_port, RESULT(48) => 
                           A_neg_shifted_by1_0_48_port, RESULT(47) => 
                           A_neg_shifted_by1_0_47_port, RESULT(46) => 
                           A_neg_shifted_by1_0_46_port, RESULT(45) => 
                           A_neg_shifted_by1_0_45_port, RESULT(44) => 
                           A_neg_shifted_by1_0_44_port, RESULT(43) => 
                           A_neg_shifted_by1_0_43_port, RESULT(42) => 
                           A_neg_shifted_by1_0_42_port, RESULT(41) => 
                           A_neg_shifted_by1_0_41_port, RESULT(40) => 
                           A_neg_shifted_by1_0_40_port, RESULT(39) => 
                           A_neg_shifted_by1_0_39_port, RESULT(38) => 
                           A_neg_shifted_by1_0_38_port, RESULT(37) => 
                           A_neg_shifted_by1_0_37_port, RESULT(36) => 
                           A_neg_shifted_by1_0_36_port, RESULT(35) => 
                           A_neg_shifted_by1_0_35_port, RESULT(34) => 
                           A_neg_shifted_by1_0_34_port, RESULT(33) => 
                           A_neg_shifted_by1_0_33_port, RESULT(32) => 
                           A_neg_shifted_by1_0_32_port, RESULT(31) => 
                           A_neg_shifted_by1_0_31_port, RESULT(30) => 
                           A_neg_shifted_by1_0_30_port, RESULT(29) => 
                           A_neg_shifted_by1_0_29_port, RESULT(28) => 
                           A_neg_shifted_by1_0_28_port, RESULT(27) => 
                           A_neg_shifted_by1_0_27_port, RESULT(26) => 
                           A_neg_shifted_by1_0_26_port, RESULT(25) => 
                           A_neg_shifted_by1_0_25_port, RESULT(24) => 
                           A_neg_shifted_by1_0_24_port, RESULT(23) => 
                           A_neg_shifted_by1_0_23_port, RESULT(22) => 
                           A_neg_shifted_by1_0_22_port, RESULT(21) => 
                           A_neg_shifted_by1_0_21_port, RESULT(20) => 
                           A_neg_shifted_by1_0_20_port, RESULT(19) => 
                           A_neg_shifted_by1_0_19_port, RESULT(18) => 
                           A_neg_shifted_by1_0_18_port, RESULT(17) => 
                           A_neg_shifted_by1_0_17_port, RESULT(16) => 
                           A_neg_shifted_by1_0_16_port, RESULT(15) => 
                           A_neg_shifted_by1_0_15_port, RESULT(14) => 
                           A_neg_shifted_by1_0_14_port, RESULT(13) => 
                           A_neg_shifted_by1_0_13_port, RESULT(12) => 
                           A_neg_shifted_by1_0_12_port, RESULT(11) => 
                           A_neg_shifted_by1_0_11_port, RESULT(10) => 
                           A_neg_shifted_by1_0_10_port, RESULT(9) => 
                           A_neg_shifted_by1_0_9_port, RESULT(8) => 
                           A_neg_shifted_by1_0_8_port, RESULT(7) => 
                           A_neg_shifted_by1_0_7_port, RESULT(6) => 
                           A_neg_shifted_by1_0_6_port, RESULT(5) => 
                           A_neg_shifted_by1_0_5_port, RESULT(4) => 
                           A_neg_shifted_by1_0_4_port, RESULT(3) => 
                           A_neg_shifted_by1_0_3_port, RESULT(2) => 
                           A_neg_shifted_by1_0_2_port, RESULT(1) => 
                           A_neg_shifted_by1_0_1_port, RESULT(0) => n_1172);
   SHIFTERi_1_0 : Shifter_NBIT64_15 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_0_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_0_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_0_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_0_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_0_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_0_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_0_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_0_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_0_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_0_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_0_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_0_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_0_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_0_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_0_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_0_48_port, TO_SHIFT(47) => n207, 
                           TO_SHIFT(46) => A_neg_shifted_by2_0_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_0_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_0_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_0_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_0_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_0_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_0_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_0_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_0_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_0_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_0_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_0_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_0_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_0_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_0_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_0_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_0_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_0_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_0_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_0_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_0_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_0_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_0_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_0_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_0_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_0_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_0_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_0_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_0_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_0_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_0_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_0_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_0_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_0_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_0_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_0_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_0_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_0_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_0_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_0_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_0_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_0_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_0_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_0_3_port, 
                           TO_SHIFT(2) => n187, TO_SHIFT(1) => 
                           A_neg_shifted_by2_0_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_0_0_port, RESULT(127) => 
                           A_neg_shifted_by2_1_63_port, RESULT(126) => 
                           A_neg_shifted_by2_1_62_port, RESULT(125) => 
                           A_neg_shifted_by2_1_61_port, RESULT(124) => 
                           A_neg_shifted_by2_1_60_port, RESULT(123) => 
                           A_neg_shifted_by2_1_59_port, RESULT(122) => 
                           A_neg_shifted_by2_1_58_port, RESULT(121) => 
                           A_neg_shifted_by2_1_57_port, RESULT(120) => 
                           A_neg_shifted_by2_1_56_port, RESULT(119) => 
                           A_neg_shifted_by2_1_55_port, RESULT(118) => 
                           A_neg_shifted_by2_1_54_port, RESULT(117) => 
                           A_neg_shifted_by2_1_53_port, RESULT(116) => 
                           A_neg_shifted_by2_1_52_port, RESULT(115) => 
                           A_neg_shifted_by2_1_51_port, RESULT(114) => 
                           A_neg_shifted_by2_1_50_port, RESULT(113) => 
                           A_neg_shifted_by2_1_49_port, RESULT(112) => 
                           A_neg_shifted_by2_1_48_port, RESULT(111) => 
                           A_neg_shifted_by2_1_47_port, RESULT(110) => 
                           A_neg_shifted_by2_1_46_port, RESULT(109) => 
                           A_neg_shifted_by2_1_45_port, RESULT(108) => 
                           A_neg_shifted_by2_1_44_port, RESULT(107) => 
                           A_neg_shifted_by2_1_43_port, RESULT(106) => 
                           A_neg_shifted_by2_1_42_port, RESULT(105) => 
                           A_neg_shifted_by2_1_41_port, RESULT(104) => 
                           A_neg_shifted_by2_1_40_port, RESULT(103) => 
                           A_neg_shifted_by2_1_39_port, RESULT(102) => 
                           A_neg_shifted_by2_1_38_port, RESULT(101) => 
                           A_neg_shifted_by2_1_37_port, RESULT(100) => 
                           A_neg_shifted_by2_1_36_port, RESULT(99) => 
                           A_neg_shifted_by2_1_35_port, RESULT(98) => 
                           A_neg_shifted_by2_1_34_port, RESULT(97) => 
                           A_neg_shifted_by2_1_33_port, RESULT(96) => 
                           A_neg_shifted_by2_1_32_port, RESULT(95) => 
                           A_neg_shifted_by2_1_31_port, RESULT(94) => 
                           A_neg_shifted_by2_1_30_port, RESULT(93) => 
                           A_neg_shifted_by2_1_29_port, RESULT(92) => 
                           A_neg_shifted_by2_1_28_port, RESULT(91) => 
                           A_neg_shifted_by2_1_27_port, RESULT(90) => 
                           A_neg_shifted_by2_1_26_port, RESULT(89) => 
                           A_neg_shifted_by2_1_25_port, RESULT(88) => 
                           A_neg_shifted_by2_1_24_port, RESULT(87) => 
                           A_neg_shifted_by2_1_23_port, RESULT(86) => 
                           A_neg_shifted_by2_1_22_port, RESULT(85) => 
                           A_neg_shifted_by2_1_21_port, RESULT(84) => 
                           A_neg_shifted_by2_1_20_port, RESULT(83) => 
                           A_neg_shifted_by2_1_19_port, RESULT(82) => 
                           A_neg_shifted_by2_1_18_port, RESULT(81) => 
                           A_neg_shifted_by2_1_17_port, RESULT(80) => 
                           A_neg_shifted_by2_1_16_port, RESULT(79) => 
                           A_neg_shifted_by2_1_15_port, RESULT(78) => 
                           A_neg_shifted_by2_1_14_port, RESULT(77) => 
                           A_neg_shifted_by2_1_13_port, RESULT(76) => 
                           A_neg_shifted_by2_1_12_port, RESULT(75) => 
                           A_neg_shifted_by2_1_11_port, RESULT(74) => 
                           A_neg_shifted_by2_1_10_port, RESULT(73) => 
                           A_neg_shifted_by2_1_9_port, RESULT(72) => 
                           A_neg_shifted_by2_1_8_port, RESULT(71) => 
                           A_neg_shifted_by2_1_7_port, RESULT(70) => 
                           A_neg_shifted_by2_1_6_port, RESULT(69) => 
                           A_neg_shifted_by2_1_5_port, RESULT(68) => 
                           A_neg_shifted_by2_1_4_port, RESULT(67) => 
                           A_neg_shifted_by2_1_3_port, RESULT(66) => 
                           A_neg_shifted_by2_1_2_port, RESULT(65) => n_1173, 
                           RESULT(64) => n_1174, RESULT(63) => 
                           A_neg_shifted_by1_1_63_port, RESULT(62) => 
                           A_neg_shifted_by1_1_62_port, RESULT(61) => 
                           A_neg_shifted_by1_1_61_port, RESULT(60) => 
                           A_neg_shifted_by1_1_60_port, RESULT(59) => 
                           A_neg_shifted_by1_1_59_port, RESULT(58) => 
                           A_neg_shifted_by1_1_58_port, RESULT(57) => 
                           A_neg_shifted_by1_1_57_port, RESULT(56) => 
                           A_neg_shifted_by1_1_56_port, RESULT(55) => 
                           A_neg_shifted_by1_1_55_port, RESULT(54) => 
                           A_neg_shifted_by1_1_54_port, RESULT(53) => 
                           A_neg_shifted_by1_1_53_port, RESULT(52) => 
                           A_neg_shifted_by1_1_52_port, RESULT(51) => 
                           A_neg_shifted_by1_1_51_port, RESULT(50) => 
                           A_neg_shifted_by1_1_50_port, RESULT(49) => 
                           A_neg_shifted_by1_1_49_port, RESULT(48) => 
                           A_neg_shifted_by1_1_48_port, RESULT(47) => 
                           A_neg_shifted_by1_1_47_port, RESULT(46) => 
                           A_neg_shifted_by1_1_46_port, RESULT(45) => 
                           A_neg_shifted_by1_1_45_port, RESULT(44) => 
                           A_neg_shifted_by1_1_44_port, RESULT(43) => 
                           A_neg_shifted_by1_1_43_port, RESULT(42) => 
                           A_neg_shifted_by1_1_42_port, RESULT(41) => 
                           A_neg_shifted_by1_1_41_port, RESULT(40) => 
                           A_neg_shifted_by1_1_40_port, RESULT(39) => 
                           A_neg_shifted_by1_1_39_port, RESULT(38) => 
                           A_neg_shifted_by1_1_38_port, RESULT(37) => 
                           A_neg_shifted_by1_1_37_port, RESULT(36) => 
                           A_neg_shifted_by1_1_36_port, RESULT(35) => 
                           A_neg_shifted_by1_1_35_port, RESULT(34) => 
                           A_neg_shifted_by1_1_34_port, RESULT(33) => 
                           A_neg_shifted_by1_1_33_port, RESULT(32) => 
                           A_neg_shifted_by1_1_32_port, RESULT(31) => 
                           A_neg_shifted_by1_1_31_port, RESULT(30) => 
                           A_neg_shifted_by1_1_30_port, RESULT(29) => 
                           A_neg_shifted_by1_1_29_port, RESULT(28) => 
                           A_neg_shifted_by1_1_28_port, RESULT(27) => 
                           A_neg_shifted_by1_1_27_port, RESULT(26) => 
                           A_neg_shifted_by1_1_26_port, RESULT(25) => 
                           A_neg_shifted_by1_1_25_port, RESULT(24) => 
                           A_neg_shifted_by1_1_24_port, RESULT(23) => 
                           A_neg_shifted_by1_1_23_port, RESULT(22) => 
                           A_neg_shifted_by1_1_22_port, RESULT(21) => 
                           A_neg_shifted_by1_1_21_port, RESULT(20) => 
                           A_neg_shifted_by1_1_20_port, RESULT(19) => 
                           A_neg_shifted_by1_1_19_port, RESULT(18) => 
                           A_neg_shifted_by1_1_18_port, RESULT(17) => 
                           A_neg_shifted_by1_1_17_port, RESULT(16) => 
                           A_neg_shifted_by1_1_16_port, RESULT(15) => 
                           A_neg_shifted_by1_1_15_port, RESULT(14) => 
                           A_neg_shifted_by1_1_14_port, RESULT(13) => 
                           A_neg_shifted_by1_1_13_port, RESULT(12) => 
                           A_neg_shifted_by1_1_12_port, RESULT(11) => 
                           A_neg_shifted_by1_1_11_port, RESULT(10) => 
                           A_neg_shifted_by1_1_10_port, RESULT(9) => 
                           A_neg_shifted_by1_1_9_port, RESULT(8) => 
                           A_neg_shifted_by1_1_8_port, RESULT(7) => 
                           A_neg_shifted_by1_1_7_port, RESULT(6) => 
                           A_neg_shifted_by1_1_6_port, RESULT(5) => 
                           A_neg_shifted_by1_1_5_port, RESULT(4) => 
                           A_neg_shifted_by1_1_4_port, RESULT(3) => 
                           A_neg_shifted_by1_1_3_port, RESULT(2) => 
                           A_neg_shifted_by1_1_2_port, RESULT(1) => 
                           A_neg_shifted_by1_1_1_port, RESULT(0) => n_1175);
   SHIFTERi_2_0 : Shifter_NBIT64_14 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_1_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_1_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_1_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_1_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_1_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_1_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_1_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_1_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_1_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_1_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_1_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_1_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_1_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_1_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_1_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_1_48_port, TO_SHIFT(47) => n206, 
                           TO_SHIFT(46) => A_neg_shifted_by2_1_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_1_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_1_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_1_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_1_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_1_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_1_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_1_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_1_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_1_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_1_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_1_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_1_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_1_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_1_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_1_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_1_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_1_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_1_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_1_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_1_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_1_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_1_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_1_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_1_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_1_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_1_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_1_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_1_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_1_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_1_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_1_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_1_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_1_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_1_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_1_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_1_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_1_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_1_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_1_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_1_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_1_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_1_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_1_3_port, 
                           TO_SHIFT(2) => A_neg_shifted_by2_1_2_port, 
                           TO_SHIFT(1) => A_neg_shifted_by2_1_1_port, 
                           TO_SHIFT(0) => A_neg_shifted_by2_1_0_port, 
                           RESULT(127) => A_neg_shifted_by2_2_63_port, 
                           RESULT(126) => A_neg_shifted_by2_2_62_port, 
                           RESULT(125) => A_neg_shifted_by2_2_61_port, 
                           RESULT(124) => A_neg_shifted_by2_2_60_port, 
                           RESULT(123) => A_neg_shifted_by2_2_59_port, 
                           RESULT(122) => A_neg_shifted_by2_2_58_port, 
                           RESULT(121) => A_neg_shifted_by2_2_57_port, 
                           RESULT(120) => A_neg_shifted_by2_2_56_port, 
                           RESULT(119) => A_neg_shifted_by2_2_55_port, 
                           RESULT(118) => A_neg_shifted_by2_2_54_port, 
                           RESULT(117) => A_neg_shifted_by2_2_53_port, 
                           RESULT(116) => A_neg_shifted_by2_2_52_port, 
                           RESULT(115) => A_neg_shifted_by2_2_51_port, 
                           RESULT(114) => A_neg_shifted_by2_2_50_port, 
                           RESULT(113) => A_neg_shifted_by2_2_49_port, 
                           RESULT(112) => A_neg_shifted_by2_2_48_port, 
                           RESULT(111) => A_neg_shifted_by2_2_47_port, 
                           RESULT(110) => A_neg_shifted_by2_2_46_port, 
                           RESULT(109) => A_neg_shifted_by2_2_45_port, 
                           RESULT(108) => A_neg_shifted_by2_2_44_port, 
                           RESULT(107) => A_neg_shifted_by2_2_43_port, 
                           RESULT(106) => A_neg_shifted_by2_2_42_port, 
                           RESULT(105) => A_neg_shifted_by2_2_41_port, 
                           RESULT(104) => A_neg_shifted_by2_2_40_port, 
                           RESULT(103) => A_neg_shifted_by2_2_39_port, 
                           RESULT(102) => A_neg_shifted_by2_2_38_port, 
                           RESULT(101) => A_neg_shifted_by2_2_37_port, 
                           RESULT(100) => A_neg_shifted_by2_2_36_port, 
                           RESULT(99) => A_neg_shifted_by2_2_35_port, 
                           RESULT(98) => A_neg_shifted_by2_2_34_port, 
                           RESULT(97) => A_neg_shifted_by2_2_33_port, 
                           RESULT(96) => A_neg_shifted_by2_2_32_port, 
                           RESULT(95) => A_neg_shifted_by2_2_31_port, 
                           RESULT(94) => A_neg_shifted_by2_2_30_port, 
                           RESULT(93) => A_neg_shifted_by2_2_29_port, 
                           RESULT(92) => A_neg_shifted_by2_2_28_port, 
                           RESULT(91) => A_neg_shifted_by2_2_27_port, 
                           RESULT(90) => A_neg_shifted_by2_2_26_port, 
                           RESULT(89) => A_neg_shifted_by2_2_25_port, 
                           RESULT(88) => A_neg_shifted_by2_2_24_port, 
                           RESULT(87) => A_neg_shifted_by2_2_23_port, 
                           RESULT(86) => A_neg_shifted_by2_2_22_port, 
                           RESULT(85) => A_neg_shifted_by2_2_21_port, 
                           RESULT(84) => A_neg_shifted_by2_2_20_port, 
                           RESULT(83) => A_neg_shifted_by2_2_19_port, 
                           RESULT(82) => A_neg_shifted_by2_2_18_port, 
                           RESULT(81) => A_neg_shifted_by2_2_17_port, 
                           RESULT(80) => A_neg_shifted_by2_2_16_port, 
                           RESULT(79) => A_neg_shifted_by2_2_15_port, 
                           RESULT(78) => A_neg_shifted_by2_2_14_port, 
                           RESULT(77) => A_neg_shifted_by2_2_13_port, 
                           RESULT(76) => A_neg_shifted_by2_2_12_port, 
                           RESULT(75) => A_neg_shifted_by2_2_11_port, 
                           RESULT(74) => A_neg_shifted_by2_2_10_port, 
                           RESULT(73) => A_neg_shifted_by2_2_9_port, RESULT(72)
                           => A_neg_shifted_by2_2_8_port, RESULT(71) => 
                           A_neg_shifted_by2_2_7_port, RESULT(70) => 
                           A_neg_shifted_by2_2_6_port, RESULT(69) => 
                           A_neg_shifted_by2_2_5_port, RESULT(68) => 
                           A_neg_shifted_by2_2_4_port, RESULT(67) => 
                           A_neg_shifted_by2_2_3_port, RESULT(66) => 
                           A_neg_shifted_by2_2_2_port, RESULT(65) => n_1176, 
                           RESULT(64) => n_1177, RESULT(63) => 
                           A_neg_shifted_by1_2_63_port, RESULT(62) => 
                           A_neg_shifted_by1_2_62_port, RESULT(61) => 
                           A_neg_shifted_by1_2_61_port, RESULT(60) => 
                           A_neg_shifted_by1_2_60_port, RESULT(59) => 
                           A_neg_shifted_by1_2_59_port, RESULT(58) => 
                           A_neg_shifted_by1_2_58_port, RESULT(57) => 
                           A_neg_shifted_by1_2_57_port, RESULT(56) => 
                           A_neg_shifted_by1_2_56_port, RESULT(55) => 
                           A_neg_shifted_by1_2_55_port, RESULT(54) => 
                           A_neg_shifted_by1_2_54_port, RESULT(53) => 
                           A_neg_shifted_by1_2_53_port, RESULT(52) => 
                           A_neg_shifted_by1_2_52_port, RESULT(51) => 
                           A_neg_shifted_by1_2_51_port, RESULT(50) => 
                           A_neg_shifted_by1_2_50_port, RESULT(49) => 
                           A_neg_shifted_by1_2_49_port, RESULT(48) => 
                           A_neg_shifted_by1_2_48_port, RESULT(47) => 
                           A_neg_shifted_by1_2_47_port, RESULT(46) => 
                           A_neg_shifted_by1_2_46_port, RESULT(45) => 
                           A_neg_shifted_by1_2_45_port, RESULT(44) => 
                           A_neg_shifted_by1_2_44_port, RESULT(43) => 
                           A_neg_shifted_by1_2_43_port, RESULT(42) => 
                           A_neg_shifted_by1_2_42_port, RESULT(41) => 
                           A_neg_shifted_by1_2_41_port, RESULT(40) => 
                           A_neg_shifted_by1_2_40_port, RESULT(39) => 
                           A_neg_shifted_by1_2_39_port, RESULT(38) => 
                           A_neg_shifted_by1_2_38_port, RESULT(37) => 
                           A_neg_shifted_by1_2_37_port, RESULT(36) => 
                           A_neg_shifted_by1_2_36_port, RESULT(35) => 
                           A_neg_shifted_by1_2_35_port, RESULT(34) => 
                           A_neg_shifted_by1_2_34_port, RESULT(33) => 
                           A_neg_shifted_by1_2_33_port, RESULT(32) => 
                           A_neg_shifted_by1_2_32_port, RESULT(31) => 
                           A_neg_shifted_by1_2_31_port, RESULT(30) => 
                           A_neg_shifted_by1_2_30_port, RESULT(29) => 
                           A_neg_shifted_by1_2_29_port, RESULT(28) => 
                           A_neg_shifted_by1_2_28_port, RESULT(27) => 
                           A_neg_shifted_by1_2_27_port, RESULT(26) => 
                           A_neg_shifted_by1_2_26_port, RESULT(25) => 
                           A_neg_shifted_by1_2_25_port, RESULT(24) => 
                           A_neg_shifted_by1_2_24_port, RESULT(23) => 
                           A_neg_shifted_by1_2_23_port, RESULT(22) => 
                           A_neg_shifted_by1_2_22_port, RESULT(21) => 
                           A_neg_shifted_by1_2_21_port, RESULT(20) => 
                           A_neg_shifted_by1_2_20_port, RESULT(19) => 
                           A_neg_shifted_by1_2_19_port, RESULT(18) => 
                           A_neg_shifted_by1_2_18_port, RESULT(17) => 
                           A_neg_shifted_by1_2_17_port, RESULT(16) => 
                           A_neg_shifted_by1_2_16_port, RESULT(15) => 
                           A_neg_shifted_by1_2_15_port, RESULT(14) => 
                           A_neg_shifted_by1_2_14_port, RESULT(13) => 
                           A_neg_shifted_by1_2_13_port, RESULT(12) => 
                           A_neg_shifted_by1_2_12_port, RESULT(11) => 
                           A_neg_shifted_by1_2_11_port, RESULT(10) => 
                           A_neg_shifted_by1_2_10_port, RESULT(9) => 
                           A_neg_shifted_by1_2_9_port, RESULT(8) => 
                           A_neg_shifted_by1_2_8_port, RESULT(7) => 
                           A_neg_shifted_by1_2_7_port, RESULT(6) => 
                           A_neg_shifted_by1_2_6_port, RESULT(5) => 
                           A_neg_shifted_by1_2_5_port, RESULT(4) => 
                           A_neg_shifted_by1_2_4_port, RESULT(3) => 
                           A_neg_shifted_by1_2_3_port, RESULT(2) => 
                           A_neg_shifted_by1_2_2_port, RESULT(1) => 
                           A_neg_shifted_by1_2_1_port, RESULT(0) => n_1178);
   SHIFTERi_3_0 : Shifter_NBIT64_13 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_2_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_2_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_2_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_2_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_2_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_2_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_2_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_2_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_2_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_2_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_2_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_2_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_2_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_2_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_2_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_2_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_2_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_2_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_2_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_2_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_2_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_2_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_2_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_2_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_2_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_2_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_2_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_2_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_2_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_2_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_2_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_2_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_2_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_2_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_2_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_2_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_2_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_2_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_2_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_2_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_2_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_2_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_2_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_2_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_2_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_2_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_2_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_2_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_2_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_2_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_2_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_2_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_2_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_2_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_2_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_2_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_2_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_2_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_2_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_2_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_2_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_2_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_2_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_2_0_port, RESULT(127) => 
                           A_neg_shifted_by2_3_63_port, RESULT(126) => 
                           A_neg_shifted_by2_3_62_port, RESULT(125) => 
                           A_neg_shifted_by2_3_61_port, RESULT(124) => 
                           A_neg_shifted_by2_3_60_port, RESULT(123) => 
                           A_neg_shifted_by2_3_59_port, RESULT(122) => 
                           A_neg_shifted_by2_3_58_port, RESULT(121) => 
                           A_neg_shifted_by2_3_57_port, RESULT(120) => 
                           A_neg_shifted_by2_3_56_port, RESULT(119) => 
                           A_neg_shifted_by2_3_55_port, RESULT(118) => 
                           A_neg_shifted_by2_3_54_port, RESULT(117) => 
                           A_neg_shifted_by2_3_53_port, RESULT(116) => 
                           A_neg_shifted_by2_3_52_port, RESULT(115) => 
                           A_neg_shifted_by2_3_51_port, RESULT(114) => 
                           A_neg_shifted_by2_3_50_port, RESULT(113) => 
                           A_neg_shifted_by2_3_49_port, RESULT(112) => 
                           A_neg_shifted_by2_3_48_port, RESULT(111) => 
                           A_neg_shifted_by2_3_47_port, RESULT(110) => 
                           A_neg_shifted_by2_3_46_port, RESULT(109) => 
                           A_neg_shifted_by2_3_45_port, RESULT(108) => 
                           A_neg_shifted_by2_3_44_port, RESULT(107) => 
                           A_neg_shifted_by2_3_43_port, RESULT(106) => 
                           A_neg_shifted_by2_3_42_port, RESULT(105) => 
                           A_neg_shifted_by2_3_41_port, RESULT(104) => 
                           A_neg_shifted_by2_3_40_port, RESULT(103) => 
                           A_neg_shifted_by2_3_39_port, RESULT(102) => 
                           A_neg_shifted_by2_3_38_port, RESULT(101) => 
                           A_neg_shifted_by2_3_37_port, RESULT(100) => 
                           A_neg_shifted_by2_3_36_port, RESULT(99) => 
                           A_neg_shifted_by2_3_35_port, RESULT(98) => 
                           A_neg_shifted_by2_3_34_port, RESULT(97) => 
                           A_neg_shifted_by2_3_33_port, RESULT(96) => 
                           A_neg_shifted_by2_3_32_port, RESULT(95) => 
                           A_neg_shifted_by2_3_31_port, RESULT(94) => 
                           A_neg_shifted_by2_3_30_port, RESULT(93) => 
                           A_neg_shifted_by2_3_29_port, RESULT(92) => 
                           A_neg_shifted_by2_3_28_port, RESULT(91) => 
                           A_neg_shifted_by2_3_27_port, RESULT(90) => 
                           A_neg_shifted_by2_3_26_port, RESULT(89) => 
                           A_neg_shifted_by2_3_25_port, RESULT(88) => 
                           A_neg_shifted_by2_3_24_port, RESULT(87) => 
                           A_neg_shifted_by2_3_23_port, RESULT(86) => 
                           A_neg_shifted_by2_3_22_port, RESULT(85) => 
                           A_neg_shifted_by2_3_21_port, RESULT(84) => 
                           A_neg_shifted_by2_3_20_port, RESULT(83) => 
                           A_neg_shifted_by2_3_19_port, RESULT(82) => 
                           A_neg_shifted_by2_3_18_port, RESULT(81) => 
                           A_neg_shifted_by2_3_17_port, RESULT(80) => 
                           A_neg_shifted_by2_3_16_port, RESULT(79) => 
                           A_neg_shifted_by2_3_15_port, RESULT(78) => 
                           A_neg_shifted_by2_3_14_port, RESULT(77) => 
                           A_neg_shifted_by2_3_13_port, RESULT(76) => 
                           A_neg_shifted_by2_3_12_port, RESULT(75) => 
                           A_neg_shifted_by2_3_11_port, RESULT(74) => 
                           A_neg_shifted_by2_3_10_port, RESULT(73) => 
                           A_neg_shifted_by2_3_9_port, RESULT(72) => 
                           A_neg_shifted_by2_3_8_port, RESULT(71) => 
                           A_neg_shifted_by2_3_7_port, RESULT(70) => 
                           A_neg_shifted_by2_3_6_port, RESULT(69) => 
                           A_neg_shifted_by2_3_5_port, RESULT(68) => 
                           A_neg_shifted_by2_3_4_port, RESULT(67) => 
                           A_neg_shifted_by2_3_3_port, RESULT(66) => 
                           A_neg_shifted_by2_3_2_port, RESULT(65) => n_1179, 
                           RESULT(64) => n_1180, RESULT(63) => 
                           A_neg_shifted_by1_3_63_port, RESULT(62) => 
                           A_neg_shifted_by1_3_62_port, RESULT(61) => 
                           A_neg_shifted_by1_3_61_port, RESULT(60) => 
                           A_neg_shifted_by1_3_60_port, RESULT(59) => 
                           A_neg_shifted_by1_3_59_port, RESULT(58) => 
                           A_neg_shifted_by1_3_58_port, RESULT(57) => 
                           A_neg_shifted_by1_3_57_port, RESULT(56) => 
                           A_neg_shifted_by1_3_56_port, RESULT(55) => 
                           A_neg_shifted_by1_3_55_port, RESULT(54) => 
                           A_neg_shifted_by1_3_54_port, RESULT(53) => 
                           A_neg_shifted_by1_3_53_port, RESULT(52) => 
                           A_neg_shifted_by1_3_52_port, RESULT(51) => 
                           A_neg_shifted_by1_3_51_port, RESULT(50) => 
                           A_neg_shifted_by1_3_50_port, RESULT(49) => 
                           A_neg_shifted_by1_3_49_port, RESULT(48) => 
                           A_neg_shifted_by1_3_48_port, RESULT(47) => 
                           A_neg_shifted_by1_3_47_port, RESULT(46) => 
                           A_neg_shifted_by1_3_46_port, RESULT(45) => 
                           A_neg_shifted_by1_3_45_port, RESULT(44) => 
                           A_neg_shifted_by1_3_44_port, RESULT(43) => 
                           A_neg_shifted_by1_3_43_port, RESULT(42) => 
                           A_neg_shifted_by1_3_42_port, RESULT(41) => 
                           A_neg_shifted_by1_3_41_port, RESULT(40) => 
                           A_neg_shifted_by1_3_40_port, RESULT(39) => 
                           A_neg_shifted_by1_3_39_port, RESULT(38) => 
                           A_neg_shifted_by1_3_38_port, RESULT(37) => 
                           A_neg_shifted_by1_3_37_port, RESULT(36) => 
                           A_neg_shifted_by1_3_36_port, RESULT(35) => 
                           A_neg_shifted_by1_3_35_port, RESULT(34) => 
                           A_neg_shifted_by1_3_34_port, RESULT(33) => 
                           A_neg_shifted_by1_3_33_port, RESULT(32) => 
                           A_neg_shifted_by1_3_32_port, RESULT(31) => 
                           A_neg_shifted_by1_3_31_port, RESULT(30) => 
                           A_neg_shifted_by1_3_30_port, RESULT(29) => 
                           A_neg_shifted_by1_3_29_port, RESULT(28) => 
                           A_neg_shifted_by1_3_28_port, RESULT(27) => 
                           A_neg_shifted_by1_3_27_port, RESULT(26) => 
                           A_neg_shifted_by1_3_26_port, RESULT(25) => 
                           A_neg_shifted_by1_3_25_port, RESULT(24) => 
                           A_neg_shifted_by1_3_24_port, RESULT(23) => 
                           A_neg_shifted_by1_3_23_port, RESULT(22) => 
                           A_neg_shifted_by1_3_22_port, RESULT(21) => 
                           A_neg_shifted_by1_3_21_port, RESULT(20) => 
                           A_neg_shifted_by1_3_20_port, RESULT(19) => 
                           A_neg_shifted_by1_3_19_port, RESULT(18) => 
                           A_neg_shifted_by1_3_18_port, RESULT(17) => 
                           A_neg_shifted_by1_3_17_port, RESULT(16) => 
                           A_neg_shifted_by1_3_16_port, RESULT(15) => 
                           A_neg_shifted_by1_3_15_port, RESULT(14) => 
                           A_neg_shifted_by1_3_14_port, RESULT(13) => 
                           A_neg_shifted_by1_3_13_port, RESULT(12) => 
                           A_neg_shifted_by1_3_12_port, RESULT(11) => 
                           A_neg_shifted_by1_3_11_port, RESULT(10) => 
                           A_neg_shifted_by1_3_10_port, RESULT(9) => 
                           A_neg_shifted_by1_3_9_port, RESULT(8) => 
                           A_neg_shifted_by1_3_8_port, RESULT(7) => 
                           A_neg_shifted_by1_3_7_port, RESULT(6) => 
                           A_neg_shifted_by1_3_6_port, RESULT(5) => 
                           A_neg_shifted_by1_3_5_port, RESULT(4) => 
                           A_neg_shifted_by1_3_4_port, RESULT(3) => 
                           A_neg_shifted_by1_3_3_port, RESULT(2) => 
                           A_neg_shifted_by1_3_2_port, RESULT(1) => 
                           A_neg_shifted_by1_3_1_port, RESULT(0) => n_1181);
   SHIFTERi_4_0 : Shifter_NBIT64_12 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_3_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_3_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_3_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_3_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_3_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_3_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_3_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_3_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_3_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_3_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_3_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_3_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_3_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_3_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_3_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_3_48_port, TO_SHIFT(47) => n205, 
                           TO_SHIFT(46) => A_neg_shifted_by2_3_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_3_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_3_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_3_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_3_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_3_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_3_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_3_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_3_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_3_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_3_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_3_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_3_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_3_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_3_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_3_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_3_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_3_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_3_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_3_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_3_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_3_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_3_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_3_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_3_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_3_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_3_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_3_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_3_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_3_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_3_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_3_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_3_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_3_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_3_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_3_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_3_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_3_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_3_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_3_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_3_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_3_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_3_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_3_3_port, 
                           TO_SHIFT(2) => A_neg_shifted_by2_3_2_port, 
                           TO_SHIFT(1) => A_neg_shifted_by2_3_1_port, 
                           TO_SHIFT(0) => A_neg_shifted_by2_3_0_port, 
                           RESULT(127) => A_neg_shifted_by2_4_63_port, 
                           RESULT(126) => A_neg_shifted_by2_4_62_port, 
                           RESULT(125) => A_neg_shifted_by2_4_61_port, 
                           RESULT(124) => A_neg_shifted_by2_4_60_port, 
                           RESULT(123) => A_neg_shifted_by2_4_59_port, 
                           RESULT(122) => A_neg_shifted_by2_4_58_port, 
                           RESULT(121) => A_neg_shifted_by2_4_57_port, 
                           RESULT(120) => A_neg_shifted_by2_4_56_port, 
                           RESULT(119) => A_neg_shifted_by2_4_55_port, 
                           RESULT(118) => A_neg_shifted_by2_4_54_port, 
                           RESULT(117) => A_neg_shifted_by2_4_53_port, 
                           RESULT(116) => A_neg_shifted_by2_4_52_port, 
                           RESULT(115) => A_neg_shifted_by2_4_51_port, 
                           RESULT(114) => A_neg_shifted_by2_4_50_port, 
                           RESULT(113) => A_neg_shifted_by2_4_49_port, 
                           RESULT(112) => A_neg_shifted_by2_4_48_port, 
                           RESULT(111) => A_neg_shifted_by2_4_47_port, 
                           RESULT(110) => A_neg_shifted_by2_4_46_port, 
                           RESULT(109) => A_neg_shifted_by2_4_45_port, 
                           RESULT(108) => A_neg_shifted_by2_4_44_port, 
                           RESULT(107) => A_neg_shifted_by2_4_43_port, 
                           RESULT(106) => A_neg_shifted_by2_4_42_port, 
                           RESULT(105) => A_neg_shifted_by2_4_41_port, 
                           RESULT(104) => A_neg_shifted_by2_4_40_port, 
                           RESULT(103) => A_neg_shifted_by2_4_39_port, 
                           RESULT(102) => A_neg_shifted_by2_4_38_port, 
                           RESULT(101) => A_neg_shifted_by2_4_37_port, 
                           RESULT(100) => A_neg_shifted_by2_4_36_port, 
                           RESULT(99) => A_neg_shifted_by2_4_35_port, 
                           RESULT(98) => A_neg_shifted_by2_4_34_port, 
                           RESULT(97) => A_neg_shifted_by2_4_33_port, 
                           RESULT(96) => A_neg_shifted_by2_4_32_port, 
                           RESULT(95) => A_neg_shifted_by2_4_31_port, 
                           RESULT(94) => A_neg_shifted_by2_4_30_port, 
                           RESULT(93) => A_neg_shifted_by2_4_29_port, 
                           RESULT(92) => A_neg_shifted_by2_4_28_port, 
                           RESULT(91) => A_neg_shifted_by2_4_27_port, 
                           RESULT(90) => A_neg_shifted_by2_4_26_port, 
                           RESULT(89) => A_neg_shifted_by2_4_25_port, 
                           RESULT(88) => A_neg_shifted_by2_4_24_port, 
                           RESULT(87) => A_neg_shifted_by2_4_23_port, 
                           RESULT(86) => A_neg_shifted_by2_4_22_port, 
                           RESULT(85) => A_neg_shifted_by2_4_21_port, 
                           RESULT(84) => A_neg_shifted_by2_4_20_port, 
                           RESULT(83) => A_neg_shifted_by2_4_19_port, 
                           RESULT(82) => A_neg_shifted_by2_4_18_port, 
                           RESULT(81) => A_neg_shifted_by2_4_17_port, 
                           RESULT(80) => A_neg_shifted_by2_4_16_port, 
                           RESULT(79) => A_neg_shifted_by2_4_15_port, 
                           RESULT(78) => A_neg_shifted_by2_4_14_port, 
                           RESULT(77) => A_neg_shifted_by2_4_13_port, 
                           RESULT(76) => A_neg_shifted_by2_4_12_port, 
                           RESULT(75) => A_neg_shifted_by2_4_11_port, 
                           RESULT(74) => A_neg_shifted_by2_4_10_port, 
                           RESULT(73) => A_neg_shifted_by2_4_9_port, RESULT(72)
                           => A_neg_shifted_by2_4_8_port, RESULT(71) => 
                           A_neg_shifted_by2_4_7_port, RESULT(70) => 
                           A_neg_shifted_by2_4_6_port, RESULT(69) => 
                           A_neg_shifted_by2_4_5_port, RESULT(68) => 
                           A_neg_shifted_by2_4_4_port, RESULT(67) => 
                           A_neg_shifted_by2_4_3_port, RESULT(66) => 
                           A_neg_shifted_by2_4_2_port, RESULT(65) => n_1182, 
                           RESULT(64) => n_1183, RESULT(63) => 
                           A_neg_shifted_by1_4_63_port, RESULT(62) => 
                           A_neg_shifted_by1_4_62_port, RESULT(61) => 
                           A_neg_shifted_by1_4_61_port, RESULT(60) => 
                           A_neg_shifted_by1_4_60_port, RESULT(59) => 
                           A_neg_shifted_by1_4_59_port, RESULT(58) => 
                           A_neg_shifted_by1_4_58_port, RESULT(57) => 
                           A_neg_shifted_by1_4_57_port, RESULT(56) => 
                           A_neg_shifted_by1_4_56_port, RESULT(55) => 
                           A_neg_shifted_by1_4_55_port, RESULT(54) => 
                           A_neg_shifted_by1_4_54_port, RESULT(53) => 
                           A_neg_shifted_by1_4_53_port, RESULT(52) => 
                           A_neg_shifted_by1_4_52_port, RESULT(51) => 
                           A_neg_shifted_by1_4_51_port, RESULT(50) => 
                           A_neg_shifted_by1_4_50_port, RESULT(49) => 
                           A_neg_shifted_by1_4_49_port, RESULT(48) => 
                           A_neg_shifted_by1_4_48_port, RESULT(47) => 
                           A_neg_shifted_by1_4_47_port, RESULT(46) => 
                           A_neg_shifted_by1_4_46_port, RESULT(45) => 
                           A_neg_shifted_by1_4_45_port, RESULT(44) => 
                           A_neg_shifted_by1_4_44_port, RESULT(43) => 
                           A_neg_shifted_by1_4_43_port, RESULT(42) => 
                           A_neg_shifted_by1_4_42_port, RESULT(41) => 
                           A_neg_shifted_by1_4_41_port, RESULT(40) => 
                           A_neg_shifted_by1_4_40_port, RESULT(39) => 
                           A_neg_shifted_by1_4_39_port, RESULT(38) => 
                           A_neg_shifted_by1_4_38_port, RESULT(37) => 
                           A_neg_shifted_by1_4_37_port, RESULT(36) => 
                           A_neg_shifted_by1_4_36_port, RESULT(35) => 
                           A_neg_shifted_by1_4_35_port, RESULT(34) => 
                           A_neg_shifted_by1_4_34_port, RESULT(33) => 
                           A_neg_shifted_by1_4_33_port, RESULT(32) => 
                           A_neg_shifted_by1_4_32_port, RESULT(31) => 
                           A_neg_shifted_by1_4_31_port, RESULT(30) => 
                           A_neg_shifted_by1_4_30_port, RESULT(29) => 
                           A_neg_shifted_by1_4_29_port, RESULT(28) => 
                           A_neg_shifted_by1_4_28_port, RESULT(27) => 
                           A_neg_shifted_by1_4_27_port, RESULT(26) => 
                           A_neg_shifted_by1_4_26_port, RESULT(25) => 
                           A_neg_shifted_by1_4_25_port, RESULT(24) => 
                           A_neg_shifted_by1_4_24_port, RESULT(23) => 
                           A_neg_shifted_by1_4_23_port, RESULT(22) => 
                           A_neg_shifted_by1_4_22_port, RESULT(21) => 
                           A_neg_shifted_by1_4_21_port, RESULT(20) => 
                           A_neg_shifted_by1_4_20_port, RESULT(19) => 
                           A_neg_shifted_by1_4_19_port, RESULT(18) => 
                           A_neg_shifted_by1_4_18_port, RESULT(17) => 
                           A_neg_shifted_by1_4_17_port, RESULT(16) => 
                           A_neg_shifted_by1_4_16_port, RESULT(15) => 
                           A_neg_shifted_by1_4_15_port, RESULT(14) => 
                           A_neg_shifted_by1_4_14_port, RESULT(13) => 
                           A_neg_shifted_by1_4_13_port, RESULT(12) => 
                           A_neg_shifted_by1_4_12_port, RESULT(11) => 
                           A_neg_shifted_by1_4_11_port, RESULT(10) => 
                           A_neg_shifted_by1_4_10_port, RESULT(9) => 
                           A_neg_shifted_by1_4_9_port, RESULT(8) => 
                           A_neg_shifted_by1_4_8_port, RESULT(7) => 
                           A_neg_shifted_by1_4_7_port, RESULT(6) => 
                           A_neg_shifted_by1_4_6_port, RESULT(5) => 
                           A_neg_shifted_by1_4_5_port, RESULT(4) => 
                           A_neg_shifted_by1_4_4_port, RESULT(3) => 
                           A_neg_shifted_by1_4_3_port, RESULT(2) => 
                           A_neg_shifted_by1_4_2_port, RESULT(1) => 
                           A_neg_shifted_by1_4_1_port, RESULT(0) => n_1184);
   SHIFTERi_5_0 : Shifter_NBIT64_11 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_4_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_4_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_4_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_4_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_4_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_4_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_4_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_4_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_4_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_4_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_4_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_4_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_4_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_4_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_4_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_4_48_port, TO_SHIFT(47) => n204, 
                           TO_SHIFT(46) => A_neg_shifted_by2_4_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_4_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_4_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_4_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_4_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_4_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_4_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_4_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_4_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_4_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_4_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_4_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_4_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_4_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_4_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_4_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_4_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_4_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_4_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_4_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_4_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_4_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_4_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_4_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_4_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_4_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_4_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_4_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_4_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_4_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_4_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_4_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_4_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_4_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_4_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_4_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_4_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_4_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_4_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_4_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_4_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_4_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_4_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_4_3_port, 
                           TO_SHIFT(2) => A_neg_shifted_by2_4_2_port, 
                           TO_SHIFT(1) => A_neg_shifted_by2_4_1_port, 
                           TO_SHIFT(0) => A_neg_shifted_by2_4_0_port, 
                           RESULT(127) => A_neg_shifted_by2_5_63_port, 
                           RESULT(126) => A_neg_shifted_by2_5_62_port, 
                           RESULT(125) => A_neg_shifted_by2_5_61_port, 
                           RESULT(124) => A_neg_shifted_by2_5_60_port, 
                           RESULT(123) => A_neg_shifted_by2_5_59_port, 
                           RESULT(122) => A_neg_shifted_by2_5_58_port, 
                           RESULT(121) => A_neg_shifted_by2_5_57_port, 
                           RESULT(120) => A_neg_shifted_by2_5_56_port, 
                           RESULT(119) => A_neg_shifted_by2_5_55_port, 
                           RESULT(118) => A_neg_shifted_by2_5_54_port, 
                           RESULT(117) => A_neg_shifted_by2_5_53_port, 
                           RESULT(116) => A_neg_shifted_by2_5_52_port, 
                           RESULT(115) => A_neg_shifted_by2_5_51_port, 
                           RESULT(114) => A_neg_shifted_by2_5_50_port, 
                           RESULT(113) => A_neg_shifted_by2_5_49_port, 
                           RESULT(112) => A_neg_shifted_by2_5_48_port, 
                           RESULT(111) => A_neg_shifted_by2_5_47_port, 
                           RESULT(110) => A_neg_shifted_by2_5_46_port, 
                           RESULT(109) => A_neg_shifted_by2_5_45_port, 
                           RESULT(108) => A_neg_shifted_by2_5_44_port, 
                           RESULT(107) => A_neg_shifted_by2_5_43_port, 
                           RESULT(106) => A_neg_shifted_by2_5_42_port, 
                           RESULT(105) => A_neg_shifted_by2_5_41_port, 
                           RESULT(104) => A_neg_shifted_by2_5_40_port, 
                           RESULT(103) => A_neg_shifted_by2_5_39_port, 
                           RESULT(102) => A_neg_shifted_by2_5_38_port, 
                           RESULT(101) => A_neg_shifted_by2_5_37_port, 
                           RESULT(100) => A_neg_shifted_by2_5_36_port, 
                           RESULT(99) => A_neg_shifted_by2_5_35_port, 
                           RESULT(98) => A_neg_shifted_by2_5_34_port, 
                           RESULT(97) => A_neg_shifted_by2_5_33_port, 
                           RESULT(96) => A_neg_shifted_by2_5_32_port, 
                           RESULT(95) => A_neg_shifted_by2_5_31_port, 
                           RESULT(94) => A_neg_shifted_by2_5_30_port, 
                           RESULT(93) => A_neg_shifted_by2_5_29_port, 
                           RESULT(92) => A_neg_shifted_by2_5_28_port, 
                           RESULT(91) => A_neg_shifted_by2_5_27_port, 
                           RESULT(90) => A_neg_shifted_by2_5_26_port, 
                           RESULT(89) => A_neg_shifted_by2_5_25_port, 
                           RESULT(88) => A_neg_shifted_by2_5_24_port, 
                           RESULT(87) => A_neg_shifted_by2_5_23_port, 
                           RESULT(86) => A_neg_shifted_by2_5_22_port, 
                           RESULT(85) => A_neg_shifted_by2_5_21_port, 
                           RESULT(84) => A_neg_shifted_by2_5_20_port, 
                           RESULT(83) => A_neg_shifted_by2_5_19_port, 
                           RESULT(82) => A_neg_shifted_by2_5_18_port, 
                           RESULT(81) => A_neg_shifted_by2_5_17_port, 
                           RESULT(80) => A_neg_shifted_by2_5_16_port, 
                           RESULT(79) => A_neg_shifted_by2_5_15_port, 
                           RESULT(78) => A_neg_shifted_by2_5_14_port, 
                           RESULT(77) => A_neg_shifted_by2_5_13_port, 
                           RESULT(76) => A_neg_shifted_by2_5_12_port, 
                           RESULT(75) => A_neg_shifted_by2_5_11_port, 
                           RESULT(74) => A_neg_shifted_by2_5_10_port, 
                           RESULT(73) => A_neg_shifted_by2_5_9_port, RESULT(72)
                           => A_neg_shifted_by2_5_8_port, RESULT(71) => 
                           A_neg_shifted_by2_5_7_port, RESULT(70) => 
                           A_neg_shifted_by2_5_6_port, RESULT(69) => 
                           A_neg_shifted_by2_5_5_port, RESULT(68) => 
                           A_neg_shifted_by2_5_4_port, RESULT(67) => 
                           A_neg_shifted_by2_5_3_port, RESULT(66) => 
                           A_neg_shifted_by2_5_2_port, RESULT(65) => n_1185, 
                           RESULT(64) => n_1186, RESULT(63) => 
                           A_neg_shifted_by1_5_63_port, RESULT(62) => 
                           A_neg_shifted_by1_5_62_port, RESULT(61) => 
                           A_neg_shifted_by1_5_61_port, RESULT(60) => 
                           A_neg_shifted_by1_5_60_port, RESULT(59) => 
                           A_neg_shifted_by1_5_59_port, RESULT(58) => 
                           A_neg_shifted_by1_5_58_port, RESULT(57) => 
                           A_neg_shifted_by1_5_57_port, RESULT(56) => 
                           A_neg_shifted_by1_5_56_port, RESULT(55) => 
                           A_neg_shifted_by1_5_55_port, RESULT(54) => 
                           A_neg_shifted_by1_5_54_port, RESULT(53) => 
                           A_neg_shifted_by1_5_53_port, RESULT(52) => 
                           A_neg_shifted_by1_5_52_port, RESULT(51) => 
                           A_neg_shifted_by1_5_51_port, RESULT(50) => 
                           A_neg_shifted_by1_5_50_port, RESULT(49) => 
                           A_neg_shifted_by1_5_49_port, RESULT(48) => 
                           A_neg_shifted_by1_5_48_port, RESULT(47) => 
                           A_neg_shifted_by1_5_47_port, RESULT(46) => 
                           A_neg_shifted_by1_5_46_port, RESULT(45) => 
                           A_neg_shifted_by1_5_45_port, RESULT(44) => 
                           A_neg_shifted_by1_5_44_port, RESULT(43) => 
                           A_neg_shifted_by1_5_43_port, RESULT(42) => 
                           A_neg_shifted_by1_5_42_port, RESULT(41) => 
                           A_neg_shifted_by1_5_41_port, RESULT(40) => 
                           A_neg_shifted_by1_5_40_port, RESULT(39) => 
                           A_neg_shifted_by1_5_39_port, RESULT(38) => 
                           A_neg_shifted_by1_5_38_port, RESULT(37) => 
                           A_neg_shifted_by1_5_37_port, RESULT(36) => 
                           A_neg_shifted_by1_5_36_port, RESULT(35) => 
                           A_neg_shifted_by1_5_35_port, RESULT(34) => 
                           A_neg_shifted_by1_5_34_port, RESULT(33) => 
                           A_neg_shifted_by1_5_33_port, RESULT(32) => 
                           A_neg_shifted_by1_5_32_port, RESULT(31) => 
                           A_neg_shifted_by1_5_31_port, RESULT(30) => 
                           A_neg_shifted_by1_5_30_port, RESULT(29) => 
                           A_neg_shifted_by1_5_29_port, RESULT(28) => 
                           A_neg_shifted_by1_5_28_port, RESULT(27) => 
                           A_neg_shifted_by1_5_27_port, RESULT(26) => 
                           A_neg_shifted_by1_5_26_port, RESULT(25) => 
                           A_neg_shifted_by1_5_25_port, RESULT(24) => 
                           A_neg_shifted_by1_5_24_port, RESULT(23) => 
                           A_neg_shifted_by1_5_23_port, RESULT(22) => 
                           A_neg_shifted_by1_5_22_port, RESULT(21) => 
                           A_neg_shifted_by1_5_21_port, RESULT(20) => 
                           A_neg_shifted_by1_5_20_port, RESULT(19) => 
                           A_neg_shifted_by1_5_19_port, RESULT(18) => 
                           A_neg_shifted_by1_5_18_port, RESULT(17) => 
                           A_neg_shifted_by1_5_17_port, RESULT(16) => 
                           A_neg_shifted_by1_5_16_port, RESULT(15) => 
                           A_neg_shifted_by1_5_15_port, RESULT(14) => 
                           A_neg_shifted_by1_5_14_port, RESULT(13) => 
                           A_neg_shifted_by1_5_13_port, RESULT(12) => 
                           A_neg_shifted_by1_5_12_port, RESULT(11) => 
                           A_neg_shifted_by1_5_11_port, RESULT(10) => 
                           A_neg_shifted_by1_5_10_port, RESULT(9) => 
                           A_neg_shifted_by1_5_9_port, RESULT(8) => 
                           A_neg_shifted_by1_5_8_port, RESULT(7) => 
                           A_neg_shifted_by1_5_7_port, RESULT(6) => 
                           A_neg_shifted_by1_5_6_port, RESULT(5) => 
                           A_neg_shifted_by1_5_5_port, RESULT(4) => 
                           A_neg_shifted_by1_5_4_port, RESULT(3) => 
                           A_neg_shifted_by1_5_3_port, RESULT(2) => 
                           A_neg_shifted_by1_5_2_port, RESULT(1) => 
                           A_neg_shifted_by1_5_1_port, RESULT(0) => n_1187);
   SHIFTERi_6_0 : Shifter_NBIT64_10 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_5_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_5_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_5_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_5_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_5_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_5_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_5_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_5_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_5_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_5_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_5_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_5_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_5_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_5_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_5_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_5_48_port, TO_SHIFT(47) => n203, 
                           TO_SHIFT(46) => A_neg_shifted_by2_5_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_5_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_5_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_5_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_5_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_5_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_5_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_5_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_5_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_5_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_5_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_5_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_5_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_5_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_5_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_5_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_5_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_5_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_5_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_5_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_5_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_5_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_5_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_5_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_5_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_5_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_5_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_5_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_5_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_5_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_5_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_5_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_5_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_5_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_5_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_5_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_5_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_5_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_5_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_5_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_5_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_5_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_5_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_5_3_port, 
                           TO_SHIFT(2) => A_neg_shifted_by2_5_2_port, 
                           TO_SHIFT(1) => A_neg_shifted_by2_5_1_port, 
                           TO_SHIFT(0) => A_neg_shifted_by2_5_0_port, 
                           RESULT(127) => A_neg_shifted_by2_6_63_port, 
                           RESULT(126) => A_neg_shifted_by2_6_62_port, 
                           RESULT(125) => A_neg_shifted_by2_6_61_port, 
                           RESULT(124) => A_neg_shifted_by2_6_60_port, 
                           RESULT(123) => A_neg_shifted_by2_6_59_port, 
                           RESULT(122) => A_neg_shifted_by2_6_58_port, 
                           RESULT(121) => A_neg_shifted_by2_6_57_port, 
                           RESULT(120) => A_neg_shifted_by2_6_56_port, 
                           RESULT(119) => A_neg_shifted_by2_6_55_port, 
                           RESULT(118) => A_neg_shifted_by2_6_54_port, 
                           RESULT(117) => A_neg_shifted_by2_6_53_port, 
                           RESULT(116) => A_neg_shifted_by2_6_52_port, 
                           RESULT(115) => A_neg_shifted_by2_6_51_port, 
                           RESULT(114) => A_neg_shifted_by2_6_50_port, 
                           RESULT(113) => A_neg_shifted_by2_6_49_port, 
                           RESULT(112) => A_neg_shifted_by2_6_48_port, 
                           RESULT(111) => A_neg_shifted_by2_6_47_port, 
                           RESULT(110) => A_neg_shifted_by2_6_46_port, 
                           RESULT(109) => A_neg_shifted_by2_6_45_port, 
                           RESULT(108) => A_neg_shifted_by2_6_44_port, 
                           RESULT(107) => A_neg_shifted_by2_6_43_port, 
                           RESULT(106) => A_neg_shifted_by2_6_42_port, 
                           RESULT(105) => A_neg_shifted_by2_6_41_port, 
                           RESULT(104) => A_neg_shifted_by2_6_40_port, 
                           RESULT(103) => A_neg_shifted_by2_6_39_port, 
                           RESULT(102) => A_neg_shifted_by2_6_38_port, 
                           RESULT(101) => A_neg_shifted_by2_6_37_port, 
                           RESULT(100) => A_neg_shifted_by2_6_36_port, 
                           RESULT(99) => A_neg_shifted_by2_6_35_port, 
                           RESULT(98) => A_neg_shifted_by2_6_34_port, 
                           RESULT(97) => A_neg_shifted_by2_6_33_port, 
                           RESULT(96) => A_neg_shifted_by2_6_32_port, 
                           RESULT(95) => A_neg_shifted_by2_6_31_port, 
                           RESULT(94) => A_neg_shifted_by2_6_30_port, 
                           RESULT(93) => A_neg_shifted_by2_6_29_port, 
                           RESULT(92) => A_neg_shifted_by2_6_28_port, 
                           RESULT(91) => A_neg_shifted_by2_6_27_port, 
                           RESULT(90) => A_neg_shifted_by2_6_26_port, 
                           RESULT(89) => A_neg_shifted_by2_6_25_port, 
                           RESULT(88) => A_neg_shifted_by2_6_24_port, 
                           RESULT(87) => A_neg_shifted_by2_6_23_port, 
                           RESULT(86) => A_neg_shifted_by2_6_22_port, 
                           RESULT(85) => A_neg_shifted_by2_6_21_port, 
                           RESULT(84) => A_neg_shifted_by2_6_20_port, 
                           RESULT(83) => A_neg_shifted_by2_6_19_port, 
                           RESULT(82) => A_neg_shifted_by2_6_18_port, 
                           RESULT(81) => A_neg_shifted_by2_6_17_port, 
                           RESULT(80) => A_neg_shifted_by2_6_16_port, 
                           RESULT(79) => A_neg_shifted_by2_6_15_port, 
                           RESULT(78) => A_neg_shifted_by2_6_14_port, 
                           RESULT(77) => A_neg_shifted_by2_6_13_port, 
                           RESULT(76) => A_neg_shifted_by2_6_12_port, 
                           RESULT(75) => A_neg_shifted_by2_6_11_port, 
                           RESULT(74) => A_neg_shifted_by2_6_10_port, 
                           RESULT(73) => A_neg_shifted_by2_6_9_port, RESULT(72)
                           => A_neg_shifted_by2_6_8_port, RESULT(71) => 
                           A_neg_shifted_by2_6_7_port, RESULT(70) => 
                           A_neg_shifted_by2_6_6_port, RESULT(69) => 
                           A_neg_shifted_by2_6_5_port, RESULT(68) => 
                           A_neg_shifted_by2_6_4_port, RESULT(67) => 
                           A_neg_shifted_by2_6_3_port, RESULT(66) => 
                           A_neg_shifted_by2_6_2_port, RESULT(65) => n_1188, 
                           RESULT(64) => n_1189, RESULT(63) => 
                           A_neg_shifted_by1_6_63_port, RESULT(62) => 
                           A_neg_shifted_by1_6_62_port, RESULT(61) => 
                           A_neg_shifted_by1_6_61_port, RESULT(60) => 
                           A_neg_shifted_by1_6_60_port, RESULT(59) => 
                           A_neg_shifted_by1_6_59_port, RESULT(58) => 
                           A_neg_shifted_by1_6_58_port, RESULT(57) => 
                           A_neg_shifted_by1_6_57_port, RESULT(56) => 
                           A_neg_shifted_by1_6_56_port, RESULT(55) => 
                           A_neg_shifted_by1_6_55_port, RESULT(54) => 
                           A_neg_shifted_by1_6_54_port, RESULT(53) => 
                           A_neg_shifted_by1_6_53_port, RESULT(52) => 
                           A_neg_shifted_by1_6_52_port, RESULT(51) => 
                           A_neg_shifted_by1_6_51_port, RESULT(50) => 
                           A_neg_shifted_by1_6_50_port, RESULT(49) => 
                           A_neg_shifted_by1_6_49_port, RESULT(48) => 
                           A_neg_shifted_by1_6_48_port, RESULT(47) => 
                           A_neg_shifted_by1_6_47_port, RESULT(46) => 
                           A_neg_shifted_by1_6_46_port, RESULT(45) => 
                           A_neg_shifted_by1_6_45_port, RESULT(44) => 
                           A_neg_shifted_by1_6_44_port, RESULT(43) => 
                           A_neg_shifted_by1_6_43_port, RESULT(42) => 
                           A_neg_shifted_by1_6_42_port, RESULT(41) => 
                           A_neg_shifted_by1_6_41_port, RESULT(40) => 
                           A_neg_shifted_by1_6_40_port, RESULT(39) => 
                           A_neg_shifted_by1_6_39_port, RESULT(38) => 
                           A_neg_shifted_by1_6_38_port, RESULT(37) => 
                           A_neg_shifted_by1_6_37_port, RESULT(36) => 
                           A_neg_shifted_by1_6_36_port, RESULT(35) => 
                           A_neg_shifted_by1_6_35_port, RESULT(34) => 
                           A_neg_shifted_by1_6_34_port, RESULT(33) => 
                           A_neg_shifted_by1_6_33_port, RESULT(32) => 
                           A_neg_shifted_by1_6_32_port, RESULT(31) => 
                           A_neg_shifted_by1_6_31_port, RESULT(30) => 
                           A_neg_shifted_by1_6_30_port, RESULT(29) => 
                           A_neg_shifted_by1_6_29_port, RESULT(28) => 
                           A_neg_shifted_by1_6_28_port, RESULT(27) => 
                           A_neg_shifted_by1_6_27_port, RESULT(26) => 
                           A_neg_shifted_by1_6_26_port, RESULT(25) => 
                           A_neg_shifted_by1_6_25_port, RESULT(24) => 
                           A_neg_shifted_by1_6_24_port, RESULT(23) => 
                           A_neg_shifted_by1_6_23_port, RESULT(22) => 
                           A_neg_shifted_by1_6_22_port, RESULT(21) => 
                           A_neg_shifted_by1_6_21_port, RESULT(20) => 
                           A_neg_shifted_by1_6_20_port, RESULT(19) => 
                           A_neg_shifted_by1_6_19_port, RESULT(18) => 
                           A_neg_shifted_by1_6_18_port, RESULT(17) => 
                           A_neg_shifted_by1_6_17_port, RESULT(16) => 
                           A_neg_shifted_by1_6_16_port, RESULT(15) => 
                           A_neg_shifted_by1_6_15_port, RESULT(14) => 
                           A_neg_shifted_by1_6_14_port, RESULT(13) => 
                           A_neg_shifted_by1_6_13_port, RESULT(12) => 
                           A_neg_shifted_by1_6_12_port, RESULT(11) => 
                           A_neg_shifted_by1_6_11_port, RESULT(10) => 
                           A_neg_shifted_by1_6_10_port, RESULT(9) => 
                           A_neg_shifted_by1_6_9_port, RESULT(8) => 
                           A_neg_shifted_by1_6_8_port, RESULT(7) => 
                           A_neg_shifted_by1_6_7_port, RESULT(6) => 
                           A_neg_shifted_by1_6_6_port, RESULT(5) => 
                           A_neg_shifted_by1_6_5_port, RESULT(4) => 
                           A_neg_shifted_by1_6_4_port, RESULT(3) => 
                           A_neg_shifted_by1_6_3_port, RESULT(2) => 
                           A_neg_shifted_by1_6_2_port, RESULT(1) => 
                           A_neg_shifted_by1_6_1_port, RESULT(0) => n_1190);
   SHIFTERi_7_0 : Shifter_NBIT64_9 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_6_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_6_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_6_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_6_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_6_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_6_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_6_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_6_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_6_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_6_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_6_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_6_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_6_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_6_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_6_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_6_48_port, TO_SHIFT(47) => n202, 
                           TO_SHIFT(46) => A_neg_shifted_by2_6_46_port, 
                           TO_SHIFT(45) => A_neg_shifted_by2_6_45_port, 
                           TO_SHIFT(44) => A_neg_shifted_by2_6_44_port, 
                           TO_SHIFT(43) => A_neg_shifted_by2_6_43_port, 
                           TO_SHIFT(42) => A_neg_shifted_by2_6_42_port, 
                           TO_SHIFT(41) => A_neg_shifted_by2_6_41_port, 
                           TO_SHIFT(40) => A_neg_shifted_by2_6_40_port, 
                           TO_SHIFT(39) => A_neg_shifted_by2_6_39_port, 
                           TO_SHIFT(38) => A_neg_shifted_by2_6_38_port, 
                           TO_SHIFT(37) => A_neg_shifted_by2_6_37_port, 
                           TO_SHIFT(36) => A_neg_shifted_by2_6_36_port, 
                           TO_SHIFT(35) => A_neg_shifted_by2_6_35_port, 
                           TO_SHIFT(34) => A_neg_shifted_by2_6_34_port, 
                           TO_SHIFT(33) => A_neg_shifted_by2_6_33_port, 
                           TO_SHIFT(32) => A_neg_shifted_by2_6_32_port, 
                           TO_SHIFT(31) => A_neg_shifted_by2_6_31_port, 
                           TO_SHIFT(30) => A_neg_shifted_by2_6_30_port, 
                           TO_SHIFT(29) => A_neg_shifted_by2_6_29_port, 
                           TO_SHIFT(28) => A_neg_shifted_by2_6_28_port, 
                           TO_SHIFT(27) => A_neg_shifted_by2_6_27_port, 
                           TO_SHIFT(26) => A_neg_shifted_by2_6_26_port, 
                           TO_SHIFT(25) => A_neg_shifted_by2_6_25_port, 
                           TO_SHIFT(24) => A_neg_shifted_by2_6_24_port, 
                           TO_SHIFT(23) => A_neg_shifted_by2_6_23_port, 
                           TO_SHIFT(22) => A_neg_shifted_by2_6_22_port, 
                           TO_SHIFT(21) => A_neg_shifted_by2_6_21_port, 
                           TO_SHIFT(20) => A_neg_shifted_by2_6_20_port, 
                           TO_SHIFT(19) => A_neg_shifted_by2_6_19_port, 
                           TO_SHIFT(18) => A_neg_shifted_by2_6_18_port, 
                           TO_SHIFT(17) => A_neg_shifted_by2_6_17_port, 
                           TO_SHIFT(16) => A_neg_shifted_by2_6_16_port, 
                           TO_SHIFT(15) => A_neg_shifted_by2_6_15_port, 
                           TO_SHIFT(14) => A_neg_shifted_by2_6_14_port, 
                           TO_SHIFT(13) => A_neg_shifted_by2_6_13_port, 
                           TO_SHIFT(12) => A_neg_shifted_by2_6_12_port, 
                           TO_SHIFT(11) => A_neg_shifted_by2_6_11_port, 
                           TO_SHIFT(10) => A_neg_shifted_by2_6_10_port, 
                           TO_SHIFT(9) => A_neg_shifted_by2_6_9_port, 
                           TO_SHIFT(8) => A_neg_shifted_by2_6_8_port, 
                           TO_SHIFT(7) => A_neg_shifted_by2_6_7_port, 
                           TO_SHIFT(6) => A_neg_shifted_by2_6_6_port, 
                           TO_SHIFT(5) => A_neg_shifted_by2_6_5_port, 
                           TO_SHIFT(4) => A_neg_shifted_by2_6_4_port, 
                           TO_SHIFT(3) => A_neg_shifted_by2_6_3_port, 
                           TO_SHIFT(2) => A_neg_shifted_by2_6_2_port, 
                           TO_SHIFT(1) => A_neg_shifted_by2_6_1_port, 
                           TO_SHIFT(0) => A_neg_shifted_by2_6_0_port, 
                           RESULT(127) => A_neg_shifted_by2_7_63_port, 
                           RESULT(126) => A_neg_shifted_by2_7_62_port, 
                           RESULT(125) => A_neg_shifted_by2_7_61_port, 
                           RESULT(124) => A_neg_shifted_by2_7_60_port, 
                           RESULT(123) => A_neg_shifted_by2_7_59_port, 
                           RESULT(122) => A_neg_shifted_by2_7_58_port, 
                           RESULT(121) => A_neg_shifted_by2_7_57_port, 
                           RESULT(120) => A_neg_shifted_by2_7_56_port, 
                           RESULT(119) => A_neg_shifted_by2_7_55_port, 
                           RESULT(118) => A_neg_shifted_by2_7_54_port, 
                           RESULT(117) => A_neg_shifted_by2_7_53_port, 
                           RESULT(116) => A_neg_shifted_by2_7_52_port, 
                           RESULT(115) => A_neg_shifted_by2_7_51_port, 
                           RESULT(114) => A_neg_shifted_by2_7_50_port, 
                           RESULT(113) => A_neg_shifted_by2_7_49_port, 
                           RESULT(112) => A_neg_shifted_by2_7_48_port, 
                           RESULT(111) => A_neg_shifted_by2_7_47_port, 
                           RESULT(110) => A_neg_shifted_by2_7_46_port, 
                           RESULT(109) => A_neg_shifted_by2_7_45_port, 
                           RESULT(108) => A_neg_shifted_by2_7_44_port, 
                           RESULT(107) => A_neg_shifted_by2_7_43_port, 
                           RESULT(106) => A_neg_shifted_by2_7_42_port, 
                           RESULT(105) => A_neg_shifted_by2_7_41_port, 
                           RESULT(104) => A_neg_shifted_by2_7_40_port, 
                           RESULT(103) => A_neg_shifted_by2_7_39_port, 
                           RESULT(102) => A_neg_shifted_by2_7_38_port, 
                           RESULT(101) => A_neg_shifted_by2_7_37_port, 
                           RESULT(100) => A_neg_shifted_by2_7_36_port, 
                           RESULT(99) => A_neg_shifted_by2_7_35_port, 
                           RESULT(98) => A_neg_shifted_by2_7_34_port, 
                           RESULT(97) => A_neg_shifted_by2_7_33_port, 
                           RESULT(96) => A_neg_shifted_by2_7_32_port, 
                           RESULT(95) => A_neg_shifted_by2_7_31_port, 
                           RESULT(94) => A_neg_shifted_by2_7_30_port, 
                           RESULT(93) => A_neg_shifted_by2_7_29_port, 
                           RESULT(92) => A_neg_shifted_by2_7_28_port, 
                           RESULT(91) => A_neg_shifted_by2_7_27_port, 
                           RESULT(90) => A_neg_shifted_by2_7_26_port, 
                           RESULT(89) => A_neg_shifted_by2_7_25_port, 
                           RESULT(88) => A_neg_shifted_by2_7_24_port, 
                           RESULT(87) => A_neg_shifted_by2_7_23_port, 
                           RESULT(86) => A_neg_shifted_by2_7_22_port, 
                           RESULT(85) => A_neg_shifted_by2_7_21_port, 
                           RESULT(84) => A_neg_shifted_by2_7_20_port, 
                           RESULT(83) => A_neg_shifted_by2_7_19_port, 
                           RESULT(82) => A_neg_shifted_by2_7_18_port, 
                           RESULT(81) => A_neg_shifted_by2_7_17_port, 
                           RESULT(80) => A_neg_shifted_by2_7_16_port, 
                           RESULT(79) => A_neg_shifted_by2_7_15_port, 
                           RESULT(78) => A_neg_shifted_by2_7_14_port, 
                           RESULT(77) => A_neg_shifted_by2_7_13_port, 
                           RESULT(76) => A_neg_shifted_by2_7_12_port, 
                           RESULT(75) => A_neg_shifted_by2_7_11_port, 
                           RESULT(74) => A_neg_shifted_by2_7_10_port, 
                           RESULT(73) => A_neg_shifted_by2_7_9_port, RESULT(72)
                           => A_neg_shifted_by2_7_8_port, RESULT(71) => 
                           A_neg_shifted_by2_7_7_port, RESULT(70) => 
                           A_neg_shifted_by2_7_6_port, RESULT(69) => 
                           A_neg_shifted_by2_7_5_port, RESULT(68) => 
                           A_neg_shifted_by2_7_4_port, RESULT(67) => 
                           A_neg_shifted_by2_7_3_port, RESULT(66) => 
                           A_neg_shifted_by2_7_2_port, RESULT(65) => n_1191, 
                           RESULT(64) => n_1192, RESULT(63) => 
                           A_neg_shifted_by1_7_63_port, RESULT(62) => 
                           A_neg_shifted_by1_7_62_port, RESULT(61) => 
                           A_neg_shifted_by1_7_61_port, RESULT(60) => 
                           A_neg_shifted_by1_7_60_port, RESULT(59) => 
                           A_neg_shifted_by1_7_59_port, RESULT(58) => 
                           A_neg_shifted_by1_7_58_port, RESULT(57) => 
                           A_neg_shifted_by1_7_57_port, RESULT(56) => 
                           A_neg_shifted_by1_7_56_port, RESULT(55) => 
                           A_neg_shifted_by1_7_55_port, RESULT(54) => 
                           A_neg_shifted_by1_7_54_port, RESULT(53) => 
                           A_neg_shifted_by1_7_53_port, RESULT(52) => 
                           A_neg_shifted_by1_7_52_port, RESULT(51) => 
                           A_neg_shifted_by1_7_51_port, RESULT(50) => 
                           A_neg_shifted_by1_7_50_port, RESULT(49) => 
                           A_neg_shifted_by1_7_49_port, RESULT(48) => 
                           A_neg_shifted_by1_7_48_port, RESULT(47) => 
                           A_neg_shifted_by1_7_47_port, RESULT(46) => 
                           A_neg_shifted_by1_7_46_port, RESULT(45) => 
                           A_neg_shifted_by1_7_45_port, RESULT(44) => 
                           A_neg_shifted_by1_7_44_port, RESULT(43) => 
                           A_neg_shifted_by1_7_43_port, RESULT(42) => 
                           A_neg_shifted_by1_7_42_port, RESULT(41) => 
                           A_neg_shifted_by1_7_41_port, RESULT(40) => 
                           A_neg_shifted_by1_7_40_port, RESULT(39) => 
                           A_neg_shifted_by1_7_39_port, RESULT(38) => 
                           A_neg_shifted_by1_7_38_port, RESULT(37) => 
                           A_neg_shifted_by1_7_37_port, RESULT(36) => 
                           A_neg_shifted_by1_7_36_port, RESULT(35) => 
                           A_neg_shifted_by1_7_35_port, RESULT(34) => 
                           A_neg_shifted_by1_7_34_port, RESULT(33) => 
                           A_neg_shifted_by1_7_33_port, RESULT(32) => 
                           A_neg_shifted_by1_7_32_port, RESULT(31) => 
                           A_neg_shifted_by1_7_31_port, RESULT(30) => 
                           A_neg_shifted_by1_7_30_port, RESULT(29) => 
                           A_neg_shifted_by1_7_29_port, RESULT(28) => 
                           A_neg_shifted_by1_7_28_port, RESULT(27) => 
                           A_neg_shifted_by1_7_27_port, RESULT(26) => 
                           A_neg_shifted_by1_7_26_port, RESULT(25) => 
                           A_neg_shifted_by1_7_25_port, RESULT(24) => 
                           A_neg_shifted_by1_7_24_port, RESULT(23) => 
                           A_neg_shifted_by1_7_23_port, RESULT(22) => 
                           A_neg_shifted_by1_7_22_port, RESULT(21) => 
                           A_neg_shifted_by1_7_21_port, RESULT(20) => 
                           A_neg_shifted_by1_7_20_port, RESULT(19) => 
                           A_neg_shifted_by1_7_19_port, RESULT(18) => 
                           A_neg_shifted_by1_7_18_port, RESULT(17) => 
                           A_neg_shifted_by1_7_17_port, RESULT(16) => 
                           A_neg_shifted_by1_7_16_port, RESULT(15) => 
                           A_neg_shifted_by1_7_15_port, RESULT(14) => 
                           A_neg_shifted_by1_7_14_port, RESULT(13) => 
                           A_neg_shifted_by1_7_13_port, RESULT(12) => 
                           A_neg_shifted_by1_7_12_port, RESULT(11) => 
                           A_neg_shifted_by1_7_11_port, RESULT(10) => 
                           A_neg_shifted_by1_7_10_port, RESULT(9) => 
                           A_neg_shifted_by1_7_9_port, RESULT(8) => 
                           A_neg_shifted_by1_7_8_port, RESULT(7) => 
                           A_neg_shifted_by1_7_7_port, RESULT(6) => 
                           A_neg_shifted_by1_7_6_port, RESULT(5) => 
                           A_neg_shifted_by1_7_5_port, RESULT(4) => 
                           A_neg_shifted_by1_7_4_port, RESULT(3) => 
                           A_neg_shifted_by1_7_3_port, RESULT(2) => 
                           A_neg_shifted_by1_7_2_port, RESULT(1) => 
                           A_neg_shifted_by1_7_1_port, RESULT(0) => n_1193);
   SHIFTERi_8_0 : Shifter_NBIT64_8 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_7_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_7_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_7_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_7_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_7_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_7_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_7_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_7_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_7_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_7_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_7_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_7_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_7_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_7_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_7_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_7_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_7_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_7_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_7_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_7_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_7_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_7_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_7_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_7_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_7_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_7_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_7_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_7_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_7_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_7_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_7_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_7_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_7_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_7_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_7_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_7_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_7_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_7_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_7_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_7_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_7_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_7_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_7_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_7_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_7_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_7_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_7_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_7_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_7_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_7_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_7_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_7_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_7_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_7_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_7_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_7_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_7_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_7_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_7_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_7_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_7_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_7_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_7_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_7_0_port, RESULT(127) => 
                           A_neg_shifted_by2_8_63_port, RESULT(126) => 
                           A_neg_shifted_by2_8_62_port, RESULT(125) => 
                           A_neg_shifted_by2_8_61_port, RESULT(124) => 
                           A_neg_shifted_by2_8_60_port, RESULT(123) => 
                           A_neg_shifted_by2_8_59_port, RESULT(122) => 
                           A_neg_shifted_by2_8_58_port, RESULT(121) => 
                           A_neg_shifted_by2_8_57_port, RESULT(120) => 
                           A_neg_shifted_by2_8_56_port, RESULT(119) => 
                           A_neg_shifted_by2_8_55_port, RESULT(118) => 
                           A_neg_shifted_by2_8_54_port, RESULT(117) => 
                           A_neg_shifted_by2_8_53_port, RESULT(116) => 
                           A_neg_shifted_by2_8_52_port, RESULT(115) => 
                           A_neg_shifted_by2_8_51_port, RESULT(114) => 
                           A_neg_shifted_by2_8_50_port, RESULT(113) => 
                           A_neg_shifted_by2_8_49_port, RESULT(112) => 
                           A_neg_shifted_by2_8_48_port, RESULT(111) => 
                           A_neg_shifted_by2_8_47_port, RESULT(110) => 
                           A_neg_shifted_by2_8_46_port, RESULT(109) => 
                           A_neg_shifted_by2_8_45_port, RESULT(108) => 
                           A_neg_shifted_by2_8_44_port, RESULT(107) => 
                           A_neg_shifted_by2_8_43_port, RESULT(106) => 
                           A_neg_shifted_by2_8_42_port, RESULT(105) => 
                           A_neg_shifted_by2_8_41_port, RESULT(104) => 
                           A_neg_shifted_by2_8_40_port, RESULT(103) => 
                           A_neg_shifted_by2_8_39_port, RESULT(102) => 
                           A_neg_shifted_by2_8_38_port, RESULT(101) => 
                           A_neg_shifted_by2_8_37_port, RESULT(100) => 
                           A_neg_shifted_by2_8_36_port, RESULT(99) => 
                           A_neg_shifted_by2_8_35_port, RESULT(98) => 
                           A_neg_shifted_by2_8_34_port, RESULT(97) => 
                           A_neg_shifted_by2_8_33_port, RESULT(96) => 
                           A_neg_shifted_by2_8_32_port, RESULT(95) => 
                           A_neg_shifted_by2_8_31_port, RESULT(94) => 
                           A_neg_shifted_by2_8_30_port, RESULT(93) => 
                           A_neg_shifted_by2_8_29_port, RESULT(92) => 
                           A_neg_shifted_by2_8_28_port, RESULT(91) => 
                           A_neg_shifted_by2_8_27_port, RESULT(90) => 
                           A_neg_shifted_by2_8_26_port, RESULT(89) => 
                           A_neg_shifted_by2_8_25_port, RESULT(88) => 
                           A_neg_shifted_by2_8_24_port, RESULT(87) => 
                           A_neg_shifted_by2_8_23_port, RESULT(86) => 
                           A_neg_shifted_by2_8_22_port, RESULT(85) => 
                           A_neg_shifted_by2_8_21_port, RESULT(84) => 
                           A_neg_shifted_by2_8_20_port, RESULT(83) => 
                           A_neg_shifted_by2_8_19_port, RESULT(82) => 
                           A_neg_shifted_by2_8_18_port, RESULT(81) => 
                           A_neg_shifted_by2_8_17_port, RESULT(80) => 
                           A_neg_shifted_by2_8_16_port, RESULT(79) => 
                           A_neg_shifted_by2_8_15_port, RESULT(78) => 
                           A_neg_shifted_by2_8_14_port, RESULT(77) => 
                           A_neg_shifted_by2_8_13_port, RESULT(76) => 
                           A_neg_shifted_by2_8_12_port, RESULT(75) => 
                           A_neg_shifted_by2_8_11_port, RESULT(74) => 
                           A_neg_shifted_by2_8_10_port, RESULT(73) => 
                           A_neg_shifted_by2_8_9_port, RESULT(72) => 
                           A_neg_shifted_by2_8_8_port, RESULT(71) => 
                           A_neg_shifted_by2_8_7_port, RESULT(70) => 
                           A_neg_shifted_by2_8_6_port, RESULT(69) => 
                           A_neg_shifted_by2_8_5_port, RESULT(68) => 
                           A_neg_shifted_by2_8_4_port, RESULT(67) => 
                           A_neg_shifted_by2_8_3_port, RESULT(66) => 
                           A_neg_shifted_by2_8_2_port, RESULT(65) => n_1194, 
                           RESULT(64) => n_1195, RESULT(63) => 
                           A_neg_shifted_by1_8_63_port, RESULT(62) => 
                           A_neg_shifted_by1_8_62_port, RESULT(61) => 
                           A_neg_shifted_by1_8_61_port, RESULT(60) => 
                           A_neg_shifted_by1_8_60_port, RESULT(59) => 
                           A_neg_shifted_by1_8_59_port, RESULT(58) => 
                           A_neg_shifted_by1_8_58_port, RESULT(57) => 
                           A_neg_shifted_by1_8_57_port, RESULT(56) => 
                           A_neg_shifted_by1_8_56_port, RESULT(55) => 
                           A_neg_shifted_by1_8_55_port, RESULT(54) => 
                           A_neg_shifted_by1_8_54_port, RESULT(53) => 
                           A_neg_shifted_by1_8_53_port, RESULT(52) => 
                           A_neg_shifted_by1_8_52_port, RESULT(51) => 
                           A_neg_shifted_by1_8_51_port, RESULT(50) => 
                           A_neg_shifted_by1_8_50_port, RESULT(49) => 
                           A_neg_shifted_by1_8_49_port, RESULT(48) => 
                           A_neg_shifted_by1_8_48_port, RESULT(47) => 
                           A_neg_shifted_by1_8_47_port, RESULT(46) => 
                           A_neg_shifted_by1_8_46_port, RESULT(45) => 
                           A_neg_shifted_by1_8_45_port, RESULT(44) => 
                           A_neg_shifted_by1_8_44_port, RESULT(43) => 
                           A_neg_shifted_by1_8_43_port, RESULT(42) => 
                           A_neg_shifted_by1_8_42_port, RESULT(41) => 
                           A_neg_shifted_by1_8_41_port, RESULT(40) => 
                           A_neg_shifted_by1_8_40_port, RESULT(39) => 
                           A_neg_shifted_by1_8_39_port, RESULT(38) => 
                           A_neg_shifted_by1_8_38_port, RESULT(37) => 
                           A_neg_shifted_by1_8_37_port, RESULT(36) => 
                           A_neg_shifted_by1_8_36_port, RESULT(35) => 
                           A_neg_shifted_by1_8_35_port, RESULT(34) => 
                           A_neg_shifted_by1_8_34_port, RESULT(33) => 
                           A_neg_shifted_by1_8_33_port, RESULT(32) => 
                           A_neg_shifted_by1_8_32_port, RESULT(31) => 
                           A_neg_shifted_by1_8_31_port, RESULT(30) => 
                           A_neg_shifted_by1_8_30_port, RESULT(29) => 
                           A_neg_shifted_by1_8_29_port, RESULT(28) => 
                           A_neg_shifted_by1_8_28_port, RESULT(27) => 
                           A_neg_shifted_by1_8_27_port, RESULT(26) => 
                           A_neg_shifted_by1_8_26_port, RESULT(25) => 
                           A_neg_shifted_by1_8_25_port, RESULT(24) => 
                           A_neg_shifted_by1_8_24_port, RESULT(23) => 
                           A_neg_shifted_by1_8_23_port, RESULT(22) => 
                           A_neg_shifted_by1_8_22_port, RESULT(21) => 
                           A_neg_shifted_by1_8_21_port, RESULT(20) => 
                           A_neg_shifted_by1_8_20_port, RESULT(19) => 
                           A_neg_shifted_by1_8_19_port, RESULT(18) => 
                           A_neg_shifted_by1_8_18_port, RESULT(17) => 
                           A_neg_shifted_by1_8_17_port, RESULT(16) => 
                           A_neg_shifted_by1_8_16_port, RESULT(15) => 
                           A_neg_shifted_by1_8_15_port, RESULT(14) => 
                           A_neg_shifted_by1_8_14_port, RESULT(13) => 
                           A_neg_shifted_by1_8_13_port, RESULT(12) => 
                           A_neg_shifted_by1_8_12_port, RESULT(11) => 
                           A_neg_shifted_by1_8_11_port, RESULT(10) => 
                           A_neg_shifted_by1_8_10_port, RESULT(9) => 
                           A_neg_shifted_by1_8_9_port, RESULT(8) => 
                           A_neg_shifted_by1_8_8_port, RESULT(7) => 
                           A_neg_shifted_by1_8_7_port, RESULT(6) => 
                           A_neg_shifted_by1_8_6_port, RESULT(5) => 
                           A_neg_shifted_by1_8_5_port, RESULT(4) => 
                           A_neg_shifted_by1_8_4_port, RESULT(3) => 
                           A_neg_shifted_by1_8_3_port, RESULT(2) => 
                           A_neg_shifted_by1_8_2_port, RESULT(1) => 
                           A_neg_shifted_by1_8_1_port, RESULT(0) => n_1196);
   SHIFTERi_9_0 : Shifter_NBIT64_7 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_8_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_8_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_8_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_8_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_8_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_8_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_8_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_8_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_8_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_8_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_8_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_8_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_8_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_8_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_8_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_8_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_8_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_8_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_8_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_8_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_8_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_8_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_8_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_8_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_8_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_8_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_8_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_8_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_8_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_8_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_8_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_8_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_8_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_8_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_8_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_8_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_8_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_8_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_8_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_8_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_8_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_8_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_8_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_8_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_8_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_8_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_8_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_8_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_8_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_8_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_8_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_8_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_8_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_8_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_8_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_8_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_8_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_8_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_8_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_8_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_8_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_8_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_8_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_8_0_port, RESULT(127) => 
                           A_neg_shifted_by2_9_63_port, RESULT(126) => 
                           A_neg_shifted_by2_9_62_port, RESULT(125) => 
                           A_neg_shifted_by2_9_61_port, RESULT(124) => 
                           A_neg_shifted_by2_9_60_port, RESULT(123) => 
                           A_neg_shifted_by2_9_59_port, RESULT(122) => 
                           A_neg_shifted_by2_9_58_port, RESULT(121) => 
                           A_neg_shifted_by2_9_57_port, RESULT(120) => 
                           A_neg_shifted_by2_9_56_port, RESULT(119) => 
                           A_neg_shifted_by2_9_55_port, RESULT(118) => 
                           A_neg_shifted_by2_9_54_port, RESULT(117) => 
                           A_neg_shifted_by2_9_53_port, RESULT(116) => 
                           A_neg_shifted_by2_9_52_port, RESULT(115) => 
                           A_neg_shifted_by2_9_51_port, RESULT(114) => 
                           A_neg_shifted_by2_9_50_port, RESULT(113) => 
                           A_neg_shifted_by2_9_49_port, RESULT(112) => 
                           A_neg_shifted_by2_9_48_port, RESULT(111) => 
                           A_neg_shifted_by2_9_47_port, RESULT(110) => 
                           A_neg_shifted_by2_9_46_port, RESULT(109) => 
                           A_neg_shifted_by2_9_45_port, RESULT(108) => 
                           A_neg_shifted_by2_9_44_port, RESULT(107) => 
                           A_neg_shifted_by2_9_43_port, RESULT(106) => 
                           A_neg_shifted_by2_9_42_port, RESULT(105) => 
                           A_neg_shifted_by2_9_41_port, RESULT(104) => 
                           A_neg_shifted_by2_9_40_port, RESULT(103) => 
                           A_neg_shifted_by2_9_39_port, RESULT(102) => 
                           A_neg_shifted_by2_9_38_port, RESULT(101) => 
                           A_neg_shifted_by2_9_37_port, RESULT(100) => 
                           A_neg_shifted_by2_9_36_port, RESULT(99) => 
                           A_neg_shifted_by2_9_35_port, RESULT(98) => 
                           A_neg_shifted_by2_9_34_port, RESULT(97) => 
                           A_neg_shifted_by2_9_33_port, RESULT(96) => 
                           A_neg_shifted_by2_9_32_port, RESULT(95) => 
                           A_neg_shifted_by2_9_31_port, RESULT(94) => 
                           A_neg_shifted_by2_9_30_port, RESULT(93) => 
                           A_neg_shifted_by2_9_29_port, RESULT(92) => 
                           A_neg_shifted_by2_9_28_port, RESULT(91) => 
                           A_neg_shifted_by2_9_27_port, RESULT(90) => 
                           A_neg_shifted_by2_9_26_port, RESULT(89) => 
                           A_neg_shifted_by2_9_25_port, RESULT(88) => 
                           A_neg_shifted_by2_9_24_port, RESULT(87) => 
                           A_neg_shifted_by2_9_23_port, RESULT(86) => 
                           A_neg_shifted_by2_9_22_port, RESULT(85) => 
                           A_neg_shifted_by2_9_21_port, RESULT(84) => 
                           A_neg_shifted_by2_9_20_port, RESULT(83) => 
                           A_neg_shifted_by2_9_19_port, RESULT(82) => 
                           A_neg_shifted_by2_9_18_port, RESULT(81) => 
                           A_neg_shifted_by2_9_17_port, RESULT(80) => 
                           A_neg_shifted_by2_9_16_port, RESULT(79) => 
                           A_neg_shifted_by2_9_15_port, RESULT(78) => 
                           A_neg_shifted_by2_9_14_port, RESULT(77) => 
                           A_neg_shifted_by2_9_13_port, RESULT(76) => 
                           A_neg_shifted_by2_9_12_port, RESULT(75) => 
                           A_neg_shifted_by2_9_11_port, RESULT(74) => 
                           A_neg_shifted_by2_9_10_port, RESULT(73) => 
                           A_neg_shifted_by2_9_9_port, RESULT(72) => 
                           A_neg_shifted_by2_9_8_port, RESULT(71) => 
                           A_neg_shifted_by2_9_7_port, RESULT(70) => 
                           A_neg_shifted_by2_9_6_port, RESULT(69) => 
                           A_neg_shifted_by2_9_5_port, RESULT(68) => 
                           A_neg_shifted_by2_9_4_port, RESULT(67) => 
                           A_neg_shifted_by2_9_3_port, RESULT(66) => 
                           A_neg_shifted_by2_9_2_port, RESULT(65) => n_1197, 
                           RESULT(64) => n_1198, RESULT(63) => 
                           A_neg_shifted_by1_9_63_port, RESULT(62) => 
                           A_neg_shifted_by1_9_62_port, RESULT(61) => 
                           A_neg_shifted_by1_9_61_port, RESULT(60) => 
                           A_neg_shifted_by1_9_60_port, RESULT(59) => 
                           A_neg_shifted_by1_9_59_port, RESULT(58) => 
                           A_neg_shifted_by1_9_58_port, RESULT(57) => 
                           A_neg_shifted_by1_9_57_port, RESULT(56) => 
                           A_neg_shifted_by1_9_56_port, RESULT(55) => 
                           A_neg_shifted_by1_9_55_port, RESULT(54) => 
                           A_neg_shifted_by1_9_54_port, RESULT(53) => 
                           A_neg_shifted_by1_9_53_port, RESULT(52) => 
                           A_neg_shifted_by1_9_52_port, RESULT(51) => 
                           A_neg_shifted_by1_9_51_port, RESULT(50) => 
                           A_neg_shifted_by1_9_50_port, RESULT(49) => 
                           A_neg_shifted_by1_9_49_port, RESULT(48) => 
                           A_neg_shifted_by1_9_48_port, RESULT(47) => 
                           A_neg_shifted_by1_9_47_port, RESULT(46) => 
                           A_neg_shifted_by1_9_46_port, RESULT(45) => 
                           A_neg_shifted_by1_9_45_port, RESULT(44) => 
                           A_neg_shifted_by1_9_44_port, RESULT(43) => 
                           A_neg_shifted_by1_9_43_port, RESULT(42) => 
                           A_neg_shifted_by1_9_42_port, RESULT(41) => 
                           A_neg_shifted_by1_9_41_port, RESULT(40) => 
                           A_neg_shifted_by1_9_40_port, RESULT(39) => 
                           A_neg_shifted_by1_9_39_port, RESULT(38) => 
                           A_neg_shifted_by1_9_38_port, RESULT(37) => 
                           A_neg_shifted_by1_9_37_port, RESULT(36) => 
                           A_neg_shifted_by1_9_36_port, RESULT(35) => 
                           A_neg_shifted_by1_9_35_port, RESULT(34) => 
                           A_neg_shifted_by1_9_34_port, RESULT(33) => 
                           A_neg_shifted_by1_9_33_port, RESULT(32) => 
                           A_neg_shifted_by1_9_32_port, RESULT(31) => 
                           A_neg_shifted_by1_9_31_port, RESULT(30) => 
                           A_neg_shifted_by1_9_30_port, RESULT(29) => 
                           A_neg_shifted_by1_9_29_port, RESULT(28) => 
                           A_neg_shifted_by1_9_28_port, RESULT(27) => 
                           A_neg_shifted_by1_9_27_port, RESULT(26) => 
                           A_neg_shifted_by1_9_26_port, RESULT(25) => 
                           A_neg_shifted_by1_9_25_port, RESULT(24) => 
                           A_neg_shifted_by1_9_24_port, RESULT(23) => 
                           A_neg_shifted_by1_9_23_port, RESULT(22) => 
                           A_neg_shifted_by1_9_22_port, RESULT(21) => 
                           A_neg_shifted_by1_9_21_port, RESULT(20) => 
                           A_neg_shifted_by1_9_20_port, RESULT(19) => 
                           A_neg_shifted_by1_9_19_port, RESULT(18) => 
                           A_neg_shifted_by1_9_18_port, RESULT(17) => 
                           A_neg_shifted_by1_9_17_port, RESULT(16) => 
                           A_neg_shifted_by1_9_16_port, RESULT(15) => 
                           A_neg_shifted_by1_9_15_port, RESULT(14) => 
                           A_neg_shifted_by1_9_14_port, RESULT(13) => 
                           A_neg_shifted_by1_9_13_port, RESULT(12) => 
                           A_neg_shifted_by1_9_12_port, RESULT(11) => 
                           A_neg_shifted_by1_9_11_port, RESULT(10) => 
                           A_neg_shifted_by1_9_10_port, RESULT(9) => 
                           A_neg_shifted_by1_9_9_port, RESULT(8) => 
                           A_neg_shifted_by1_9_8_port, RESULT(7) => 
                           A_neg_shifted_by1_9_7_port, RESULT(6) => 
                           A_neg_shifted_by1_9_6_port, RESULT(5) => 
                           A_neg_shifted_by1_9_5_port, RESULT(4) => 
                           A_neg_shifted_by1_9_4_port, RESULT(3) => 
                           A_neg_shifted_by1_9_3_port, RESULT(2) => 
                           A_neg_shifted_by1_9_2_port, RESULT(1) => 
                           A_neg_shifted_by1_9_1_port, RESULT(0) => n_1199);
   SHIFTERi_10_0 : Shifter_NBIT64_6 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_9_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_9_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_9_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_9_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_9_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_9_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_9_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_9_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_9_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_9_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_9_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_9_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_9_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_9_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_9_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_9_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_9_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_9_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_9_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_9_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_9_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_9_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_9_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_9_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_9_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_9_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_9_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_9_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_9_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_9_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_9_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_9_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_9_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_9_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_9_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_9_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_9_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_9_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_9_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_9_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_9_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_9_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_9_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_9_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_9_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_9_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_9_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_9_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_9_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_9_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_9_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_9_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_9_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_9_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_9_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_9_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_9_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_9_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_9_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_9_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_9_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_9_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_9_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_9_0_port, RESULT(127) => 
                           A_neg_shifted_by2_10_63_port, RESULT(126) => 
                           A_neg_shifted_by2_10_62_port, RESULT(125) => 
                           A_neg_shifted_by2_10_61_port, RESULT(124) => 
                           A_neg_shifted_by2_10_60_port, RESULT(123) => 
                           A_neg_shifted_by2_10_59_port, RESULT(122) => 
                           A_neg_shifted_by2_10_58_port, RESULT(121) => 
                           A_neg_shifted_by2_10_57_port, RESULT(120) => 
                           A_neg_shifted_by2_10_56_port, RESULT(119) => 
                           A_neg_shifted_by2_10_55_port, RESULT(118) => 
                           A_neg_shifted_by2_10_54_port, RESULT(117) => 
                           A_neg_shifted_by2_10_53_port, RESULT(116) => 
                           A_neg_shifted_by2_10_52_port, RESULT(115) => 
                           A_neg_shifted_by2_10_51_port, RESULT(114) => 
                           A_neg_shifted_by2_10_50_port, RESULT(113) => 
                           A_neg_shifted_by2_10_49_port, RESULT(112) => 
                           A_neg_shifted_by2_10_48_port, RESULT(111) => 
                           A_neg_shifted_by2_10_47_port, RESULT(110) => 
                           A_neg_shifted_by2_10_46_port, RESULT(109) => 
                           A_neg_shifted_by2_10_45_port, RESULT(108) => 
                           A_neg_shifted_by2_10_44_port, RESULT(107) => 
                           A_neg_shifted_by2_10_43_port, RESULT(106) => 
                           A_neg_shifted_by2_10_42_port, RESULT(105) => 
                           A_neg_shifted_by2_10_41_port, RESULT(104) => 
                           A_neg_shifted_by2_10_40_port, RESULT(103) => 
                           A_neg_shifted_by2_10_39_port, RESULT(102) => 
                           A_neg_shifted_by2_10_38_port, RESULT(101) => 
                           A_neg_shifted_by2_10_37_port, RESULT(100) => 
                           A_neg_shifted_by2_10_36_port, RESULT(99) => 
                           A_neg_shifted_by2_10_35_port, RESULT(98) => 
                           A_neg_shifted_by2_10_34_port, RESULT(97) => 
                           A_neg_shifted_by2_10_33_port, RESULT(96) => 
                           A_neg_shifted_by2_10_32_port, RESULT(95) => 
                           A_neg_shifted_by2_10_31_port, RESULT(94) => 
                           A_neg_shifted_by2_10_30_port, RESULT(93) => 
                           A_neg_shifted_by2_10_29_port, RESULT(92) => 
                           A_neg_shifted_by2_10_28_port, RESULT(91) => 
                           A_neg_shifted_by2_10_27_port, RESULT(90) => 
                           A_neg_shifted_by2_10_26_port, RESULT(89) => 
                           A_neg_shifted_by2_10_25_port, RESULT(88) => 
                           A_neg_shifted_by2_10_24_port, RESULT(87) => 
                           A_neg_shifted_by2_10_23_port, RESULT(86) => 
                           A_neg_shifted_by2_10_22_port, RESULT(85) => 
                           A_neg_shifted_by2_10_21_port, RESULT(84) => 
                           A_neg_shifted_by2_10_20_port, RESULT(83) => 
                           A_neg_shifted_by2_10_19_port, RESULT(82) => 
                           A_neg_shifted_by2_10_18_port, RESULT(81) => 
                           A_neg_shifted_by2_10_17_port, RESULT(80) => 
                           A_neg_shifted_by2_10_16_port, RESULT(79) => 
                           A_neg_shifted_by2_10_15_port, RESULT(78) => 
                           A_neg_shifted_by2_10_14_port, RESULT(77) => 
                           A_neg_shifted_by2_10_13_port, RESULT(76) => 
                           A_neg_shifted_by2_10_12_port, RESULT(75) => 
                           A_neg_shifted_by2_10_11_port, RESULT(74) => 
                           A_neg_shifted_by2_10_10_port, RESULT(73) => 
                           A_neg_shifted_by2_10_9_port, RESULT(72) => 
                           A_neg_shifted_by2_10_8_port, RESULT(71) => 
                           A_neg_shifted_by2_10_7_port, RESULT(70) => 
                           A_neg_shifted_by2_10_6_port, RESULT(69) => 
                           A_neg_shifted_by2_10_5_port, RESULT(68) => 
                           A_neg_shifted_by2_10_4_port, RESULT(67) => 
                           A_neg_shifted_by2_10_3_port, RESULT(66) => 
                           A_neg_shifted_by2_10_2_port, RESULT(65) => n_1200, 
                           RESULT(64) => n_1201, RESULT(63) => 
                           A_neg_shifted_by1_10_63_port, RESULT(62) => 
                           A_neg_shifted_by1_10_62_port, RESULT(61) => 
                           A_neg_shifted_by1_10_61_port, RESULT(60) => 
                           A_neg_shifted_by1_10_60_port, RESULT(59) => 
                           A_neg_shifted_by1_10_59_port, RESULT(58) => 
                           A_neg_shifted_by1_10_58_port, RESULT(57) => 
                           A_neg_shifted_by1_10_57_port, RESULT(56) => 
                           A_neg_shifted_by1_10_56_port, RESULT(55) => 
                           A_neg_shifted_by1_10_55_port, RESULT(54) => 
                           A_neg_shifted_by1_10_54_port, RESULT(53) => 
                           A_neg_shifted_by1_10_53_port, RESULT(52) => 
                           A_neg_shifted_by1_10_52_port, RESULT(51) => 
                           A_neg_shifted_by1_10_51_port, RESULT(50) => 
                           A_neg_shifted_by1_10_50_port, RESULT(49) => 
                           A_neg_shifted_by1_10_49_port, RESULT(48) => 
                           A_neg_shifted_by1_10_48_port, RESULT(47) => 
                           A_neg_shifted_by1_10_47_port, RESULT(46) => 
                           A_neg_shifted_by1_10_46_port, RESULT(45) => 
                           A_neg_shifted_by1_10_45_port, RESULT(44) => 
                           A_neg_shifted_by1_10_44_port, RESULT(43) => 
                           A_neg_shifted_by1_10_43_port, RESULT(42) => 
                           A_neg_shifted_by1_10_42_port, RESULT(41) => 
                           A_neg_shifted_by1_10_41_port, RESULT(40) => 
                           A_neg_shifted_by1_10_40_port, RESULT(39) => 
                           A_neg_shifted_by1_10_39_port, RESULT(38) => 
                           A_neg_shifted_by1_10_38_port, RESULT(37) => 
                           A_neg_shifted_by1_10_37_port, RESULT(36) => 
                           A_neg_shifted_by1_10_36_port, RESULT(35) => 
                           A_neg_shifted_by1_10_35_port, RESULT(34) => 
                           A_neg_shifted_by1_10_34_port, RESULT(33) => 
                           A_neg_shifted_by1_10_33_port, RESULT(32) => 
                           A_neg_shifted_by1_10_32_port, RESULT(31) => 
                           A_neg_shifted_by1_10_31_port, RESULT(30) => 
                           A_neg_shifted_by1_10_30_port, RESULT(29) => 
                           A_neg_shifted_by1_10_29_port, RESULT(28) => 
                           A_neg_shifted_by1_10_28_port, RESULT(27) => 
                           A_neg_shifted_by1_10_27_port, RESULT(26) => 
                           A_neg_shifted_by1_10_26_port, RESULT(25) => 
                           A_neg_shifted_by1_10_25_port, RESULT(24) => 
                           A_neg_shifted_by1_10_24_port, RESULT(23) => 
                           A_neg_shifted_by1_10_23_port, RESULT(22) => 
                           A_neg_shifted_by1_10_22_port, RESULT(21) => 
                           A_neg_shifted_by1_10_21_port, RESULT(20) => 
                           A_neg_shifted_by1_10_20_port, RESULT(19) => 
                           A_neg_shifted_by1_10_19_port, RESULT(18) => 
                           A_neg_shifted_by1_10_18_port, RESULT(17) => 
                           A_neg_shifted_by1_10_17_port, RESULT(16) => 
                           A_neg_shifted_by1_10_16_port, RESULT(15) => 
                           A_neg_shifted_by1_10_15_port, RESULT(14) => 
                           A_neg_shifted_by1_10_14_port, RESULT(13) => 
                           A_neg_shifted_by1_10_13_port, RESULT(12) => 
                           A_neg_shifted_by1_10_12_port, RESULT(11) => 
                           A_neg_shifted_by1_10_11_port, RESULT(10) => 
                           A_neg_shifted_by1_10_10_port, RESULT(9) => 
                           A_neg_shifted_by1_10_9_port, RESULT(8) => 
                           A_neg_shifted_by1_10_8_port, RESULT(7) => 
                           A_neg_shifted_by1_10_7_port, RESULT(6) => 
                           A_neg_shifted_by1_10_6_port, RESULT(5) => 
                           A_neg_shifted_by1_10_5_port, RESULT(4) => 
                           A_neg_shifted_by1_10_4_port, RESULT(3) => 
                           A_neg_shifted_by1_10_3_port, RESULT(2) => 
                           A_neg_shifted_by1_10_2_port, RESULT(1) => 
                           A_neg_shifted_by1_10_1_port, RESULT(0) => n_1202);
   SHIFTERi_11_0 : Shifter_NBIT64_5 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_10_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_10_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_10_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_10_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_10_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_10_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_10_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_10_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_10_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_10_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_10_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_10_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_10_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_10_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_10_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_10_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_10_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_10_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_10_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_10_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_10_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_10_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_10_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_10_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_10_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_10_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_10_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_10_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_10_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_10_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_10_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_10_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_10_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_10_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_10_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_10_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_10_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_10_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_10_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_10_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_10_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_10_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_10_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_10_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_10_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_10_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_10_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_10_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_10_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_10_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_10_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_10_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_10_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_10_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_10_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_10_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_10_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_10_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_10_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_10_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_10_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_10_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_10_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_10_0_port, RESULT(127) => 
                           A_neg_shifted_by2_11_63_port, RESULT(126) => 
                           A_neg_shifted_by2_11_62_port, RESULT(125) => 
                           A_neg_shifted_by2_11_61_port, RESULT(124) => 
                           A_neg_shifted_by2_11_60_port, RESULT(123) => 
                           A_neg_shifted_by2_11_59_port, RESULT(122) => 
                           A_neg_shifted_by2_11_58_port, RESULT(121) => 
                           A_neg_shifted_by2_11_57_port, RESULT(120) => 
                           A_neg_shifted_by2_11_56_port, RESULT(119) => 
                           A_neg_shifted_by2_11_55_port, RESULT(118) => 
                           A_neg_shifted_by2_11_54_port, RESULT(117) => 
                           A_neg_shifted_by2_11_53_port, RESULT(116) => 
                           A_neg_shifted_by2_11_52_port, RESULT(115) => 
                           A_neg_shifted_by2_11_51_port, RESULT(114) => 
                           A_neg_shifted_by2_11_50_port, RESULT(113) => 
                           A_neg_shifted_by2_11_49_port, RESULT(112) => 
                           A_neg_shifted_by2_11_48_port, RESULT(111) => 
                           A_neg_shifted_by2_11_47_port, RESULT(110) => 
                           A_neg_shifted_by2_11_46_port, RESULT(109) => 
                           A_neg_shifted_by2_11_45_port, RESULT(108) => 
                           A_neg_shifted_by2_11_44_port, RESULT(107) => 
                           A_neg_shifted_by2_11_43_port, RESULT(106) => 
                           A_neg_shifted_by2_11_42_port, RESULT(105) => 
                           A_neg_shifted_by2_11_41_port, RESULT(104) => 
                           A_neg_shifted_by2_11_40_port, RESULT(103) => 
                           A_neg_shifted_by2_11_39_port, RESULT(102) => 
                           A_neg_shifted_by2_11_38_port, RESULT(101) => 
                           A_neg_shifted_by2_11_37_port, RESULT(100) => 
                           A_neg_shifted_by2_11_36_port, RESULT(99) => 
                           A_neg_shifted_by2_11_35_port, RESULT(98) => 
                           A_neg_shifted_by2_11_34_port, RESULT(97) => 
                           A_neg_shifted_by2_11_33_port, RESULT(96) => 
                           A_neg_shifted_by2_11_32_port, RESULT(95) => 
                           A_neg_shifted_by2_11_31_port, RESULT(94) => 
                           A_neg_shifted_by2_11_30_port, RESULT(93) => 
                           A_neg_shifted_by2_11_29_port, RESULT(92) => 
                           A_neg_shifted_by2_11_28_port, RESULT(91) => 
                           A_neg_shifted_by2_11_27_port, RESULT(90) => 
                           A_neg_shifted_by2_11_26_port, RESULT(89) => 
                           A_neg_shifted_by2_11_25_port, RESULT(88) => 
                           A_neg_shifted_by2_11_24_port, RESULT(87) => 
                           A_neg_shifted_by2_11_23_port, RESULT(86) => 
                           A_neg_shifted_by2_11_22_port, RESULT(85) => 
                           A_neg_shifted_by2_11_21_port, RESULT(84) => 
                           A_neg_shifted_by2_11_20_port, RESULT(83) => 
                           A_neg_shifted_by2_11_19_port, RESULT(82) => 
                           A_neg_shifted_by2_11_18_port, RESULT(81) => 
                           A_neg_shifted_by2_11_17_port, RESULT(80) => 
                           A_neg_shifted_by2_11_16_port, RESULT(79) => 
                           A_neg_shifted_by2_11_15_port, RESULT(78) => 
                           A_neg_shifted_by2_11_14_port, RESULT(77) => 
                           A_neg_shifted_by2_11_13_port, RESULT(76) => 
                           A_neg_shifted_by2_11_12_port, RESULT(75) => 
                           A_neg_shifted_by2_11_11_port, RESULT(74) => 
                           A_neg_shifted_by2_11_10_port, RESULT(73) => 
                           A_neg_shifted_by2_11_9_port, RESULT(72) => 
                           A_neg_shifted_by2_11_8_port, RESULT(71) => 
                           A_neg_shifted_by2_11_7_port, RESULT(70) => 
                           A_neg_shifted_by2_11_6_port, RESULT(69) => 
                           A_neg_shifted_by2_11_5_port, RESULT(68) => 
                           A_neg_shifted_by2_11_4_port, RESULT(67) => 
                           A_neg_shifted_by2_11_3_port, RESULT(66) => 
                           A_neg_shifted_by2_11_2_port, RESULT(65) => n_1203, 
                           RESULT(64) => n_1204, RESULT(63) => 
                           A_neg_shifted_by1_11_63_port, RESULT(62) => 
                           A_neg_shifted_by1_11_62_port, RESULT(61) => 
                           A_neg_shifted_by1_11_61_port, RESULT(60) => 
                           A_neg_shifted_by1_11_60_port, RESULT(59) => 
                           A_neg_shifted_by1_11_59_port, RESULT(58) => 
                           A_neg_shifted_by1_11_58_port, RESULT(57) => 
                           A_neg_shifted_by1_11_57_port, RESULT(56) => 
                           A_neg_shifted_by1_11_56_port, RESULT(55) => 
                           A_neg_shifted_by1_11_55_port, RESULT(54) => 
                           A_neg_shifted_by1_11_54_port, RESULT(53) => 
                           A_neg_shifted_by1_11_53_port, RESULT(52) => 
                           A_neg_shifted_by1_11_52_port, RESULT(51) => 
                           A_neg_shifted_by1_11_51_port, RESULT(50) => 
                           A_neg_shifted_by1_11_50_port, RESULT(49) => 
                           A_neg_shifted_by1_11_49_port, RESULT(48) => 
                           A_neg_shifted_by1_11_48_port, RESULT(47) => 
                           A_neg_shifted_by1_11_47_port, RESULT(46) => 
                           A_neg_shifted_by1_11_46_port, RESULT(45) => 
                           A_neg_shifted_by1_11_45_port, RESULT(44) => 
                           A_neg_shifted_by1_11_44_port, RESULT(43) => 
                           A_neg_shifted_by1_11_43_port, RESULT(42) => 
                           A_neg_shifted_by1_11_42_port, RESULT(41) => 
                           A_neg_shifted_by1_11_41_port, RESULT(40) => 
                           A_neg_shifted_by1_11_40_port, RESULT(39) => 
                           A_neg_shifted_by1_11_39_port, RESULT(38) => 
                           A_neg_shifted_by1_11_38_port, RESULT(37) => 
                           A_neg_shifted_by1_11_37_port, RESULT(36) => 
                           A_neg_shifted_by1_11_36_port, RESULT(35) => 
                           A_neg_shifted_by1_11_35_port, RESULT(34) => 
                           A_neg_shifted_by1_11_34_port, RESULT(33) => 
                           A_neg_shifted_by1_11_33_port, RESULT(32) => 
                           A_neg_shifted_by1_11_32_port, RESULT(31) => 
                           A_neg_shifted_by1_11_31_port, RESULT(30) => 
                           A_neg_shifted_by1_11_30_port, RESULT(29) => 
                           A_neg_shifted_by1_11_29_port, RESULT(28) => 
                           A_neg_shifted_by1_11_28_port, RESULT(27) => 
                           A_neg_shifted_by1_11_27_port, RESULT(26) => 
                           A_neg_shifted_by1_11_26_port, RESULT(25) => 
                           A_neg_shifted_by1_11_25_port, RESULT(24) => 
                           A_neg_shifted_by1_11_24_port, RESULT(23) => 
                           A_neg_shifted_by1_11_23_port, RESULT(22) => 
                           A_neg_shifted_by1_11_22_port, RESULT(21) => 
                           A_neg_shifted_by1_11_21_port, RESULT(20) => 
                           A_neg_shifted_by1_11_20_port, RESULT(19) => 
                           A_neg_shifted_by1_11_19_port, RESULT(18) => 
                           A_neg_shifted_by1_11_18_port, RESULT(17) => 
                           A_neg_shifted_by1_11_17_port, RESULT(16) => 
                           A_neg_shifted_by1_11_16_port, RESULT(15) => 
                           A_neg_shifted_by1_11_15_port, RESULT(14) => 
                           A_neg_shifted_by1_11_14_port, RESULT(13) => 
                           A_neg_shifted_by1_11_13_port, RESULT(12) => 
                           A_neg_shifted_by1_11_12_port, RESULT(11) => 
                           A_neg_shifted_by1_11_11_port, RESULT(10) => 
                           A_neg_shifted_by1_11_10_port, RESULT(9) => 
                           A_neg_shifted_by1_11_9_port, RESULT(8) => 
                           A_neg_shifted_by1_11_8_port, RESULT(7) => 
                           A_neg_shifted_by1_11_7_port, RESULT(6) => 
                           A_neg_shifted_by1_11_6_port, RESULT(5) => 
                           A_neg_shifted_by1_11_5_port, RESULT(4) => 
                           A_neg_shifted_by1_11_4_port, RESULT(3) => 
                           A_neg_shifted_by1_11_3_port, RESULT(2) => 
                           A_neg_shifted_by1_11_2_port, RESULT(1) => 
                           A_neg_shifted_by1_11_1_port, RESULT(0) => n_1205);
   SHIFTERi_12_0 : Shifter_NBIT64_4 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_11_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_11_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_11_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_11_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_11_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_11_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_11_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_11_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_11_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_11_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_11_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_11_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_11_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_11_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_11_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_11_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_11_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_11_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_11_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_11_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_11_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_11_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_11_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_11_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_11_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_11_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_11_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_11_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_11_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_11_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_11_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_11_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_11_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_11_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_11_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_11_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_11_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_11_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_11_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_11_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_11_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_11_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_11_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_11_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_11_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_11_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_11_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_11_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_11_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_11_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_11_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_11_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_11_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_11_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_11_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_11_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_11_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_11_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_11_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_11_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_11_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_11_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_11_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_11_0_port, RESULT(127) => 
                           A_neg_shifted_by2_12_63_port, RESULT(126) => 
                           A_neg_shifted_by2_12_62_port, RESULT(125) => 
                           A_neg_shifted_by2_12_61_port, RESULT(124) => 
                           A_neg_shifted_by2_12_60_port, RESULT(123) => 
                           A_neg_shifted_by2_12_59_port, RESULT(122) => 
                           A_neg_shifted_by2_12_58_port, RESULT(121) => 
                           A_neg_shifted_by2_12_57_port, RESULT(120) => 
                           A_neg_shifted_by2_12_56_port, RESULT(119) => 
                           A_neg_shifted_by2_12_55_port, RESULT(118) => 
                           A_neg_shifted_by2_12_54_port, RESULT(117) => 
                           A_neg_shifted_by2_12_53_port, RESULT(116) => 
                           A_neg_shifted_by2_12_52_port, RESULT(115) => 
                           A_neg_shifted_by2_12_51_port, RESULT(114) => 
                           A_neg_shifted_by2_12_50_port, RESULT(113) => 
                           A_neg_shifted_by2_12_49_port, RESULT(112) => 
                           A_neg_shifted_by2_12_48_port, RESULT(111) => 
                           A_neg_shifted_by2_12_47_port, RESULT(110) => 
                           A_neg_shifted_by2_12_46_port, RESULT(109) => 
                           A_neg_shifted_by2_12_45_port, RESULT(108) => 
                           A_neg_shifted_by2_12_44_port, RESULT(107) => 
                           A_neg_shifted_by2_12_43_port, RESULT(106) => 
                           A_neg_shifted_by2_12_42_port, RESULT(105) => 
                           A_neg_shifted_by2_12_41_port, RESULT(104) => 
                           A_neg_shifted_by2_12_40_port, RESULT(103) => 
                           A_neg_shifted_by2_12_39_port, RESULT(102) => 
                           A_neg_shifted_by2_12_38_port, RESULT(101) => 
                           A_neg_shifted_by2_12_37_port, RESULT(100) => 
                           A_neg_shifted_by2_12_36_port, RESULT(99) => 
                           A_neg_shifted_by2_12_35_port, RESULT(98) => 
                           A_neg_shifted_by2_12_34_port, RESULT(97) => 
                           A_neg_shifted_by2_12_33_port, RESULT(96) => 
                           A_neg_shifted_by2_12_32_port, RESULT(95) => 
                           A_neg_shifted_by2_12_31_port, RESULT(94) => 
                           A_neg_shifted_by2_12_30_port, RESULT(93) => 
                           A_neg_shifted_by2_12_29_port, RESULT(92) => 
                           A_neg_shifted_by2_12_28_port, RESULT(91) => 
                           A_neg_shifted_by2_12_27_port, RESULT(90) => 
                           A_neg_shifted_by2_12_26_port, RESULT(89) => 
                           A_neg_shifted_by2_12_25_port, RESULT(88) => 
                           A_neg_shifted_by2_12_24_port, RESULT(87) => 
                           A_neg_shifted_by2_12_23_port, RESULT(86) => 
                           A_neg_shifted_by2_12_22_port, RESULT(85) => 
                           A_neg_shifted_by2_12_21_port, RESULT(84) => 
                           A_neg_shifted_by2_12_20_port, RESULT(83) => 
                           A_neg_shifted_by2_12_19_port, RESULT(82) => 
                           A_neg_shifted_by2_12_18_port, RESULT(81) => 
                           A_neg_shifted_by2_12_17_port, RESULT(80) => 
                           A_neg_shifted_by2_12_16_port, RESULT(79) => 
                           A_neg_shifted_by2_12_15_port, RESULT(78) => 
                           A_neg_shifted_by2_12_14_port, RESULT(77) => 
                           A_neg_shifted_by2_12_13_port, RESULT(76) => 
                           A_neg_shifted_by2_12_12_port, RESULT(75) => 
                           A_neg_shifted_by2_12_11_port, RESULT(74) => 
                           A_neg_shifted_by2_12_10_port, RESULT(73) => 
                           A_neg_shifted_by2_12_9_port, RESULT(72) => 
                           A_neg_shifted_by2_12_8_port, RESULT(71) => 
                           A_neg_shifted_by2_12_7_port, RESULT(70) => 
                           A_neg_shifted_by2_12_6_port, RESULT(69) => 
                           A_neg_shifted_by2_12_5_port, RESULT(68) => 
                           A_neg_shifted_by2_12_4_port, RESULT(67) => 
                           A_neg_shifted_by2_12_3_port, RESULT(66) => 
                           A_neg_shifted_by2_12_2_port, RESULT(65) => n_1206, 
                           RESULT(64) => n_1207, RESULT(63) => 
                           A_neg_shifted_by1_12_63_port, RESULT(62) => 
                           A_neg_shifted_by1_12_62_port, RESULT(61) => 
                           A_neg_shifted_by1_12_61_port, RESULT(60) => 
                           A_neg_shifted_by1_12_60_port, RESULT(59) => 
                           A_neg_shifted_by1_12_59_port, RESULT(58) => 
                           A_neg_shifted_by1_12_58_port, RESULT(57) => 
                           A_neg_shifted_by1_12_57_port, RESULT(56) => 
                           A_neg_shifted_by1_12_56_port, RESULT(55) => 
                           A_neg_shifted_by1_12_55_port, RESULT(54) => 
                           A_neg_shifted_by1_12_54_port, RESULT(53) => 
                           A_neg_shifted_by1_12_53_port, RESULT(52) => 
                           A_neg_shifted_by1_12_52_port, RESULT(51) => 
                           A_neg_shifted_by1_12_51_port, RESULT(50) => 
                           A_neg_shifted_by1_12_50_port, RESULT(49) => 
                           A_neg_shifted_by1_12_49_port, RESULT(48) => 
                           A_neg_shifted_by1_12_48_port, RESULT(47) => 
                           A_neg_shifted_by1_12_47_port, RESULT(46) => 
                           A_neg_shifted_by1_12_46_port, RESULT(45) => 
                           A_neg_shifted_by1_12_45_port, RESULT(44) => 
                           A_neg_shifted_by1_12_44_port, RESULT(43) => 
                           A_neg_shifted_by1_12_43_port, RESULT(42) => 
                           A_neg_shifted_by1_12_42_port, RESULT(41) => 
                           A_neg_shifted_by1_12_41_port, RESULT(40) => 
                           A_neg_shifted_by1_12_40_port, RESULT(39) => 
                           A_neg_shifted_by1_12_39_port, RESULT(38) => 
                           A_neg_shifted_by1_12_38_port, RESULT(37) => 
                           A_neg_shifted_by1_12_37_port, RESULT(36) => 
                           A_neg_shifted_by1_12_36_port, RESULT(35) => 
                           A_neg_shifted_by1_12_35_port, RESULT(34) => 
                           A_neg_shifted_by1_12_34_port, RESULT(33) => 
                           A_neg_shifted_by1_12_33_port, RESULT(32) => 
                           A_neg_shifted_by1_12_32_port, RESULT(31) => 
                           A_neg_shifted_by1_12_31_port, RESULT(30) => 
                           A_neg_shifted_by1_12_30_port, RESULT(29) => 
                           A_neg_shifted_by1_12_29_port, RESULT(28) => 
                           A_neg_shifted_by1_12_28_port, RESULT(27) => 
                           A_neg_shifted_by1_12_27_port, RESULT(26) => 
                           A_neg_shifted_by1_12_26_port, RESULT(25) => 
                           A_neg_shifted_by1_12_25_port, RESULT(24) => 
                           A_neg_shifted_by1_12_24_port, RESULT(23) => 
                           A_neg_shifted_by1_12_23_port, RESULT(22) => 
                           A_neg_shifted_by1_12_22_port, RESULT(21) => 
                           A_neg_shifted_by1_12_21_port, RESULT(20) => 
                           A_neg_shifted_by1_12_20_port, RESULT(19) => 
                           A_neg_shifted_by1_12_19_port, RESULT(18) => 
                           A_neg_shifted_by1_12_18_port, RESULT(17) => 
                           A_neg_shifted_by1_12_17_port, RESULT(16) => 
                           A_neg_shifted_by1_12_16_port, RESULT(15) => 
                           A_neg_shifted_by1_12_15_port, RESULT(14) => 
                           A_neg_shifted_by1_12_14_port, RESULT(13) => 
                           A_neg_shifted_by1_12_13_port, RESULT(12) => 
                           A_neg_shifted_by1_12_12_port, RESULT(11) => 
                           A_neg_shifted_by1_12_11_port, RESULT(10) => 
                           A_neg_shifted_by1_12_10_port, RESULT(9) => 
                           A_neg_shifted_by1_12_9_port, RESULT(8) => 
                           A_neg_shifted_by1_12_8_port, RESULT(7) => 
                           A_neg_shifted_by1_12_7_port, RESULT(6) => 
                           A_neg_shifted_by1_12_6_port, RESULT(5) => 
                           A_neg_shifted_by1_12_5_port, RESULT(4) => 
                           A_neg_shifted_by1_12_4_port, RESULT(3) => 
                           A_neg_shifted_by1_12_3_port, RESULT(2) => 
                           A_neg_shifted_by1_12_2_port, RESULT(1) => 
                           A_neg_shifted_by1_12_1_port, RESULT(0) => n_1208);
   SHIFTERi_13_0 : Shifter_NBIT64_3 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_12_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_12_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_12_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_12_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_12_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_12_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_12_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_12_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_12_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_12_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_12_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_12_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_12_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_12_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_12_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_12_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_12_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_12_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_12_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_12_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_12_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_12_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_12_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_12_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_12_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_12_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_12_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_12_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_12_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_12_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_12_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_12_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_12_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_12_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_12_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_12_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_12_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_12_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_12_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_12_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_12_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_12_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_12_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_12_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_12_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_12_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_12_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_12_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_12_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_12_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_12_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_12_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_12_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_12_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_12_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_12_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_12_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_12_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_12_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_12_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_12_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_12_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_12_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_12_0_port, RESULT(127) => 
                           A_neg_shifted_by2_13_63_port, RESULT(126) => 
                           A_neg_shifted_by2_13_62_port, RESULT(125) => 
                           A_neg_shifted_by2_13_61_port, RESULT(124) => 
                           A_neg_shifted_by2_13_60_port, RESULT(123) => 
                           A_neg_shifted_by2_13_59_port, RESULT(122) => 
                           A_neg_shifted_by2_13_58_port, RESULT(121) => 
                           A_neg_shifted_by2_13_57_port, RESULT(120) => 
                           A_neg_shifted_by2_13_56_port, RESULT(119) => 
                           A_neg_shifted_by2_13_55_port, RESULT(118) => 
                           A_neg_shifted_by2_13_54_port, RESULT(117) => 
                           A_neg_shifted_by2_13_53_port, RESULT(116) => 
                           A_neg_shifted_by2_13_52_port, RESULT(115) => 
                           A_neg_shifted_by2_13_51_port, RESULT(114) => 
                           A_neg_shifted_by2_13_50_port, RESULT(113) => 
                           A_neg_shifted_by2_13_49_port, RESULT(112) => 
                           A_neg_shifted_by2_13_48_port, RESULT(111) => 
                           A_neg_shifted_by2_13_47_port, RESULT(110) => 
                           A_neg_shifted_by2_13_46_port, RESULT(109) => 
                           A_neg_shifted_by2_13_45_port, RESULT(108) => 
                           A_neg_shifted_by2_13_44_port, RESULT(107) => 
                           A_neg_shifted_by2_13_43_port, RESULT(106) => 
                           A_neg_shifted_by2_13_42_port, RESULT(105) => 
                           A_neg_shifted_by2_13_41_port, RESULT(104) => 
                           A_neg_shifted_by2_13_40_port, RESULT(103) => 
                           A_neg_shifted_by2_13_39_port, RESULT(102) => 
                           A_neg_shifted_by2_13_38_port, RESULT(101) => 
                           A_neg_shifted_by2_13_37_port, RESULT(100) => 
                           A_neg_shifted_by2_13_36_port, RESULT(99) => 
                           A_neg_shifted_by2_13_35_port, RESULT(98) => 
                           A_neg_shifted_by2_13_34_port, RESULT(97) => 
                           A_neg_shifted_by2_13_33_port, RESULT(96) => 
                           A_neg_shifted_by2_13_32_port, RESULT(95) => 
                           A_neg_shifted_by2_13_31_port, RESULT(94) => 
                           A_neg_shifted_by2_13_30_port, RESULT(93) => 
                           A_neg_shifted_by2_13_29_port, RESULT(92) => 
                           A_neg_shifted_by2_13_28_port, RESULT(91) => 
                           A_neg_shifted_by2_13_27_port, RESULT(90) => 
                           A_neg_shifted_by2_13_26_port, RESULT(89) => 
                           A_neg_shifted_by2_13_25_port, RESULT(88) => 
                           A_neg_shifted_by2_13_24_port, RESULT(87) => 
                           A_neg_shifted_by2_13_23_port, RESULT(86) => 
                           A_neg_shifted_by2_13_22_port, RESULT(85) => 
                           A_neg_shifted_by2_13_21_port, RESULT(84) => 
                           A_neg_shifted_by2_13_20_port, RESULT(83) => 
                           A_neg_shifted_by2_13_19_port, RESULT(82) => 
                           A_neg_shifted_by2_13_18_port, RESULT(81) => 
                           A_neg_shifted_by2_13_17_port, RESULT(80) => 
                           A_neg_shifted_by2_13_16_port, RESULT(79) => 
                           A_neg_shifted_by2_13_15_port, RESULT(78) => 
                           A_neg_shifted_by2_13_14_port, RESULT(77) => 
                           A_neg_shifted_by2_13_13_port, RESULT(76) => 
                           A_neg_shifted_by2_13_12_port, RESULT(75) => 
                           A_neg_shifted_by2_13_11_port, RESULT(74) => 
                           A_neg_shifted_by2_13_10_port, RESULT(73) => 
                           A_neg_shifted_by2_13_9_port, RESULT(72) => 
                           A_neg_shifted_by2_13_8_port, RESULT(71) => 
                           A_neg_shifted_by2_13_7_port, RESULT(70) => 
                           A_neg_shifted_by2_13_6_port, RESULT(69) => 
                           A_neg_shifted_by2_13_5_port, RESULT(68) => 
                           A_neg_shifted_by2_13_4_port, RESULT(67) => 
                           A_neg_shifted_by2_13_3_port, RESULT(66) => 
                           A_neg_shifted_by2_13_2_port, RESULT(65) => n_1209, 
                           RESULT(64) => n_1210, RESULT(63) => 
                           A_neg_shifted_by1_13_63_port, RESULT(62) => 
                           A_neg_shifted_by1_13_62_port, RESULT(61) => 
                           A_neg_shifted_by1_13_61_port, RESULT(60) => 
                           A_neg_shifted_by1_13_60_port, RESULT(59) => 
                           A_neg_shifted_by1_13_59_port, RESULT(58) => 
                           A_neg_shifted_by1_13_58_port, RESULT(57) => 
                           A_neg_shifted_by1_13_57_port, RESULT(56) => 
                           A_neg_shifted_by1_13_56_port, RESULT(55) => 
                           A_neg_shifted_by1_13_55_port, RESULT(54) => 
                           A_neg_shifted_by1_13_54_port, RESULT(53) => 
                           A_neg_shifted_by1_13_53_port, RESULT(52) => 
                           A_neg_shifted_by1_13_52_port, RESULT(51) => 
                           A_neg_shifted_by1_13_51_port, RESULT(50) => 
                           A_neg_shifted_by1_13_50_port, RESULT(49) => 
                           A_neg_shifted_by1_13_49_port, RESULT(48) => 
                           A_neg_shifted_by1_13_48_port, RESULT(47) => 
                           A_neg_shifted_by1_13_47_port, RESULT(46) => 
                           A_neg_shifted_by1_13_46_port, RESULT(45) => 
                           A_neg_shifted_by1_13_45_port, RESULT(44) => 
                           A_neg_shifted_by1_13_44_port, RESULT(43) => 
                           A_neg_shifted_by1_13_43_port, RESULT(42) => 
                           A_neg_shifted_by1_13_42_port, RESULT(41) => 
                           A_neg_shifted_by1_13_41_port, RESULT(40) => 
                           A_neg_shifted_by1_13_40_port, RESULT(39) => 
                           A_neg_shifted_by1_13_39_port, RESULT(38) => 
                           A_neg_shifted_by1_13_38_port, RESULT(37) => 
                           A_neg_shifted_by1_13_37_port, RESULT(36) => 
                           A_neg_shifted_by1_13_36_port, RESULT(35) => 
                           A_neg_shifted_by1_13_35_port, RESULT(34) => 
                           A_neg_shifted_by1_13_34_port, RESULT(33) => 
                           A_neg_shifted_by1_13_33_port, RESULT(32) => 
                           A_neg_shifted_by1_13_32_port, RESULT(31) => 
                           A_neg_shifted_by1_13_31_port, RESULT(30) => 
                           A_neg_shifted_by1_13_30_port, RESULT(29) => 
                           A_neg_shifted_by1_13_29_port, RESULT(28) => 
                           A_neg_shifted_by1_13_28_port, RESULT(27) => 
                           A_neg_shifted_by1_13_27_port, RESULT(26) => 
                           A_neg_shifted_by1_13_26_port, RESULT(25) => 
                           A_neg_shifted_by1_13_25_port, RESULT(24) => 
                           A_neg_shifted_by1_13_24_port, RESULT(23) => 
                           A_neg_shifted_by1_13_23_port, RESULT(22) => 
                           A_neg_shifted_by1_13_22_port, RESULT(21) => 
                           A_neg_shifted_by1_13_21_port, RESULT(20) => 
                           A_neg_shifted_by1_13_20_port, RESULT(19) => 
                           A_neg_shifted_by1_13_19_port, RESULT(18) => 
                           A_neg_shifted_by1_13_18_port, RESULT(17) => 
                           A_neg_shifted_by1_13_17_port, RESULT(16) => 
                           A_neg_shifted_by1_13_16_port, RESULT(15) => 
                           A_neg_shifted_by1_13_15_port, RESULT(14) => 
                           A_neg_shifted_by1_13_14_port, RESULT(13) => 
                           A_neg_shifted_by1_13_13_port, RESULT(12) => 
                           A_neg_shifted_by1_13_12_port, RESULT(11) => 
                           A_neg_shifted_by1_13_11_port, RESULT(10) => 
                           A_neg_shifted_by1_13_10_port, RESULT(9) => 
                           A_neg_shifted_by1_13_9_port, RESULT(8) => 
                           A_neg_shifted_by1_13_8_port, RESULT(7) => 
                           A_neg_shifted_by1_13_7_port, RESULT(6) => 
                           A_neg_shifted_by1_13_6_port, RESULT(5) => 
                           A_neg_shifted_by1_13_5_port, RESULT(4) => 
                           A_neg_shifted_by1_13_4_port, RESULT(3) => 
                           A_neg_shifted_by1_13_3_port, RESULT(2) => 
                           A_neg_shifted_by1_13_2_port, RESULT(1) => 
                           A_neg_shifted_by1_13_1_port, RESULT(0) => n_1211);
   SHIFTERi_14_0 : Shifter_NBIT64_2 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_13_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_13_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_13_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_13_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_13_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_13_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_13_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_13_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_13_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_13_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_13_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_13_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_13_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_13_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_13_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_13_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_13_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_13_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_13_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_13_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_13_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_13_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_13_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_13_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_13_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_13_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_13_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_13_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_13_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_13_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_13_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_13_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_13_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_13_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_13_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_13_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_13_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_13_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_13_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_13_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_13_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_13_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_13_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_13_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_13_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_13_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_13_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_13_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_13_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_13_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_13_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_13_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_13_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_13_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_13_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_13_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_13_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_13_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_13_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_13_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_13_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_13_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_13_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_13_0_port, RESULT(127) => 
                           A_neg_shifted_by2_14_63_port, RESULT(126) => 
                           A_neg_shifted_by2_14_62_port, RESULT(125) => 
                           A_neg_shifted_by2_14_61_port, RESULT(124) => 
                           A_neg_shifted_by2_14_60_port, RESULT(123) => 
                           A_neg_shifted_by2_14_59_port, RESULT(122) => 
                           A_neg_shifted_by2_14_58_port, RESULT(121) => 
                           A_neg_shifted_by2_14_57_port, RESULT(120) => 
                           A_neg_shifted_by2_14_56_port, RESULT(119) => 
                           A_neg_shifted_by2_14_55_port, RESULT(118) => 
                           A_neg_shifted_by2_14_54_port, RESULT(117) => 
                           A_neg_shifted_by2_14_53_port, RESULT(116) => 
                           A_neg_shifted_by2_14_52_port, RESULT(115) => 
                           A_neg_shifted_by2_14_51_port, RESULT(114) => 
                           A_neg_shifted_by2_14_50_port, RESULT(113) => 
                           A_neg_shifted_by2_14_49_port, RESULT(112) => 
                           A_neg_shifted_by2_14_48_port, RESULT(111) => 
                           A_neg_shifted_by2_14_47_port, RESULT(110) => 
                           A_neg_shifted_by2_14_46_port, RESULT(109) => 
                           A_neg_shifted_by2_14_45_port, RESULT(108) => 
                           A_neg_shifted_by2_14_44_port, RESULT(107) => 
                           A_neg_shifted_by2_14_43_port, RESULT(106) => 
                           A_neg_shifted_by2_14_42_port, RESULT(105) => 
                           A_neg_shifted_by2_14_41_port, RESULT(104) => 
                           A_neg_shifted_by2_14_40_port, RESULT(103) => 
                           A_neg_shifted_by2_14_39_port, RESULT(102) => 
                           A_neg_shifted_by2_14_38_port, RESULT(101) => 
                           A_neg_shifted_by2_14_37_port, RESULT(100) => 
                           A_neg_shifted_by2_14_36_port, RESULT(99) => 
                           A_neg_shifted_by2_14_35_port, RESULT(98) => 
                           A_neg_shifted_by2_14_34_port, RESULT(97) => 
                           A_neg_shifted_by2_14_33_port, RESULT(96) => 
                           A_neg_shifted_by2_14_32_port, RESULT(95) => 
                           A_neg_shifted_by2_14_31_port, RESULT(94) => 
                           A_neg_shifted_by2_14_30_port, RESULT(93) => 
                           A_neg_shifted_by2_14_29_port, RESULT(92) => 
                           A_neg_shifted_by2_14_28_port, RESULT(91) => 
                           A_neg_shifted_by2_14_27_port, RESULT(90) => 
                           A_neg_shifted_by2_14_26_port, RESULT(89) => 
                           A_neg_shifted_by2_14_25_port, RESULT(88) => 
                           A_neg_shifted_by2_14_24_port, RESULT(87) => 
                           A_neg_shifted_by2_14_23_port, RESULT(86) => 
                           A_neg_shifted_by2_14_22_port, RESULT(85) => 
                           A_neg_shifted_by2_14_21_port, RESULT(84) => 
                           A_neg_shifted_by2_14_20_port, RESULT(83) => 
                           A_neg_shifted_by2_14_19_port, RESULT(82) => 
                           A_neg_shifted_by2_14_18_port, RESULT(81) => 
                           A_neg_shifted_by2_14_17_port, RESULT(80) => 
                           A_neg_shifted_by2_14_16_port, RESULT(79) => 
                           A_neg_shifted_by2_14_15_port, RESULT(78) => 
                           A_neg_shifted_by2_14_14_port, RESULT(77) => 
                           A_neg_shifted_by2_14_13_port, RESULT(76) => 
                           A_neg_shifted_by2_14_12_port, RESULT(75) => 
                           A_neg_shifted_by2_14_11_port, RESULT(74) => 
                           A_neg_shifted_by2_14_10_port, RESULT(73) => 
                           A_neg_shifted_by2_14_9_port, RESULT(72) => 
                           A_neg_shifted_by2_14_8_port, RESULT(71) => 
                           A_neg_shifted_by2_14_7_port, RESULT(70) => 
                           A_neg_shifted_by2_14_6_port, RESULT(69) => 
                           A_neg_shifted_by2_14_5_port, RESULT(68) => 
                           A_neg_shifted_by2_14_4_port, RESULT(67) => 
                           A_neg_shifted_by2_14_3_port, RESULT(66) => 
                           A_neg_shifted_by2_14_2_port, RESULT(65) => n_1212, 
                           RESULT(64) => n_1213, RESULT(63) => 
                           A_neg_shifted_by1_14_63_port, RESULT(62) => 
                           A_neg_shifted_by1_14_62_port, RESULT(61) => 
                           A_neg_shifted_by1_14_61_port, RESULT(60) => 
                           A_neg_shifted_by1_14_60_port, RESULT(59) => 
                           A_neg_shifted_by1_14_59_port, RESULT(58) => 
                           A_neg_shifted_by1_14_58_port, RESULT(57) => 
                           A_neg_shifted_by1_14_57_port, RESULT(56) => 
                           A_neg_shifted_by1_14_56_port, RESULT(55) => 
                           A_neg_shifted_by1_14_55_port, RESULT(54) => 
                           A_neg_shifted_by1_14_54_port, RESULT(53) => 
                           A_neg_shifted_by1_14_53_port, RESULT(52) => 
                           A_neg_shifted_by1_14_52_port, RESULT(51) => 
                           A_neg_shifted_by1_14_51_port, RESULT(50) => 
                           A_neg_shifted_by1_14_50_port, RESULT(49) => 
                           A_neg_shifted_by1_14_49_port, RESULT(48) => 
                           A_neg_shifted_by1_14_48_port, RESULT(47) => 
                           A_neg_shifted_by1_14_47_port, RESULT(46) => 
                           A_neg_shifted_by1_14_46_port, RESULT(45) => 
                           A_neg_shifted_by1_14_45_port, RESULT(44) => 
                           A_neg_shifted_by1_14_44_port, RESULT(43) => 
                           A_neg_shifted_by1_14_43_port, RESULT(42) => 
                           A_neg_shifted_by1_14_42_port, RESULT(41) => 
                           A_neg_shifted_by1_14_41_port, RESULT(40) => 
                           A_neg_shifted_by1_14_40_port, RESULT(39) => 
                           A_neg_shifted_by1_14_39_port, RESULT(38) => 
                           A_neg_shifted_by1_14_38_port, RESULT(37) => 
                           A_neg_shifted_by1_14_37_port, RESULT(36) => 
                           A_neg_shifted_by1_14_36_port, RESULT(35) => 
                           A_neg_shifted_by1_14_35_port, RESULT(34) => 
                           A_neg_shifted_by1_14_34_port, RESULT(33) => 
                           A_neg_shifted_by1_14_33_port, RESULT(32) => 
                           A_neg_shifted_by1_14_32_port, RESULT(31) => 
                           A_neg_shifted_by1_14_31_port, RESULT(30) => 
                           A_neg_shifted_by1_14_30_port, RESULT(29) => 
                           A_neg_shifted_by1_14_29_port, RESULT(28) => 
                           A_neg_shifted_by1_14_28_port, RESULT(27) => 
                           A_neg_shifted_by1_14_27_port, RESULT(26) => 
                           A_neg_shifted_by1_14_26_port, RESULT(25) => 
                           A_neg_shifted_by1_14_25_port, RESULT(24) => 
                           A_neg_shifted_by1_14_24_port, RESULT(23) => 
                           A_neg_shifted_by1_14_23_port, RESULT(22) => 
                           A_neg_shifted_by1_14_22_port, RESULT(21) => 
                           A_neg_shifted_by1_14_21_port, RESULT(20) => 
                           A_neg_shifted_by1_14_20_port, RESULT(19) => 
                           A_neg_shifted_by1_14_19_port, RESULT(18) => 
                           A_neg_shifted_by1_14_18_port, RESULT(17) => 
                           A_neg_shifted_by1_14_17_port, RESULT(16) => 
                           A_neg_shifted_by1_14_16_port, RESULT(15) => 
                           A_neg_shifted_by1_14_15_port, RESULT(14) => 
                           A_neg_shifted_by1_14_14_port, RESULT(13) => 
                           A_neg_shifted_by1_14_13_port, RESULT(12) => 
                           A_neg_shifted_by1_14_12_port, RESULT(11) => 
                           A_neg_shifted_by1_14_11_port, RESULT(10) => 
                           A_neg_shifted_by1_14_10_port, RESULT(9) => 
                           A_neg_shifted_by1_14_9_port, RESULT(8) => 
                           A_neg_shifted_by1_14_8_port, RESULT(7) => 
                           A_neg_shifted_by1_14_7_port, RESULT(6) => 
                           A_neg_shifted_by1_14_6_port, RESULT(5) => 
                           A_neg_shifted_by1_14_5_port, RESULT(4) => 
                           A_neg_shifted_by1_14_4_port, RESULT(3) => 
                           A_neg_shifted_by1_14_3_port, RESULT(2) => 
                           A_neg_shifted_by1_14_2_port, RESULT(1) => 
                           A_neg_shifted_by1_14_1_port, RESULT(0) => n_1214);
   SHIFTERi_15_0 : Shifter_NBIT64_1 port map( TO_SHIFT(63) => 
                           A_neg_shifted_by2_14_63_port, TO_SHIFT(62) => 
                           A_neg_shifted_by2_14_62_port, TO_SHIFT(61) => 
                           A_neg_shifted_by2_14_61_port, TO_SHIFT(60) => 
                           A_neg_shifted_by2_14_60_port, TO_SHIFT(59) => 
                           A_neg_shifted_by2_14_59_port, TO_SHIFT(58) => 
                           A_neg_shifted_by2_14_58_port, TO_SHIFT(57) => 
                           A_neg_shifted_by2_14_57_port, TO_SHIFT(56) => 
                           A_neg_shifted_by2_14_56_port, TO_SHIFT(55) => 
                           A_neg_shifted_by2_14_55_port, TO_SHIFT(54) => 
                           A_neg_shifted_by2_14_54_port, TO_SHIFT(53) => 
                           A_neg_shifted_by2_14_53_port, TO_SHIFT(52) => 
                           A_neg_shifted_by2_14_52_port, TO_SHIFT(51) => 
                           A_neg_shifted_by2_14_51_port, TO_SHIFT(50) => 
                           A_neg_shifted_by2_14_50_port, TO_SHIFT(49) => 
                           A_neg_shifted_by2_14_49_port, TO_SHIFT(48) => 
                           A_neg_shifted_by2_14_48_port, TO_SHIFT(47) => 
                           A_neg_shifted_by2_14_47_port, TO_SHIFT(46) => 
                           A_neg_shifted_by2_14_46_port, TO_SHIFT(45) => 
                           A_neg_shifted_by2_14_45_port, TO_SHIFT(44) => 
                           A_neg_shifted_by2_14_44_port, TO_SHIFT(43) => 
                           A_neg_shifted_by2_14_43_port, TO_SHIFT(42) => 
                           A_neg_shifted_by2_14_42_port, TO_SHIFT(41) => 
                           A_neg_shifted_by2_14_41_port, TO_SHIFT(40) => 
                           A_neg_shifted_by2_14_40_port, TO_SHIFT(39) => 
                           A_neg_shifted_by2_14_39_port, TO_SHIFT(38) => 
                           A_neg_shifted_by2_14_38_port, TO_SHIFT(37) => 
                           A_neg_shifted_by2_14_37_port, TO_SHIFT(36) => 
                           A_neg_shifted_by2_14_36_port, TO_SHIFT(35) => 
                           A_neg_shifted_by2_14_35_port, TO_SHIFT(34) => 
                           A_neg_shifted_by2_14_34_port, TO_SHIFT(33) => 
                           A_neg_shifted_by2_14_33_port, TO_SHIFT(32) => 
                           A_neg_shifted_by2_14_32_port, TO_SHIFT(31) => 
                           A_neg_shifted_by2_14_31_port, TO_SHIFT(30) => 
                           A_neg_shifted_by2_14_30_port, TO_SHIFT(29) => 
                           A_neg_shifted_by2_14_29_port, TO_SHIFT(28) => 
                           A_neg_shifted_by2_14_28_port, TO_SHIFT(27) => 
                           A_neg_shifted_by2_14_27_port, TO_SHIFT(26) => 
                           A_neg_shifted_by2_14_26_port, TO_SHIFT(25) => 
                           A_neg_shifted_by2_14_25_port, TO_SHIFT(24) => 
                           A_neg_shifted_by2_14_24_port, TO_SHIFT(23) => 
                           A_neg_shifted_by2_14_23_port, TO_SHIFT(22) => 
                           A_neg_shifted_by2_14_22_port, TO_SHIFT(21) => 
                           A_neg_shifted_by2_14_21_port, TO_SHIFT(20) => 
                           A_neg_shifted_by2_14_20_port, TO_SHIFT(19) => 
                           A_neg_shifted_by2_14_19_port, TO_SHIFT(18) => 
                           A_neg_shifted_by2_14_18_port, TO_SHIFT(17) => 
                           A_neg_shifted_by2_14_17_port, TO_SHIFT(16) => 
                           A_neg_shifted_by2_14_16_port, TO_SHIFT(15) => 
                           A_neg_shifted_by2_14_15_port, TO_SHIFT(14) => 
                           A_neg_shifted_by2_14_14_port, TO_SHIFT(13) => 
                           A_neg_shifted_by2_14_13_port, TO_SHIFT(12) => 
                           A_neg_shifted_by2_14_12_port, TO_SHIFT(11) => 
                           A_neg_shifted_by2_14_11_port, TO_SHIFT(10) => 
                           A_neg_shifted_by2_14_10_port, TO_SHIFT(9) => 
                           A_neg_shifted_by2_14_9_port, TO_SHIFT(8) => 
                           A_neg_shifted_by2_14_8_port, TO_SHIFT(7) => 
                           A_neg_shifted_by2_14_7_port, TO_SHIFT(6) => 
                           A_neg_shifted_by2_14_6_port, TO_SHIFT(5) => 
                           A_neg_shifted_by2_14_5_port, TO_SHIFT(4) => 
                           A_neg_shifted_by2_14_4_port, TO_SHIFT(3) => 
                           A_neg_shifted_by2_14_3_port, TO_SHIFT(2) => 
                           A_neg_shifted_by2_14_2_port, TO_SHIFT(1) => 
                           A_neg_shifted_by2_14_1_port, TO_SHIFT(0) => 
                           A_neg_shifted_by2_14_0_port, RESULT(127) => n_1215, 
                           RESULT(126) => n_1216, RESULT(125) => n_1217, 
                           RESULT(124) => n_1218, RESULT(123) => n_1219, 
                           RESULT(122) => n_1220, RESULT(121) => n_1221, 
                           RESULT(120) => n_1222, RESULT(119) => n_1223, 
                           RESULT(118) => n_1224, RESULT(117) => n_1225, 
                           RESULT(116) => n_1226, RESULT(115) => n_1227, 
                           RESULT(114) => n_1228, RESULT(113) => n_1229, 
                           RESULT(112) => n_1230, RESULT(111) => n_1231, 
                           RESULT(110) => n_1232, RESULT(109) => n_1233, 
                           RESULT(108) => n_1234, RESULT(107) => n_1235, 
                           RESULT(106) => n_1236, RESULT(105) => n_1237, 
                           RESULT(104) => n_1238, RESULT(103) => n_1239, 
                           RESULT(102) => n_1240, RESULT(101) => n_1241, 
                           RESULT(100) => n_1242, RESULT(99) => n_1243, 
                           RESULT(98) => n_1244, RESULT(97) => n_1245, 
                           RESULT(96) => n_1246, RESULT(95) => n_1247, 
                           RESULT(94) => n_1248, RESULT(93) => n_1249, 
                           RESULT(92) => n_1250, RESULT(91) => n_1251, 
                           RESULT(90) => n_1252, RESULT(89) => n_1253, 
                           RESULT(88) => n_1254, RESULT(87) => n_1255, 
                           RESULT(86) => n_1256, RESULT(85) => n_1257, 
                           RESULT(84) => n_1258, RESULT(83) => n_1259, 
                           RESULT(82) => n_1260, RESULT(81) => n_1261, 
                           RESULT(80) => n_1262, RESULT(79) => n_1263, 
                           RESULT(78) => n_1264, RESULT(77) => n_1265, 
                           RESULT(76) => n_1266, RESULT(75) => n_1267, 
                           RESULT(74) => n_1268, RESULT(73) => n_1269, 
                           RESULT(72) => n_1270, RESULT(71) => n_1271, 
                           RESULT(70) => n_1272, RESULT(69) => n_1273, 
                           RESULT(68) => n_1274, RESULT(67) => n_1275, 
                           RESULT(66) => n_1276, RESULT(65) => n_1277, 
                           RESULT(64) => n_1278, RESULT(63) => 
                           A_neg_shifted_by1_15_63_port, RESULT(62) => 
                           A_neg_shifted_by1_15_62_port, RESULT(61) => 
                           A_neg_shifted_by1_15_61_port, RESULT(60) => 
                           A_neg_shifted_by1_15_60_port, RESULT(59) => 
                           A_neg_shifted_by1_15_59_port, RESULT(58) => 
                           A_neg_shifted_by1_15_58_port, RESULT(57) => 
                           A_neg_shifted_by1_15_57_port, RESULT(56) => 
                           A_neg_shifted_by1_15_56_port, RESULT(55) => 
                           A_neg_shifted_by1_15_55_port, RESULT(54) => 
                           A_neg_shifted_by1_15_54_port, RESULT(53) => 
                           A_neg_shifted_by1_15_53_port, RESULT(52) => 
                           A_neg_shifted_by1_15_52_port, RESULT(51) => 
                           A_neg_shifted_by1_15_51_port, RESULT(50) => 
                           A_neg_shifted_by1_15_50_port, RESULT(49) => 
                           A_neg_shifted_by1_15_49_port, RESULT(48) => 
                           A_neg_shifted_by1_15_48_port, RESULT(47) => 
                           A_neg_shifted_by1_15_47_port, RESULT(46) => 
                           A_neg_shifted_by1_15_46_port, RESULT(45) => 
                           A_neg_shifted_by1_15_45_port, RESULT(44) => 
                           A_neg_shifted_by1_15_44_port, RESULT(43) => 
                           A_neg_shifted_by1_15_43_port, RESULT(42) => 
                           A_neg_shifted_by1_15_42_port, RESULT(41) => 
                           A_neg_shifted_by1_15_41_port, RESULT(40) => 
                           A_neg_shifted_by1_15_40_port, RESULT(39) => 
                           A_neg_shifted_by1_15_39_port, RESULT(38) => 
                           A_neg_shifted_by1_15_38_port, RESULT(37) => 
                           A_neg_shifted_by1_15_37_port, RESULT(36) => 
                           A_neg_shifted_by1_15_36_port, RESULT(35) => 
                           A_neg_shifted_by1_15_35_port, RESULT(34) => 
                           A_neg_shifted_by1_15_34_port, RESULT(33) => 
                           A_neg_shifted_by1_15_33_port, RESULT(32) => 
                           A_neg_shifted_by1_15_32_port, RESULT(31) => 
                           A_neg_shifted_by1_15_31_port, RESULT(30) => 
                           A_neg_shifted_by1_15_30_port, RESULT(29) => 
                           A_neg_shifted_by1_15_29_port, RESULT(28) => 
                           A_neg_shifted_by1_15_28_port, RESULT(27) => 
                           A_neg_shifted_by1_15_27_port, RESULT(26) => 
                           A_neg_shifted_by1_15_26_port, RESULT(25) => 
                           A_neg_shifted_by1_15_25_port, RESULT(24) => 
                           A_neg_shifted_by1_15_24_port, RESULT(23) => 
                           A_neg_shifted_by1_15_23_port, RESULT(22) => 
                           A_neg_shifted_by1_15_22_port, RESULT(21) => 
                           A_neg_shifted_by1_15_21_port, RESULT(20) => 
                           A_neg_shifted_by1_15_20_port, RESULT(19) => 
                           A_neg_shifted_by1_15_19_port, RESULT(18) => 
                           A_neg_shifted_by1_15_18_port, RESULT(17) => 
                           A_neg_shifted_by1_15_17_port, RESULT(16) => 
                           A_neg_shifted_by1_15_16_port, RESULT(15) => 
                           A_neg_shifted_by1_15_15_port, RESULT(14) => 
                           A_neg_shifted_by1_15_14_port, RESULT(13) => 
                           A_neg_shifted_by1_15_13_port, RESULT(12) => 
                           A_neg_shifted_by1_15_12_port, RESULT(11) => 
                           A_neg_shifted_by1_15_11_port, RESULT(10) => 
                           A_neg_shifted_by1_15_10_port, RESULT(9) => 
                           A_neg_shifted_by1_15_9_port, RESULT(8) => 
                           A_neg_shifted_by1_15_8_port, RESULT(7) => 
                           A_neg_shifted_by1_15_7_port, RESULT(6) => 
                           A_neg_shifted_by1_15_6_port, RESULT(5) => 
                           A_neg_shifted_by1_15_5_port, RESULT(4) => 
                           A_neg_shifted_by1_15_4_port, RESULT(3) => 
                           A_neg_shifted_by1_15_3_port, RESULT(2) => 
                           A_neg_shifted_by1_15_2_port, RESULT(1) => 
                           A_neg_shifted_by1_15_1_port, RESULT(0) => n_1279);
   MUX0_0 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_0 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => n233, INPUT(65) => n233, INPUT(66) => n233, 
                           INPUT(67) => n233, INPUT(68) => n233, INPUT(69) => 
                           n233, INPUT(70) => n233, INPUT(71) => n233, 
                           INPUT(72) => n233, INPUT(73) => n233, INPUT(74) => 
                           n233, INPUT(75) => n233, INPUT(76) => n233, 
                           INPUT(77) => n233, INPUT(78) => n233, INPUT(79) => 
                           n233, INPUT(80) => n233, INPUT(81) => n233, 
                           INPUT(82) => n233, INPUT(83) => n233, INPUT(84) => 
                           n233, INPUT(85) => n233, INPUT(86) => n233, 
                           INPUT(87) => n233, INPUT(88) => n233, INPUT(89) => 
                           n233, INPUT(90) => n233, INPUT(91) => n233, 
                           INPUT(92) => n233, INPUT(93) => n233, INPUT(94) => 
                           n233, INPUT(95) => n233, INPUT(96) => n233, 
                           INPUT(97) => n228, INPUT(98) => n226, INPUT(99) => 
                           n224, INPUT(100) => n222, INPUT(101) => n220, 
                           INPUT(102) => n218, INPUT(103) => n216, INPUT(104) 
                           => net15391, INPUT(105) => net15397, INPUT(106) => 
                           net15403, INPUT(107) => net15409, INPUT(108) => 
                           net15415, INPUT(109) => net15421, INPUT(110) => 
                           net15427, INPUT(111) => net15433, INPUT(112) => 
                           net15439, INPUT(113) => net15445, INPUT(114) => 
                           net15451, INPUT(115) => net15457, INPUT(116) => 
                           net15463, INPUT(117) => net15469, INPUT(118) => 
                           net15475, INPUT(119) => net15481, INPUT(120) => 
                           net15487, INPUT(121) => net15493, INPUT(122) => n214
                           , INPUT(123) => n212, INPUT(124) => n210, INPUT(125)
                           => n208, INPUT(126) => net15523, INPUT(127) => 
                           net15533, INPUT(128) => n200, INPUT(129) => n200, 
                           INPUT(130) => n200, INPUT(131) => n200, INPUT(132) 
                           => n200, INPUT(133) => n200, INPUT(134) => n200, 
                           INPUT(135) => n200, INPUT(136) => n200, INPUT(137) 
                           => n200, INPUT(138) => n200, INPUT(139) => n200, 
                           INPUT(140) => n200, INPUT(141) => n200, INPUT(142) 
                           => n200, INPUT(143) => n200, INPUT(144) => n200, 
                           INPUT(145) => n200, INPUT(146) => n200, INPUT(147) 
                           => n200, INPUT(148) => n200, INPUT(149) => n200, 
                           INPUT(150) => n200, INPUT(151) => n201, INPUT(152) 
                           => n201, INPUT(153) => n201, INPUT(154) => n201, 
                           INPUT(155) => n201, INPUT(156) => n201, INPUT(157) 
                           => n201, INPUT(158) => n201, INPUT(159) => n200, 
                           INPUT(160) => A_neg_tmp_31_port, INPUT(161) => 
                           A_neg_tmp_30_port, INPUT(162) => A_neg_tmp_29_port, 
                           INPUT(163) => A_neg_tmp_28_port, INPUT(164) => 
                           A_neg_tmp_27_port, INPUT(165) => A_neg_tmp_26_port, 
                           INPUT(166) => A_neg_tmp_25_port, INPUT(167) => 
                           A_neg_tmp_24_port, INPUT(168) => A_neg_tmp_23_port, 
                           INPUT(169) => A_neg_tmp_22_port, INPUT(170) => 
                           A_neg_tmp_21_port, INPUT(171) => A_neg_tmp_20_port, 
                           INPUT(172) => A_neg_tmp_19_port, INPUT(173) => 
                           A_neg_tmp_18_port, INPUT(174) => A_neg_tmp_17_port, 
                           INPUT(175) => A_neg_tmp_16_port, INPUT(176) => 
                           A_neg_tmp_15_port, INPUT(177) => A_neg_tmp_14_port, 
                           INPUT(178) => A_neg_tmp_13_port, INPUT(179) => 
                           A_neg_tmp_12_port, INPUT(180) => A_neg_tmp_11_port, 
                           INPUT(181) => A_neg_tmp_10_port, INPUT(182) => 
                           A_neg_tmp_9_port, INPUT(183) => A_neg_tmp_8_port, 
                           INPUT(184) => A_neg_tmp_7_port, INPUT(185) => 
                           A_neg_tmp_6_port, INPUT(186) => A_neg_tmp_5_port, 
                           INPUT(187) => A_neg_tmp_4_port, INPUT(188) => 
                           A_neg_tmp_3_port, INPUT(189) => A_neg_tmp_2_port, 
                           INPUT(190) => n142, INPUT(191) => A_neg_tmp_0_port, 
                           INPUT(192) => A_pos_shifted_by1_0_63_port, 
                           INPUT(193) => A_pos_shifted_by1_0_62_port, 
                           INPUT(194) => A_pos_shifted_by1_0_61_port, 
                           INPUT(195) => A_pos_shifted_by1_0_60_port, 
                           INPUT(196) => A_pos_shifted_by1_0_59_port, 
                           INPUT(197) => A_pos_shifted_by1_0_58_port, 
                           INPUT(198) => A_pos_shifted_by1_0_57_port, 
                           INPUT(199) => A_pos_shifted_by1_0_56_port, 
                           INPUT(200) => A_pos_shifted_by1_0_55_port, 
                           INPUT(201) => A_pos_shifted_by1_0_54_port, 
                           INPUT(202) => A_pos_shifted_by1_0_53_port, 
                           INPUT(203) => A_pos_shifted_by1_0_52_port, 
                           INPUT(204) => A_pos_shifted_by1_0_51_port, 
                           INPUT(205) => A_pos_shifted_by1_0_50_port, 
                           INPUT(206) => A_pos_shifted_by1_0_49_port, 
                           INPUT(207) => A_pos_shifted_by1_0_48_port, 
                           INPUT(208) => A_pos_shifted_by1_0_47_port, 
                           INPUT(209) => A_pos_shifted_by1_0_46_port, 
                           INPUT(210) => A_pos_shifted_by1_0_45_port, 
                           INPUT(211) => A_pos_shifted_by1_0_44_port, 
                           INPUT(212) => A_pos_shifted_by1_0_43_port, 
                           INPUT(213) => A_pos_shifted_by1_0_42_port, 
                           INPUT(214) => A_pos_shifted_by1_0_41_port, 
                           INPUT(215) => A_pos_shifted_by1_0_40_port, 
                           INPUT(216) => A_pos_shifted_by1_0_39_port, 
                           INPUT(217) => A_pos_shifted_by1_0_38_port, 
                           INPUT(218) => A_pos_shifted_by1_0_37_port, 
                           INPUT(219) => A_pos_shifted_by1_0_36_port, 
                           INPUT(220) => A_pos_shifted_by1_0_35_port, 
                           INPUT(221) => A_pos_shifted_by1_0_34_port, 
                           INPUT(222) => A_pos_shifted_by1_0_33_port, 
                           INPUT(223) => A_pos_shifted_by1_0_32_port, 
                           INPUT(224) => A_pos_shifted_by1_0_31_port, 
                           INPUT(225) => A_pos_shifted_by1_0_30_port, 
                           INPUT(226) => A_pos_shifted_by1_0_29_port, 
                           INPUT(227) => A_pos_shifted_by1_0_28_port, 
                           INPUT(228) => A_pos_shifted_by1_0_27_port, 
                           INPUT(229) => A_pos_shifted_by1_0_26_port, 
                           INPUT(230) => A_pos_shifted_by1_0_25_port, 
                           INPUT(231) => A_pos_shifted_by1_0_24_port, 
                           INPUT(232) => A_pos_shifted_by1_0_23_port, 
                           INPUT(233) => A_pos_shifted_by1_0_22_port, 
                           INPUT(234) => A_pos_shifted_by1_0_21_port, 
                           INPUT(235) => A_pos_shifted_by1_0_20_port, 
                           INPUT(236) => A_pos_shifted_by1_0_19_port, 
                           INPUT(237) => A_pos_shifted_by1_0_18_port, 
                           INPUT(238) => A_pos_shifted_by1_0_17_port, 
                           INPUT(239) => A_pos_shifted_by1_0_16_port, 
                           INPUT(240) => A_pos_shifted_by1_0_15_port, 
                           INPUT(241) => A_pos_shifted_by1_0_14_port, 
                           INPUT(242) => A_pos_shifted_by1_0_13_port, 
                           INPUT(243) => A_pos_shifted_by1_0_12_port, 
                           INPUT(244) => A_pos_shifted_by1_0_11_port, 
                           INPUT(245) => A_pos_shifted_by1_0_10_port, 
                           INPUT(246) => A_pos_shifted_by1_0_9_port, INPUT(247)
                           => A_pos_shifted_by1_0_8_port, INPUT(248) => 
                           A_pos_shifted_by1_0_7_port, INPUT(249) => 
                           A_pos_shifted_by1_0_6_port, INPUT(250) => 
                           A_pos_shifted_by1_0_5_port, INPUT(251) => 
                           A_pos_shifted_by1_0_4_port, INPUT(252) => 
                           A_pos_shifted_by1_0_3_port, INPUT(253) => 
                           A_pos_shifted_by1_0_2_port, INPUT(254) => 
                           A_pos_shifted_by1_0_1_port, INPUT(255) => 
                           A_pos_shifted_by1_0_0_port, INPUT(256) => 
                           A_neg_shifted_by1_0_63_port, INPUT(257) => 
                           A_neg_shifted_by1_0_62_port, INPUT(258) => 
                           A_neg_shifted_by1_0_61_port, INPUT(259) => 
                           A_neg_shifted_by1_0_60_port, INPUT(260) => 
                           A_neg_shifted_by1_0_59_port, INPUT(261) => 
                           A_neg_shifted_by1_0_58_port, INPUT(262) => 
                           A_neg_shifted_by1_0_57_port, INPUT(263) => 
                           A_neg_shifted_by1_0_56_port, INPUT(264) => 
                           A_neg_shifted_by1_0_55_port, INPUT(265) => 
                           A_neg_shifted_by1_0_54_port, INPUT(266) => 
                           A_neg_shifted_by1_0_53_port, INPUT(267) => 
                           A_neg_shifted_by1_0_52_port, INPUT(268) => 
                           A_neg_shifted_by1_0_51_port, INPUT(269) => 
                           A_neg_shifted_by1_0_50_port, INPUT(270) => 
                           A_neg_shifted_by1_0_49_port, INPUT(271) => 
                           A_neg_shifted_by1_0_48_port, INPUT(272) => 
                           A_neg_shifted_by1_0_47_port, INPUT(273) => 
                           A_neg_shifted_by1_0_46_port, INPUT(274) => 
                           A_neg_shifted_by1_0_45_port, INPUT(275) => 
                           A_neg_shifted_by1_0_44_port, INPUT(276) => 
                           A_neg_shifted_by1_0_43_port, INPUT(277) => 
                           A_neg_shifted_by1_0_42_port, INPUT(278) => 
                           A_neg_shifted_by1_0_41_port, INPUT(279) => 
                           A_neg_shifted_by1_0_40_port, INPUT(280) => 
                           A_neg_shifted_by1_0_39_port, INPUT(281) => 
                           A_neg_shifted_by1_0_38_port, INPUT(282) => 
                           A_neg_shifted_by1_0_37_port, INPUT(283) => 
                           A_neg_shifted_by1_0_36_port, INPUT(284) => 
                           A_neg_shifted_by1_0_35_port, INPUT(285) => 
                           A_neg_shifted_by1_0_34_port, INPUT(286) => 
                           A_neg_shifted_by1_0_33_port, INPUT(287) => 
                           A_neg_shifted_by1_0_32_port, INPUT(288) => 
                           A_neg_shifted_by1_0_31_port, INPUT(289) => 
                           A_neg_shifted_by1_0_30_port, INPUT(290) => 
                           A_neg_shifted_by1_0_29_port, INPUT(291) => 
                           A_neg_shifted_by1_0_28_port, INPUT(292) => 
                           A_neg_shifted_by1_0_27_port, INPUT(293) => 
                           A_neg_shifted_by1_0_26_port, INPUT(294) => 
                           A_neg_shifted_by1_0_25_port, INPUT(295) => 
                           A_neg_shifted_by1_0_24_port, INPUT(296) => 
                           A_neg_shifted_by1_0_23_port, INPUT(297) => 
                           A_neg_shifted_by1_0_22_port, INPUT(298) => 
                           A_neg_shifted_by1_0_21_port, INPUT(299) => 
                           A_neg_shifted_by1_0_20_port, INPUT(300) => 
                           A_neg_shifted_by1_0_19_port, INPUT(301) => 
                           A_neg_shifted_by1_0_18_port, INPUT(302) => 
                           A_neg_shifted_by1_0_17_port, INPUT(303) => 
                           A_neg_shifted_by1_0_16_port, INPUT(304) => 
                           A_neg_shifted_by1_0_15_port, INPUT(305) => 
                           A_neg_shifted_by1_0_14_port, INPUT(306) => 
                           A_neg_shifted_by1_0_13_port, INPUT(307) => 
                           A_neg_shifted_by1_0_12_port, INPUT(308) => 
                           A_neg_shifted_by1_0_11_port, INPUT(309) => 
                           A_neg_shifted_by1_0_10_port, INPUT(310) => 
                           A_neg_shifted_by1_0_9_port, INPUT(311) => 
                           A_neg_shifted_by1_0_8_port, INPUT(312) => 
                           A_neg_shifted_by1_0_7_port, INPUT(313) => 
                           A_neg_shifted_by1_0_6_port, INPUT(314) => 
                           A_neg_shifted_by1_0_5_port, INPUT(315) => 
                           A_neg_shifted_by1_0_4_port, INPUT(316) => 
                           A_neg_shifted_by1_0_3_port, INPUT(317) => 
                           A_neg_shifted_by1_0_2_port, INPUT(318) => 
                           A_neg_shifted_by1_0_1_port, INPUT(319) => 
                           A_neg_shifted_by1_0_0_port, SEL(0) => 
                           selection_signal_0_2_port, SEL(1) => 
                           selection_signal_0_1_port, SEL(2) => 
                           selection_signal_0_0_port, Y(0) => P_tmp_0_63_port, 
                           Y(1) => P_tmp_0_62_port, Y(2) => P_tmp_0_61_port, 
                           Y(3) => P_tmp_0_60_port, Y(4) => P_tmp_0_59_port, 
                           Y(5) => P_tmp_0_58_port, Y(6) => P_tmp_0_57_port, 
                           Y(7) => P_tmp_0_56_port, Y(8) => P_tmp_0_55_port, 
                           Y(9) => P_tmp_0_54_port, Y(10) => P_tmp_0_53_port, 
                           Y(11) => P_tmp_0_52_port, Y(12) => P_tmp_0_51_port, 
                           Y(13) => P_tmp_0_50_port, Y(14) => P_tmp_0_49_port, 
                           Y(15) => P_tmp_0_48_port, Y(16) => P_tmp_0_47_port, 
                           Y(17) => P_tmp_0_46_port, Y(18) => P_tmp_0_45_port, 
                           Y(19) => P_tmp_0_44_port, Y(20) => P_tmp_0_43_port, 
                           Y(21) => P_tmp_0_42_port, Y(22) => P_tmp_0_41_port, 
                           Y(23) => P_tmp_0_40_port, Y(24) => P_tmp_0_39_port, 
                           Y(25) => P_tmp_0_38_port, Y(26) => P_tmp_0_37_port, 
                           Y(27) => P_tmp_0_36_port, Y(28) => P_tmp_0_35_port, 
                           Y(29) => P_tmp_0_34_port, Y(30) => P_tmp_0_33_port, 
                           Y(31) => P_tmp_0_32_port, Y(32) => P_tmp_0_31_port, 
                           Y(33) => P_tmp_0_30_port, Y(34) => P_tmp_0_29_port, 
                           Y(35) => P_tmp_0_28_port, Y(36) => P_tmp_0_27_port, 
                           Y(37) => P_tmp_0_26_port, Y(38) => P_tmp_0_25_port, 
                           Y(39) => P_tmp_0_24_port, Y(40) => P_tmp_0_23_port, 
                           Y(41) => P_tmp_0_22_port, Y(42) => P_tmp_0_21_port, 
                           Y(43) => P_tmp_0_20_port, Y(44) => P_tmp_0_19_port, 
                           Y(45) => P_tmp_0_18_port, Y(46) => P_tmp_0_17_port, 
                           Y(47) => P_tmp_0_16_port, Y(48) => P_tmp_0_15_port, 
                           Y(49) => P_tmp_0_14_port, Y(50) => P_tmp_0_13_port, 
                           Y(51) => P_tmp_0_12_port, Y(52) => P_tmp_0_11_port, 
                           Y(53) => P_tmp_0_10_port, Y(54) => P_tmp_0_9_port, 
                           Y(55) => P_tmp_0_8_port, Y(56) => P_tmp_0_7_port, 
                           Y(57) => P_tmp_0_6_port, Y(58) => P_tmp_0_5_port, 
                           Y(59) => P_tmp_0_4_port, Y(60) => P_tmp_0_3_port, 
                           Y(61) => P_tmp_0_2_port, Y(62) => P_tmp_0_1_port, 
                           Y(63) => P_tmp_0_0_port);
   MUXi_1 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_15 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_0_63_port, INPUT(65) => 
                           A_pos_shifted_by2_0_62_port, INPUT(66) => 
                           A_pos_shifted_by2_0_61_port, INPUT(67) => 
                           A_pos_shifted_by2_0_60_port, INPUT(68) => 
                           A_pos_shifted_by2_0_59_port, INPUT(69) => 
                           A_pos_shifted_by2_0_58_port, INPUT(70) => 
                           A_pos_shifted_by2_0_57_port, INPUT(71) => 
                           A_pos_shifted_by2_0_56_port, INPUT(72) => 
                           A_pos_shifted_by2_0_55_port, INPUT(73) => 
                           A_pos_shifted_by2_0_54_port, INPUT(74) => 
                           A_pos_shifted_by2_0_53_port, INPUT(75) => 
                           A_pos_shifted_by2_0_52_port, INPUT(76) => 
                           A_pos_shifted_by2_0_51_port, INPUT(77) => 
                           A_pos_shifted_by2_0_50_port, INPUT(78) => 
                           A_pos_shifted_by2_0_49_port, INPUT(79) => 
                           A_pos_shifted_by2_0_48_port, INPUT(80) => n242, 
                           INPUT(81) => A_pos_shifted_by2_0_46_port, INPUT(82) 
                           => A_pos_shifted_by2_0_45_port, INPUT(83) => 
                           A_pos_shifted_by2_0_44_port, INPUT(84) => 
                           A_pos_shifted_by2_0_43_port, INPUT(85) => 
                           A_pos_shifted_by2_0_42_port, INPUT(86) => 
                           A_pos_shifted_by2_0_41_port, INPUT(87) => 
                           A_pos_shifted_by2_0_40_port, INPUT(88) => 
                           A_pos_shifted_by2_0_39_port, INPUT(89) => 
                           A_pos_shifted_by2_0_38_port, INPUT(90) => 
                           A_pos_shifted_by2_0_37_port, INPUT(91) => 
                           A_pos_shifted_by2_0_36_port, INPUT(92) => 
                           A_pos_shifted_by2_0_35_port, INPUT(93) => 
                           A_pos_shifted_by2_0_34_port, INPUT(94) => 
                           A_pos_shifted_by2_0_33_port, INPUT(95) => 
                           A_pos_shifted_by2_0_32_port, INPUT(96) => 
                           A_pos_shifted_by2_0_31_port, INPUT(97) => 
                           A_pos_shifted_by2_0_30_port, INPUT(98) => 
                           A_pos_shifted_by2_0_29_port, INPUT(99) => 
                           A_pos_shifted_by2_0_28_port, INPUT(100) => 
                           A_pos_shifted_by2_0_27_port, INPUT(101) => 
                           A_pos_shifted_by2_0_26_port, INPUT(102) => 
                           A_pos_shifted_by2_0_25_port, INPUT(103) => 
                           A_pos_shifted_by2_0_24_port, INPUT(104) => 
                           A_pos_shifted_by2_0_23_port, INPUT(105) => 
                           A_pos_shifted_by2_0_22_port, INPUT(106) => 
                           A_pos_shifted_by2_0_21_port, INPUT(107) => 
                           A_pos_shifted_by2_0_20_port, INPUT(108) => 
                           A_pos_shifted_by2_0_19_port, INPUT(109) => 
                           A_pos_shifted_by2_0_18_port, INPUT(110) => 
                           A_pos_shifted_by2_0_17_port, INPUT(111) => 
                           A_pos_shifted_by2_0_16_port, INPUT(112) => 
                           A_pos_shifted_by2_0_15_port, INPUT(113) => 
                           A_pos_shifted_by2_0_14_port, INPUT(114) => 
                           A_pos_shifted_by2_0_13_port, INPUT(115) => 
                           A_pos_shifted_by2_0_12_port, INPUT(116) => 
                           A_pos_shifted_by2_0_11_port, INPUT(117) => 
                           A_pos_shifted_by2_0_10_port, INPUT(118) => 
                           A_pos_shifted_by2_0_9_port, INPUT(119) => 
                           A_pos_shifted_by2_0_8_port, INPUT(120) => 
                           A_pos_shifted_by2_0_7_port, INPUT(121) => 
                           A_pos_shifted_by2_0_6_port, INPUT(122) => 
                           A_pos_shifted_by2_0_5_port, INPUT(123) => 
                           A_pos_shifted_by2_0_4_port, INPUT(124) => 
                           A_pos_shifted_by2_0_3_port, INPUT(125) => 
                           A_pos_shifted_by2_0_2_port, INPUT(126) => 
                           A_pos_shifted_by2_0_1_port, INPUT(127) => 
                           A_pos_shifted_by2_0_0_port, INPUT(128) => 
                           A_neg_shifted_by2_0_63_port, INPUT(129) => 
                           A_neg_shifted_by2_0_62_port, INPUT(130) => 
                           A_neg_shifted_by2_0_61_port, INPUT(131) => 
                           A_neg_shifted_by2_0_60_port, INPUT(132) => 
                           A_neg_shifted_by2_0_59_port, INPUT(133) => 
                           A_neg_shifted_by2_0_58_port, INPUT(134) => 
                           A_neg_shifted_by2_0_57_port, INPUT(135) => 
                           A_neg_shifted_by2_0_56_port, INPUT(136) => 
                           A_neg_shifted_by2_0_55_port, INPUT(137) => 
                           A_neg_shifted_by2_0_54_port, INPUT(138) => 
                           A_neg_shifted_by2_0_53_port, INPUT(139) => 
                           A_neg_shifted_by2_0_52_port, INPUT(140) => 
                           A_neg_shifted_by2_0_51_port, INPUT(141) => 
                           A_neg_shifted_by2_0_50_port, INPUT(142) => 
                           A_neg_shifted_by2_0_49_port, INPUT(143) => 
                           A_neg_shifted_by2_0_48_port, INPUT(144) => n207, 
                           INPUT(145) => A_neg_shifted_by2_0_46_port, 
                           INPUT(146) => A_neg_shifted_by2_0_45_port, 
                           INPUT(147) => A_neg_shifted_by2_0_44_port, 
                           INPUT(148) => A_neg_shifted_by2_0_43_port, 
                           INPUT(149) => A_neg_shifted_by2_0_42_port, 
                           INPUT(150) => A_neg_shifted_by2_0_41_port, 
                           INPUT(151) => A_neg_shifted_by2_0_40_port, 
                           INPUT(152) => A_neg_shifted_by2_0_39_port, 
                           INPUT(153) => A_neg_shifted_by2_0_38_port, 
                           INPUT(154) => A_neg_shifted_by2_0_37_port, 
                           INPUT(155) => A_neg_shifted_by2_0_36_port, 
                           INPUT(156) => A_neg_shifted_by2_0_35_port, 
                           INPUT(157) => A_neg_shifted_by2_0_34_port, 
                           INPUT(158) => A_neg_shifted_by2_0_33_port, 
                           INPUT(159) => A_neg_shifted_by2_0_32_port, 
                           INPUT(160) => A_neg_shifted_by2_0_31_port, 
                           INPUT(161) => A_neg_shifted_by2_0_30_port, 
                           INPUT(162) => A_neg_shifted_by2_0_29_port, 
                           INPUT(163) => A_neg_shifted_by2_0_28_port, 
                           INPUT(164) => A_neg_shifted_by2_0_27_port, 
                           INPUT(165) => A_neg_shifted_by2_0_26_port, 
                           INPUT(166) => A_neg_shifted_by2_0_25_port, 
                           INPUT(167) => A_neg_shifted_by2_0_24_port, 
                           INPUT(168) => A_neg_shifted_by2_0_23_port, 
                           INPUT(169) => A_neg_shifted_by2_0_22_port, 
                           INPUT(170) => A_neg_shifted_by2_0_21_port, 
                           INPUT(171) => A_neg_shifted_by2_0_20_port, 
                           INPUT(172) => A_neg_shifted_by2_0_19_port, 
                           INPUT(173) => A_neg_shifted_by2_0_18_port, 
                           INPUT(174) => A_neg_shifted_by2_0_17_port, 
                           INPUT(175) => A_neg_shifted_by2_0_16_port, 
                           INPUT(176) => A_neg_shifted_by2_0_15_port, 
                           INPUT(177) => A_neg_shifted_by2_0_14_port, 
                           INPUT(178) => A_neg_shifted_by2_0_13_port, 
                           INPUT(179) => A_neg_shifted_by2_0_12_port, 
                           INPUT(180) => A_neg_shifted_by2_0_11_port, 
                           INPUT(181) => A_neg_shifted_by2_0_10_port, 
                           INPUT(182) => A_neg_shifted_by2_0_9_port, INPUT(183)
                           => A_neg_shifted_by2_0_8_port, INPUT(184) => 
                           A_neg_shifted_by2_0_7_port, INPUT(185) => 
                           A_neg_shifted_by2_0_6_port, INPUT(186) => 
                           A_neg_shifted_by2_0_5_port, INPUT(187) => 
                           A_neg_shifted_by2_0_4_port, INPUT(188) => 
                           A_neg_shifted_by2_0_3_port, INPUT(189) => 
                           A_neg_shifted_by2_0_2_port, INPUT(190) => 
                           A_neg_shifted_by2_0_1_port, INPUT(191) => 
                           A_neg_shifted_by2_0_0_port, INPUT(192) => 
                           A_pos_shifted_by1_1_63_port, INPUT(193) => 
                           A_pos_shifted_by1_1_62_port, INPUT(194) => 
                           A_pos_shifted_by1_1_61_port, INPUT(195) => 
                           A_pos_shifted_by1_1_60_port, INPUT(196) => 
                           A_pos_shifted_by1_1_59_port, INPUT(197) => 
                           A_pos_shifted_by1_1_58_port, INPUT(198) => 
                           A_pos_shifted_by1_1_57_port, INPUT(199) => 
                           A_pos_shifted_by1_1_56_port, INPUT(200) => 
                           A_pos_shifted_by1_1_55_port, INPUT(201) => 
                           A_pos_shifted_by1_1_54_port, INPUT(202) => 
                           A_pos_shifted_by1_1_53_port, INPUT(203) => 
                           A_pos_shifted_by1_1_52_port, INPUT(204) => 
                           A_pos_shifted_by1_1_51_port, INPUT(205) => 
                           A_pos_shifted_by1_1_50_port, INPUT(206) => 
                           A_pos_shifted_by1_1_49_port, INPUT(207) => 
                           A_pos_shifted_by1_1_48_port, INPUT(208) => 
                           A_pos_shifted_by1_1_47_port, INPUT(209) => 
                           A_pos_shifted_by1_1_46_port, INPUT(210) => 
                           A_pos_shifted_by1_1_45_port, INPUT(211) => 
                           A_pos_shifted_by1_1_44_port, INPUT(212) => 
                           A_pos_shifted_by1_1_43_port, INPUT(213) => 
                           A_pos_shifted_by1_1_42_port, INPUT(214) => 
                           A_pos_shifted_by1_1_41_port, INPUT(215) => 
                           A_pos_shifted_by1_1_40_port, INPUT(216) => 
                           A_pos_shifted_by1_1_39_port, INPUT(217) => 
                           A_pos_shifted_by1_1_38_port, INPUT(218) => 
                           A_pos_shifted_by1_1_37_port, INPUT(219) => 
                           A_pos_shifted_by1_1_36_port, INPUT(220) => 
                           A_pos_shifted_by1_1_35_port, INPUT(221) => 
                           A_pos_shifted_by1_1_34_port, INPUT(222) => 
                           A_pos_shifted_by1_1_33_port, INPUT(223) => 
                           A_pos_shifted_by1_1_32_port, INPUT(224) => 
                           A_pos_shifted_by1_1_31_port, INPUT(225) => 
                           A_pos_shifted_by1_1_30_port, INPUT(226) => 
                           A_pos_shifted_by1_1_29_port, INPUT(227) => 
                           A_pos_shifted_by1_1_28_port, INPUT(228) => 
                           A_pos_shifted_by1_1_27_port, INPUT(229) => 
                           A_pos_shifted_by1_1_26_port, INPUT(230) => 
                           A_pos_shifted_by1_1_25_port, INPUT(231) => 
                           A_pos_shifted_by1_1_24_port, INPUT(232) => 
                           A_pos_shifted_by1_1_23_port, INPUT(233) => 
                           A_pos_shifted_by1_1_22_port, INPUT(234) => 
                           A_pos_shifted_by1_1_21_port, INPUT(235) => 
                           A_pos_shifted_by1_1_20_port, INPUT(236) => 
                           A_pos_shifted_by1_1_19_port, INPUT(237) => 
                           A_pos_shifted_by1_1_18_port, INPUT(238) => 
                           A_pos_shifted_by1_1_17_port, INPUT(239) => 
                           A_pos_shifted_by1_1_16_port, INPUT(240) => 
                           A_pos_shifted_by1_1_15_port, INPUT(241) => 
                           A_pos_shifted_by1_1_14_port, INPUT(242) => 
                           A_pos_shifted_by1_1_13_port, INPUT(243) => 
                           A_pos_shifted_by1_1_12_port, INPUT(244) => 
                           A_pos_shifted_by1_1_11_port, INPUT(245) => 
                           A_pos_shifted_by1_1_10_port, INPUT(246) => 
                           A_pos_shifted_by1_1_9_port, INPUT(247) => 
                           A_pos_shifted_by1_1_8_port, INPUT(248) => 
                           A_pos_shifted_by1_1_7_port, INPUT(249) => 
                           A_pos_shifted_by1_1_6_port, INPUT(250) => 
                           A_pos_shifted_by1_1_5_port, INPUT(251) => 
                           A_pos_shifted_by1_1_4_port, INPUT(252) => 
                           A_pos_shifted_by1_1_3_port, INPUT(253) => 
                           A_pos_shifted_by1_1_2_port, INPUT(254) => 
                           A_pos_shifted_by1_1_1_port, INPUT(255) => 
                           A_pos_shifted_by1_1_0_port, INPUT(256) => 
                           A_neg_shifted_by1_1_63_port, INPUT(257) => 
                           A_neg_shifted_by1_1_62_port, INPUT(258) => 
                           A_neg_shifted_by1_1_61_port, INPUT(259) => 
                           A_neg_shifted_by1_1_60_port, INPUT(260) => 
                           A_neg_shifted_by1_1_59_port, INPUT(261) => 
                           A_neg_shifted_by1_1_58_port, INPUT(262) => 
                           A_neg_shifted_by1_1_57_port, INPUT(263) => 
                           A_neg_shifted_by1_1_56_port, INPUT(264) => 
                           A_neg_shifted_by1_1_55_port, INPUT(265) => 
                           A_neg_shifted_by1_1_54_port, INPUT(266) => 
                           A_neg_shifted_by1_1_53_port, INPUT(267) => 
                           A_neg_shifted_by1_1_52_port, INPUT(268) => 
                           A_neg_shifted_by1_1_51_port, INPUT(269) => 
                           A_neg_shifted_by1_1_50_port, INPUT(270) => 
                           A_neg_shifted_by1_1_49_port, INPUT(271) => 
                           A_neg_shifted_by1_1_48_port, INPUT(272) => 
                           A_neg_shifted_by1_1_47_port, INPUT(273) => 
                           A_neg_shifted_by1_1_46_port, INPUT(274) => 
                           A_neg_shifted_by1_1_45_port, INPUT(275) => 
                           A_neg_shifted_by1_1_44_port, INPUT(276) => 
                           A_neg_shifted_by1_1_43_port, INPUT(277) => 
                           A_neg_shifted_by1_1_42_port, INPUT(278) => 
                           A_neg_shifted_by1_1_41_port, INPUT(279) => 
                           A_neg_shifted_by1_1_40_port, INPUT(280) => 
                           A_neg_shifted_by1_1_39_port, INPUT(281) => 
                           A_neg_shifted_by1_1_38_port, INPUT(282) => 
                           A_neg_shifted_by1_1_37_port, INPUT(283) => 
                           A_neg_shifted_by1_1_36_port, INPUT(284) => 
                           A_neg_shifted_by1_1_35_port, INPUT(285) => 
                           A_neg_shifted_by1_1_34_port, INPUT(286) => 
                           A_neg_shifted_by1_1_33_port, INPUT(287) => 
                           A_neg_shifted_by1_1_32_port, INPUT(288) => 
                           A_neg_shifted_by1_1_31_port, INPUT(289) => 
                           A_neg_shifted_by1_1_30_port, INPUT(290) => 
                           A_neg_shifted_by1_1_29_port, INPUT(291) => 
                           A_neg_shifted_by1_1_28_port, INPUT(292) => 
                           A_neg_shifted_by1_1_27_port, INPUT(293) => 
                           A_neg_shifted_by1_1_26_port, INPUT(294) => 
                           A_neg_shifted_by1_1_25_port, INPUT(295) => 
                           A_neg_shifted_by1_1_24_port, INPUT(296) => 
                           A_neg_shifted_by1_1_23_port, INPUT(297) => 
                           A_neg_shifted_by1_1_22_port, INPUT(298) => 
                           A_neg_shifted_by1_1_21_port, INPUT(299) => 
                           A_neg_shifted_by1_1_20_port, INPUT(300) => 
                           A_neg_shifted_by1_1_19_port, INPUT(301) => 
                           A_neg_shifted_by1_1_18_port, INPUT(302) => 
                           A_neg_shifted_by1_1_17_port, INPUT(303) => 
                           A_neg_shifted_by1_1_16_port, INPUT(304) => 
                           A_neg_shifted_by1_1_15_port, INPUT(305) => 
                           A_neg_shifted_by1_1_14_port, INPUT(306) => 
                           A_neg_shifted_by1_1_13_port, INPUT(307) => 
                           A_neg_shifted_by1_1_12_port, INPUT(308) => 
                           A_neg_shifted_by1_1_11_port, INPUT(309) => 
                           A_neg_shifted_by1_1_10_port, INPUT(310) => 
                           A_neg_shifted_by1_1_9_port, INPUT(311) => 
                           A_neg_shifted_by1_1_8_port, INPUT(312) => 
                           A_neg_shifted_by1_1_7_port, INPUT(313) => 
                           A_neg_shifted_by1_1_6_port, INPUT(314) => 
                           A_neg_shifted_by1_1_5_port, INPUT(315) => 
                           A_neg_shifted_by1_1_4_port, INPUT(316) => 
                           A_neg_shifted_by1_1_3_port, INPUT(317) => 
                           A_neg_shifted_by1_1_2_port, INPUT(318) => 
                           A_neg_shifted_by1_1_1_port, INPUT(319) => 
                           A_neg_shifted_by1_1_0_port, SEL(0) => 
                           selection_signal_1_2_port, SEL(1) => 
                           selection_signal_1_1_port, SEL(2) => 
                           selection_signal_1_0_port, Y(0) => OUT_MUX_1_63_port
                           , Y(1) => OUT_MUX_1_62_port, Y(2) => 
                           OUT_MUX_1_61_port, Y(3) => OUT_MUX_1_60_port, Y(4) 
                           => OUT_MUX_1_59_port, Y(5) => OUT_MUX_1_58_port, 
                           Y(6) => OUT_MUX_1_57_port, Y(7) => OUT_MUX_1_56_port
                           , Y(8) => OUT_MUX_1_55_port, Y(9) => 
                           OUT_MUX_1_54_port, Y(10) => OUT_MUX_1_53_port, Y(11)
                           => OUT_MUX_1_52_port, Y(12) => OUT_MUX_1_51_port, 
                           Y(13) => OUT_MUX_1_50_port, Y(14) => 
                           OUT_MUX_1_49_port, Y(15) => OUT_MUX_1_48_port, Y(16)
                           => OUT_MUX_1_47_port, Y(17) => OUT_MUX_1_46_port, 
                           Y(18) => OUT_MUX_1_45_port, Y(19) => 
                           OUT_MUX_1_44_port, Y(20) => OUT_MUX_1_43_port, Y(21)
                           => OUT_MUX_1_42_port, Y(22) => OUT_MUX_1_41_port, 
                           Y(23) => OUT_MUX_1_40_port, Y(24) => 
                           OUT_MUX_1_39_port, Y(25) => OUT_MUX_1_38_port, Y(26)
                           => OUT_MUX_1_37_port, Y(27) => OUT_MUX_1_36_port, 
                           Y(28) => OUT_MUX_1_35_port, Y(29) => 
                           OUT_MUX_1_34_port, Y(30) => OUT_MUX_1_33_port, Y(31)
                           => OUT_MUX_1_32_port, Y(32) => OUT_MUX_1_31_port, 
                           Y(33) => OUT_MUX_1_30_port, Y(34) => 
                           OUT_MUX_1_29_port, Y(35) => OUT_MUX_1_28_port, Y(36)
                           => OUT_MUX_1_27_port, Y(37) => OUT_MUX_1_26_port, 
                           Y(38) => OUT_MUX_1_25_port, Y(39) => 
                           OUT_MUX_1_24_port, Y(40) => OUT_MUX_1_23_port, Y(41)
                           => OUT_MUX_1_22_port, Y(42) => OUT_MUX_1_21_port, 
                           Y(43) => OUT_MUX_1_20_port, Y(44) => 
                           OUT_MUX_1_19_port, Y(45) => OUT_MUX_1_18_port, Y(46)
                           => OUT_MUX_1_17_port, Y(47) => OUT_MUX_1_16_port, 
                           Y(48) => OUT_MUX_1_15_port, Y(49) => 
                           OUT_MUX_1_14_port, Y(50) => OUT_MUX_1_13_port, Y(51)
                           => OUT_MUX_1_12_port, Y(52) => OUT_MUX_1_11_port, 
                           Y(53) => OUT_MUX_1_10_port, Y(54) => 
                           OUT_MUX_1_9_port, Y(55) => OUT_MUX_1_8_port, Y(56) 
                           => OUT_MUX_1_7_port, Y(57) => OUT_MUX_1_6_port, 
                           Y(58) => OUT_MUX_1_5_port, Y(59) => OUT_MUX_1_4_port
                           , Y(60) => OUT_MUX_1_3_port, Y(61) => 
                           OUT_MUX_1_2_port, Y(62) => OUT_MUX_1_1_port, Y(63) 
                           => OUT_MUX_1_0_port);
   MUXi_2 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_14 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_1_63_port, INPUT(65) => 
                           A_pos_shifted_by2_1_62_port, INPUT(66) => 
                           A_pos_shifted_by2_1_61_port, INPUT(67) => 
                           A_pos_shifted_by2_1_60_port, INPUT(68) => 
                           A_pos_shifted_by2_1_59_port, INPUT(69) => 
                           A_pos_shifted_by2_1_58_port, INPUT(70) => 
                           A_pos_shifted_by2_1_57_port, INPUT(71) => 
                           A_pos_shifted_by2_1_56_port, INPUT(72) => 
                           A_pos_shifted_by2_1_55_port, INPUT(73) => 
                           A_pos_shifted_by2_1_54_port, INPUT(74) => 
                           A_pos_shifted_by2_1_53_port, INPUT(75) => 
                           A_pos_shifted_by2_1_52_port, INPUT(76) => 
                           A_pos_shifted_by2_1_51_port, INPUT(77) => 
                           A_pos_shifted_by2_1_50_port, INPUT(78) => 
                           A_pos_shifted_by2_1_49_port, INPUT(79) => 
                           A_pos_shifted_by2_1_48_port, INPUT(80) => n241, 
                           INPUT(81) => A_pos_shifted_by2_1_46_port, INPUT(82) 
                           => A_pos_shifted_by2_1_45_port, INPUT(83) => 
                           A_pos_shifted_by2_1_44_port, INPUT(84) => 
                           A_pos_shifted_by2_1_43_port, INPUT(85) => 
                           A_pos_shifted_by2_1_42_port, INPUT(86) => 
                           A_pos_shifted_by2_1_41_port, INPUT(87) => 
                           A_pos_shifted_by2_1_40_port, INPUT(88) => 
                           A_pos_shifted_by2_1_39_port, INPUT(89) => 
                           A_pos_shifted_by2_1_38_port, INPUT(90) => 
                           A_pos_shifted_by2_1_37_port, INPUT(91) => 
                           A_pos_shifted_by2_1_36_port, INPUT(92) => 
                           A_pos_shifted_by2_1_35_port, INPUT(93) => 
                           A_pos_shifted_by2_1_34_port, INPUT(94) => 
                           A_pos_shifted_by2_1_33_port, INPUT(95) => 
                           A_pos_shifted_by2_1_32_port, INPUT(96) => 
                           A_pos_shifted_by2_1_31_port, INPUT(97) => 
                           A_pos_shifted_by2_1_30_port, INPUT(98) => 
                           A_pos_shifted_by2_1_29_port, INPUT(99) => 
                           A_pos_shifted_by2_1_28_port, INPUT(100) => 
                           A_pos_shifted_by2_1_27_port, INPUT(101) => 
                           A_pos_shifted_by2_1_26_port, INPUT(102) => 
                           A_pos_shifted_by2_1_25_port, INPUT(103) => 
                           A_pos_shifted_by2_1_24_port, INPUT(104) => 
                           A_pos_shifted_by2_1_23_port, INPUT(105) => 
                           A_pos_shifted_by2_1_22_port, INPUT(106) => 
                           A_pos_shifted_by2_1_21_port, INPUT(107) => 
                           A_pos_shifted_by2_1_20_port, INPUT(108) => 
                           A_pos_shifted_by2_1_19_port, INPUT(109) => 
                           A_pos_shifted_by2_1_18_port, INPUT(110) => 
                           A_pos_shifted_by2_1_17_port, INPUT(111) => 
                           A_pos_shifted_by2_1_16_port, INPUT(112) => 
                           A_pos_shifted_by2_1_15_port, INPUT(113) => 
                           A_pos_shifted_by2_1_14_port, INPUT(114) => 
                           A_pos_shifted_by2_1_13_port, INPUT(115) => 
                           A_pos_shifted_by2_1_12_port, INPUT(116) => 
                           A_pos_shifted_by2_1_11_port, INPUT(117) => 
                           A_pos_shifted_by2_1_10_port, INPUT(118) => 
                           A_pos_shifted_by2_1_9_port, INPUT(119) => 
                           A_pos_shifted_by2_1_8_port, INPUT(120) => 
                           A_pos_shifted_by2_1_7_port, INPUT(121) => 
                           A_pos_shifted_by2_1_6_port, INPUT(122) => 
                           A_pos_shifted_by2_1_5_port, INPUT(123) => 
                           A_pos_shifted_by2_1_4_port, INPUT(124) => 
                           A_pos_shifted_by2_1_3_port, INPUT(125) => 
                           A_pos_shifted_by2_1_2_port, INPUT(126) => 
                           A_pos_shifted_by2_1_1_port, INPUT(127) => 
                           A_pos_shifted_by2_1_0_port, INPUT(128) => 
                           A_neg_shifted_by2_1_63_port, INPUT(129) => 
                           A_neg_shifted_by2_1_62_port, INPUT(130) => 
                           A_neg_shifted_by2_1_61_port, INPUT(131) => 
                           A_neg_shifted_by2_1_60_port, INPUT(132) => 
                           A_neg_shifted_by2_1_59_port, INPUT(133) => 
                           A_neg_shifted_by2_1_58_port, INPUT(134) => 
                           A_neg_shifted_by2_1_57_port, INPUT(135) => 
                           A_neg_shifted_by2_1_56_port, INPUT(136) => 
                           A_neg_shifted_by2_1_55_port, INPUT(137) => 
                           A_neg_shifted_by2_1_54_port, INPUT(138) => 
                           A_neg_shifted_by2_1_53_port, INPUT(139) => 
                           A_neg_shifted_by2_1_52_port, INPUT(140) => 
                           A_neg_shifted_by2_1_51_port, INPUT(141) => 
                           A_neg_shifted_by2_1_50_port, INPUT(142) => 
                           A_neg_shifted_by2_1_49_port, INPUT(143) => 
                           A_neg_shifted_by2_1_48_port, INPUT(144) => n206, 
                           INPUT(145) => A_neg_shifted_by2_1_46_port, 
                           INPUT(146) => A_neg_shifted_by2_1_45_port, 
                           INPUT(147) => A_neg_shifted_by2_1_44_port, 
                           INPUT(148) => A_neg_shifted_by2_1_43_port, 
                           INPUT(149) => A_neg_shifted_by2_1_42_port, 
                           INPUT(150) => A_neg_shifted_by2_1_41_port, 
                           INPUT(151) => A_neg_shifted_by2_1_40_port, 
                           INPUT(152) => A_neg_shifted_by2_1_39_port, 
                           INPUT(153) => A_neg_shifted_by2_1_38_port, 
                           INPUT(154) => A_neg_shifted_by2_1_37_port, 
                           INPUT(155) => A_neg_shifted_by2_1_36_port, 
                           INPUT(156) => A_neg_shifted_by2_1_35_port, 
                           INPUT(157) => A_neg_shifted_by2_1_34_port, 
                           INPUT(158) => A_neg_shifted_by2_1_33_port, 
                           INPUT(159) => A_neg_shifted_by2_1_32_port, 
                           INPUT(160) => A_neg_shifted_by2_1_31_port, 
                           INPUT(161) => A_neg_shifted_by2_1_30_port, 
                           INPUT(162) => A_neg_shifted_by2_1_29_port, 
                           INPUT(163) => A_neg_shifted_by2_1_28_port, 
                           INPUT(164) => A_neg_shifted_by2_1_27_port, 
                           INPUT(165) => A_neg_shifted_by2_1_26_port, 
                           INPUT(166) => A_neg_shifted_by2_1_25_port, 
                           INPUT(167) => A_neg_shifted_by2_1_24_port, 
                           INPUT(168) => A_neg_shifted_by2_1_23_port, 
                           INPUT(169) => A_neg_shifted_by2_1_22_port, 
                           INPUT(170) => A_neg_shifted_by2_1_21_port, 
                           INPUT(171) => A_neg_shifted_by2_1_20_port, 
                           INPUT(172) => A_neg_shifted_by2_1_19_port, 
                           INPUT(173) => A_neg_shifted_by2_1_18_port, 
                           INPUT(174) => A_neg_shifted_by2_1_17_port, 
                           INPUT(175) => A_neg_shifted_by2_1_16_port, 
                           INPUT(176) => A_neg_shifted_by2_1_15_port, 
                           INPUT(177) => A_neg_shifted_by2_1_14_port, 
                           INPUT(178) => A_neg_shifted_by2_1_13_port, 
                           INPUT(179) => A_neg_shifted_by2_1_12_port, 
                           INPUT(180) => A_neg_shifted_by2_1_11_port, 
                           INPUT(181) => A_neg_shifted_by2_1_10_port, 
                           INPUT(182) => A_neg_shifted_by2_1_9_port, INPUT(183)
                           => A_neg_shifted_by2_1_8_port, INPUT(184) => 
                           A_neg_shifted_by2_1_7_port, INPUT(185) => 
                           A_neg_shifted_by2_1_6_port, INPUT(186) => 
                           A_neg_shifted_by2_1_5_port, INPUT(187) => 
                           A_neg_shifted_by2_1_4_port, INPUT(188) => 
                           A_neg_shifted_by2_1_3_port, INPUT(189) => 
                           A_neg_shifted_by2_1_2_port, INPUT(190) => 
                           A_neg_shifted_by2_1_1_port, INPUT(191) => 
                           A_neg_shifted_by2_1_0_port, INPUT(192) => 
                           A_pos_shifted_by1_2_63_port, INPUT(193) => 
                           A_pos_shifted_by1_2_62_port, INPUT(194) => 
                           A_pos_shifted_by1_2_61_port, INPUT(195) => 
                           A_pos_shifted_by1_2_60_port, INPUT(196) => 
                           A_pos_shifted_by1_2_59_port, INPUT(197) => 
                           A_pos_shifted_by1_2_58_port, INPUT(198) => 
                           A_pos_shifted_by1_2_57_port, INPUT(199) => 
                           A_pos_shifted_by1_2_56_port, INPUT(200) => 
                           A_pos_shifted_by1_2_55_port, INPUT(201) => 
                           A_pos_shifted_by1_2_54_port, INPUT(202) => 
                           A_pos_shifted_by1_2_53_port, INPUT(203) => 
                           A_pos_shifted_by1_2_52_port, INPUT(204) => 
                           A_pos_shifted_by1_2_51_port, INPUT(205) => 
                           A_pos_shifted_by1_2_50_port, INPUT(206) => 
                           A_pos_shifted_by1_2_49_port, INPUT(207) => 
                           A_pos_shifted_by1_2_48_port, INPUT(208) => 
                           A_pos_shifted_by1_2_47_port, INPUT(209) => 
                           A_pos_shifted_by1_2_46_port, INPUT(210) => 
                           A_pos_shifted_by1_2_45_port, INPUT(211) => 
                           A_pos_shifted_by1_2_44_port, INPUT(212) => 
                           A_pos_shifted_by1_2_43_port, INPUT(213) => 
                           A_pos_shifted_by1_2_42_port, INPUT(214) => 
                           A_pos_shifted_by1_2_41_port, INPUT(215) => 
                           A_pos_shifted_by1_2_40_port, INPUT(216) => 
                           A_pos_shifted_by1_2_39_port, INPUT(217) => 
                           A_pos_shifted_by1_2_38_port, INPUT(218) => 
                           A_pos_shifted_by1_2_37_port, INPUT(219) => 
                           A_pos_shifted_by1_2_36_port, INPUT(220) => 
                           A_pos_shifted_by1_2_35_port, INPUT(221) => 
                           A_pos_shifted_by1_2_34_port, INPUT(222) => 
                           A_pos_shifted_by1_2_33_port, INPUT(223) => 
                           A_pos_shifted_by1_2_32_port, INPUT(224) => 
                           A_pos_shifted_by1_2_31_port, INPUT(225) => 
                           A_pos_shifted_by1_2_30_port, INPUT(226) => 
                           A_pos_shifted_by1_2_29_port, INPUT(227) => 
                           A_pos_shifted_by1_2_28_port, INPUT(228) => 
                           A_pos_shifted_by1_2_27_port, INPUT(229) => 
                           A_pos_shifted_by1_2_26_port, INPUT(230) => 
                           A_pos_shifted_by1_2_25_port, INPUT(231) => 
                           A_pos_shifted_by1_2_24_port, INPUT(232) => 
                           A_pos_shifted_by1_2_23_port, INPUT(233) => 
                           A_pos_shifted_by1_2_22_port, INPUT(234) => 
                           A_pos_shifted_by1_2_21_port, INPUT(235) => 
                           A_pos_shifted_by1_2_20_port, INPUT(236) => 
                           A_pos_shifted_by1_2_19_port, INPUT(237) => 
                           A_pos_shifted_by1_2_18_port, INPUT(238) => 
                           A_pos_shifted_by1_2_17_port, INPUT(239) => 
                           A_pos_shifted_by1_2_16_port, INPUT(240) => 
                           A_pos_shifted_by1_2_15_port, INPUT(241) => 
                           A_pos_shifted_by1_2_14_port, INPUT(242) => 
                           A_pos_shifted_by1_2_13_port, INPUT(243) => 
                           A_pos_shifted_by1_2_12_port, INPUT(244) => 
                           A_pos_shifted_by1_2_11_port, INPUT(245) => 
                           A_pos_shifted_by1_2_10_port, INPUT(246) => 
                           A_pos_shifted_by1_2_9_port, INPUT(247) => 
                           A_pos_shifted_by1_2_8_port, INPUT(248) => 
                           A_pos_shifted_by1_2_7_port, INPUT(249) => 
                           A_pos_shifted_by1_2_6_port, INPUT(250) => 
                           A_pos_shifted_by1_2_5_port, INPUT(251) => 
                           A_pos_shifted_by1_2_4_port, INPUT(252) => 
                           A_pos_shifted_by1_2_3_port, INPUT(253) => 
                           A_pos_shifted_by1_2_2_port, INPUT(254) => 
                           A_pos_shifted_by1_2_1_port, INPUT(255) => 
                           A_pos_shifted_by1_2_0_port, INPUT(256) => 
                           A_neg_shifted_by1_2_63_port, INPUT(257) => 
                           A_neg_shifted_by1_2_62_port, INPUT(258) => 
                           A_neg_shifted_by1_2_61_port, INPUT(259) => 
                           A_neg_shifted_by1_2_60_port, INPUT(260) => 
                           A_neg_shifted_by1_2_59_port, INPUT(261) => 
                           A_neg_shifted_by1_2_58_port, INPUT(262) => 
                           A_neg_shifted_by1_2_57_port, INPUT(263) => 
                           A_neg_shifted_by1_2_56_port, INPUT(264) => 
                           A_neg_shifted_by1_2_55_port, INPUT(265) => 
                           A_neg_shifted_by1_2_54_port, INPUT(266) => 
                           A_neg_shifted_by1_2_53_port, INPUT(267) => 
                           A_neg_shifted_by1_2_52_port, INPUT(268) => 
                           A_neg_shifted_by1_2_51_port, INPUT(269) => 
                           A_neg_shifted_by1_2_50_port, INPUT(270) => 
                           A_neg_shifted_by1_2_49_port, INPUT(271) => 
                           A_neg_shifted_by1_2_48_port, INPUT(272) => 
                           A_neg_shifted_by1_2_47_port, INPUT(273) => 
                           A_neg_shifted_by1_2_46_port, INPUT(274) => 
                           A_neg_shifted_by1_2_45_port, INPUT(275) => 
                           A_neg_shifted_by1_2_44_port, INPUT(276) => 
                           A_neg_shifted_by1_2_43_port, INPUT(277) => 
                           A_neg_shifted_by1_2_42_port, INPUT(278) => 
                           A_neg_shifted_by1_2_41_port, INPUT(279) => 
                           A_neg_shifted_by1_2_40_port, INPUT(280) => 
                           A_neg_shifted_by1_2_39_port, INPUT(281) => 
                           A_neg_shifted_by1_2_38_port, INPUT(282) => 
                           A_neg_shifted_by1_2_37_port, INPUT(283) => 
                           A_neg_shifted_by1_2_36_port, INPUT(284) => 
                           A_neg_shifted_by1_2_35_port, INPUT(285) => 
                           A_neg_shifted_by1_2_34_port, INPUT(286) => 
                           A_neg_shifted_by1_2_33_port, INPUT(287) => 
                           A_neg_shifted_by1_2_32_port, INPUT(288) => 
                           A_neg_shifted_by1_2_31_port, INPUT(289) => 
                           A_neg_shifted_by1_2_30_port, INPUT(290) => 
                           A_neg_shifted_by1_2_29_port, INPUT(291) => 
                           A_neg_shifted_by1_2_28_port, INPUT(292) => 
                           A_neg_shifted_by1_2_27_port, INPUT(293) => 
                           A_neg_shifted_by1_2_26_port, INPUT(294) => 
                           A_neg_shifted_by1_2_25_port, INPUT(295) => 
                           A_neg_shifted_by1_2_24_port, INPUT(296) => 
                           A_neg_shifted_by1_2_23_port, INPUT(297) => 
                           A_neg_shifted_by1_2_22_port, INPUT(298) => 
                           A_neg_shifted_by1_2_21_port, INPUT(299) => 
                           A_neg_shifted_by1_2_20_port, INPUT(300) => 
                           A_neg_shifted_by1_2_19_port, INPUT(301) => 
                           A_neg_shifted_by1_2_18_port, INPUT(302) => 
                           A_neg_shifted_by1_2_17_port, INPUT(303) => 
                           A_neg_shifted_by1_2_16_port, INPUT(304) => 
                           A_neg_shifted_by1_2_15_port, INPUT(305) => 
                           A_neg_shifted_by1_2_14_port, INPUT(306) => 
                           A_neg_shifted_by1_2_13_port, INPUT(307) => 
                           A_neg_shifted_by1_2_12_port, INPUT(308) => 
                           A_neg_shifted_by1_2_11_port, INPUT(309) => 
                           A_neg_shifted_by1_2_10_port, INPUT(310) => 
                           A_neg_shifted_by1_2_9_port, INPUT(311) => 
                           A_neg_shifted_by1_2_8_port, INPUT(312) => 
                           A_neg_shifted_by1_2_7_port, INPUT(313) => 
                           A_neg_shifted_by1_2_6_port, INPUT(314) => 
                           A_neg_shifted_by1_2_5_port, INPUT(315) => 
                           A_neg_shifted_by1_2_4_port, INPUT(316) => 
                           A_neg_shifted_by1_2_3_port, INPUT(317) => 
                           A_neg_shifted_by1_2_2_port, INPUT(318) => 
                           A_neg_shifted_by1_2_1_port, INPUT(319) => 
                           A_neg_shifted_by1_2_0_port, SEL(0) => 
                           selection_signal_2_2_port, SEL(1) => 
                           selection_signal_2_1_port, SEL(2) => 
                           selection_signal_2_0_port, Y(0) => OUT_MUX_2_63_port
                           , Y(1) => OUT_MUX_2_62_port, Y(2) => 
                           OUT_MUX_2_61_port, Y(3) => OUT_MUX_2_60_port, Y(4) 
                           => OUT_MUX_2_59_port, Y(5) => OUT_MUX_2_58_port, 
                           Y(6) => OUT_MUX_2_57_port, Y(7) => OUT_MUX_2_56_port
                           , Y(8) => OUT_MUX_2_55_port, Y(9) => 
                           OUT_MUX_2_54_port, Y(10) => OUT_MUX_2_53_port, Y(11)
                           => OUT_MUX_2_52_port, Y(12) => OUT_MUX_2_51_port, 
                           Y(13) => OUT_MUX_2_50_port, Y(14) => 
                           OUT_MUX_2_49_port, Y(15) => OUT_MUX_2_48_port, Y(16)
                           => OUT_MUX_2_47_port, Y(17) => OUT_MUX_2_46_port, 
                           Y(18) => OUT_MUX_2_45_port, Y(19) => 
                           OUT_MUX_2_44_port, Y(20) => OUT_MUX_2_43_port, Y(21)
                           => OUT_MUX_2_42_port, Y(22) => OUT_MUX_2_41_port, 
                           Y(23) => OUT_MUX_2_40_port, Y(24) => 
                           OUT_MUX_2_39_port, Y(25) => OUT_MUX_2_38_port, Y(26)
                           => OUT_MUX_2_37_port, Y(27) => OUT_MUX_2_36_port, 
                           Y(28) => OUT_MUX_2_35_port, Y(29) => 
                           OUT_MUX_2_34_port, Y(30) => OUT_MUX_2_33_port, Y(31)
                           => OUT_MUX_2_32_port, Y(32) => OUT_MUX_2_31_port, 
                           Y(33) => OUT_MUX_2_30_port, Y(34) => 
                           OUT_MUX_2_29_port, Y(35) => OUT_MUX_2_28_port, Y(36)
                           => OUT_MUX_2_27_port, Y(37) => OUT_MUX_2_26_port, 
                           Y(38) => OUT_MUX_2_25_port, Y(39) => 
                           OUT_MUX_2_24_port, Y(40) => OUT_MUX_2_23_port, Y(41)
                           => OUT_MUX_2_22_port, Y(42) => OUT_MUX_2_21_port, 
                           Y(43) => OUT_MUX_2_20_port, Y(44) => 
                           OUT_MUX_2_19_port, Y(45) => OUT_MUX_2_18_port, Y(46)
                           => OUT_MUX_2_17_port, Y(47) => OUT_MUX_2_16_port, 
                           Y(48) => OUT_MUX_2_15_port, Y(49) => 
                           OUT_MUX_2_14_port, Y(50) => OUT_MUX_2_13_port, Y(51)
                           => OUT_MUX_2_12_port, Y(52) => OUT_MUX_2_11_port, 
                           Y(53) => OUT_MUX_2_10_port, Y(54) => 
                           OUT_MUX_2_9_port, Y(55) => OUT_MUX_2_8_port, Y(56) 
                           => OUT_MUX_2_7_port, Y(57) => OUT_MUX_2_6_port, 
                           Y(58) => OUT_MUX_2_5_port, Y(59) => OUT_MUX_2_4_port
                           , Y(60) => OUT_MUX_2_3_port, Y(61) => 
                           OUT_MUX_2_2_port, Y(62) => OUT_MUX_2_1_port, Y(63) 
                           => OUT_MUX_2_0_port);
   MUXi_3 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_13 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_2_63_port, INPUT(65) => 
                           A_pos_shifted_by2_2_62_port, INPUT(66) => 
                           A_pos_shifted_by2_2_61_port, INPUT(67) => 
                           A_pos_shifted_by2_2_60_port, INPUT(68) => 
                           A_pos_shifted_by2_2_59_port, INPUT(69) => 
                           A_pos_shifted_by2_2_58_port, INPUT(70) => 
                           A_pos_shifted_by2_2_57_port, INPUT(71) => 
                           A_pos_shifted_by2_2_56_port, INPUT(72) => 
                           A_pos_shifted_by2_2_55_port, INPUT(73) => 
                           A_pos_shifted_by2_2_54_port, INPUT(74) => 
                           A_pos_shifted_by2_2_53_port, INPUT(75) => 
                           A_pos_shifted_by2_2_52_port, INPUT(76) => 
                           A_pos_shifted_by2_2_51_port, INPUT(77) => 
                           A_pos_shifted_by2_2_50_port, INPUT(78) => 
                           A_pos_shifted_by2_2_49_port, INPUT(79) => 
                           A_pos_shifted_by2_2_48_port, INPUT(80) => n240, 
                           INPUT(81) => A_pos_shifted_by2_2_46_port, INPUT(82) 
                           => A_pos_shifted_by2_2_45_port, INPUT(83) => 
                           A_pos_shifted_by2_2_44_port, INPUT(84) => 
                           A_pos_shifted_by2_2_43_port, INPUT(85) => 
                           A_pos_shifted_by2_2_42_port, INPUT(86) => 
                           A_pos_shifted_by2_2_41_port, INPUT(87) => 
                           A_pos_shifted_by2_2_40_port, INPUT(88) => 
                           A_pos_shifted_by2_2_39_port, INPUT(89) => 
                           A_pos_shifted_by2_2_38_port, INPUT(90) => 
                           A_pos_shifted_by2_2_37_port, INPUT(91) => 
                           A_pos_shifted_by2_2_36_port, INPUT(92) => 
                           A_pos_shifted_by2_2_35_port, INPUT(93) => 
                           A_pos_shifted_by2_2_34_port, INPUT(94) => 
                           A_pos_shifted_by2_2_33_port, INPUT(95) => 
                           A_pos_shifted_by2_2_32_port, INPUT(96) => 
                           A_pos_shifted_by2_2_31_port, INPUT(97) => 
                           A_pos_shifted_by2_2_30_port, INPUT(98) => 
                           A_pos_shifted_by2_2_29_port, INPUT(99) => 
                           A_pos_shifted_by2_2_28_port, INPUT(100) => 
                           A_pos_shifted_by2_2_27_port, INPUT(101) => 
                           A_pos_shifted_by2_2_26_port, INPUT(102) => 
                           A_pos_shifted_by2_2_25_port, INPUT(103) => 
                           A_pos_shifted_by2_2_24_port, INPUT(104) => 
                           A_pos_shifted_by2_2_23_port, INPUT(105) => 
                           A_pos_shifted_by2_2_22_port, INPUT(106) => 
                           A_pos_shifted_by2_2_21_port, INPUT(107) => 
                           A_pos_shifted_by2_2_20_port, INPUT(108) => 
                           A_pos_shifted_by2_2_19_port, INPUT(109) => 
                           A_pos_shifted_by2_2_18_port, INPUT(110) => 
                           A_pos_shifted_by2_2_17_port, INPUT(111) => 
                           A_pos_shifted_by2_2_16_port, INPUT(112) => 
                           A_pos_shifted_by2_2_15_port, INPUT(113) => 
                           A_pos_shifted_by2_2_14_port, INPUT(114) => 
                           A_pos_shifted_by2_2_13_port, INPUT(115) => 
                           A_pos_shifted_by2_2_12_port, INPUT(116) => 
                           A_pos_shifted_by2_2_11_port, INPUT(117) => 
                           A_pos_shifted_by2_2_10_port, INPUT(118) => 
                           A_pos_shifted_by2_2_9_port, INPUT(119) => 
                           A_pos_shifted_by2_2_8_port, INPUT(120) => 
                           A_pos_shifted_by2_2_7_port, INPUT(121) => 
                           A_pos_shifted_by2_2_6_port, INPUT(122) => 
                           A_pos_shifted_by2_2_5_port, INPUT(123) => 
                           A_pos_shifted_by2_2_4_port, INPUT(124) => 
                           A_pos_shifted_by2_2_3_port, INPUT(125) => 
                           A_pos_shifted_by2_2_2_port, INPUT(126) => 
                           A_pos_shifted_by2_2_1_port, INPUT(127) => 
                           A_pos_shifted_by2_2_0_port, INPUT(128) => 
                           A_neg_shifted_by2_2_63_port, INPUT(129) => 
                           A_neg_shifted_by2_2_62_port, INPUT(130) => 
                           A_neg_shifted_by2_2_61_port, INPUT(131) => 
                           A_neg_shifted_by2_2_60_port, INPUT(132) => 
                           A_neg_shifted_by2_2_59_port, INPUT(133) => 
                           A_neg_shifted_by2_2_58_port, INPUT(134) => 
                           A_neg_shifted_by2_2_57_port, INPUT(135) => 
                           A_neg_shifted_by2_2_56_port, INPUT(136) => 
                           A_neg_shifted_by2_2_55_port, INPUT(137) => 
                           A_neg_shifted_by2_2_54_port, INPUT(138) => 
                           A_neg_shifted_by2_2_53_port, INPUT(139) => 
                           A_neg_shifted_by2_2_52_port, INPUT(140) => 
                           A_neg_shifted_by2_2_51_port, INPUT(141) => 
                           A_neg_shifted_by2_2_50_port, INPUT(142) => 
                           A_neg_shifted_by2_2_49_port, INPUT(143) => 
                           A_neg_shifted_by2_2_48_port, INPUT(144) => 
                           A_neg_shifted_by2_2_47_port, INPUT(145) => 
                           A_neg_shifted_by2_2_46_port, INPUT(146) => 
                           A_neg_shifted_by2_2_45_port, INPUT(147) => 
                           A_neg_shifted_by2_2_44_port, INPUT(148) => 
                           A_neg_shifted_by2_2_43_port, INPUT(149) => 
                           A_neg_shifted_by2_2_42_port, INPUT(150) => 
                           A_neg_shifted_by2_2_41_port, INPUT(151) => 
                           A_neg_shifted_by2_2_40_port, INPUT(152) => 
                           A_neg_shifted_by2_2_39_port, INPUT(153) => 
                           A_neg_shifted_by2_2_38_port, INPUT(154) => 
                           A_neg_shifted_by2_2_37_port, INPUT(155) => 
                           A_neg_shifted_by2_2_36_port, INPUT(156) => 
                           A_neg_shifted_by2_2_35_port, INPUT(157) => 
                           A_neg_shifted_by2_2_34_port, INPUT(158) => 
                           A_neg_shifted_by2_2_33_port, INPUT(159) => 
                           A_neg_shifted_by2_2_32_port, INPUT(160) => 
                           A_neg_shifted_by2_2_31_port, INPUT(161) => 
                           A_neg_shifted_by2_2_30_port, INPUT(162) => 
                           A_neg_shifted_by2_2_29_port, INPUT(163) => 
                           A_neg_shifted_by2_2_28_port, INPUT(164) => 
                           A_neg_shifted_by2_2_27_port, INPUT(165) => 
                           A_neg_shifted_by2_2_26_port, INPUT(166) => 
                           A_neg_shifted_by2_2_25_port, INPUT(167) => 
                           A_neg_shifted_by2_2_24_port, INPUT(168) => 
                           A_neg_shifted_by2_2_23_port, INPUT(169) => 
                           A_neg_shifted_by2_2_22_port, INPUT(170) => 
                           A_neg_shifted_by2_2_21_port, INPUT(171) => 
                           A_neg_shifted_by2_2_20_port, INPUT(172) => 
                           A_neg_shifted_by2_2_19_port, INPUT(173) => 
                           A_neg_shifted_by2_2_18_port, INPUT(174) => 
                           A_neg_shifted_by2_2_17_port, INPUT(175) => 
                           A_neg_shifted_by2_2_16_port, INPUT(176) => 
                           A_neg_shifted_by2_2_15_port, INPUT(177) => 
                           A_neg_shifted_by2_2_14_port, INPUT(178) => 
                           A_neg_shifted_by2_2_13_port, INPUT(179) => 
                           A_neg_shifted_by2_2_12_port, INPUT(180) => 
                           A_neg_shifted_by2_2_11_port, INPUT(181) => 
                           A_neg_shifted_by2_2_10_port, INPUT(182) => 
                           A_neg_shifted_by2_2_9_port, INPUT(183) => 
                           A_neg_shifted_by2_2_8_port, INPUT(184) => 
                           A_neg_shifted_by2_2_7_port, INPUT(185) => 
                           A_neg_shifted_by2_2_6_port, INPUT(186) => 
                           A_neg_shifted_by2_2_5_port, INPUT(187) => 
                           A_neg_shifted_by2_2_4_port, INPUT(188) => 
                           A_neg_shifted_by2_2_3_port, INPUT(189) => 
                           A_neg_shifted_by2_2_2_port, INPUT(190) => 
                           A_neg_shifted_by2_2_1_port, INPUT(191) => 
                           A_neg_shifted_by2_2_0_port, INPUT(192) => 
                           A_pos_shifted_by1_3_63_port, INPUT(193) => 
                           A_pos_shifted_by1_3_62_port, INPUT(194) => 
                           A_pos_shifted_by1_3_61_port, INPUT(195) => 
                           A_pos_shifted_by1_3_60_port, INPUT(196) => 
                           A_pos_shifted_by1_3_59_port, INPUT(197) => 
                           A_pos_shifted_by1_3_58_port, INPUT(198) => 
                           A_pos_shifted_by1_3_57_port, INPUT(199) => 
                           A_pos_shifted_by1_3_56_port, INPUT(200) => 
                           A_pos_shifted_by1_3_55_port, INPUT(201) => 
                           A_pos_shifted_by1_3_54_port, INPUT(202) => 
                           A_pos_shifted_by1_3_53_port, INPUT(203) => 
                           A_pos_shifted_by1_3_52_port, INPUT(204) => 
                           A_pos_shifted_by1_3_51_port, INPUT(205) => 
                           A_pos_shifted_by1_3_50_port, INPUT(206) => 
                           A_pos_shifted_by1_3_49_port, INPUT(207) => 
                           A_pos_shifted_by1_3_48_port, INPUT(208) => 
                           A_pos_shifted_by1_3_47_port, INPUT(209) => 
                           A_pos_shifted_by1_3_46_port, INPUT(210) => 
                           A_pos_shifted_by1_3_45_port, INPUT(211) => 
                           A_pos_shifted_by1_3_44_port, INPUT(212) => 
                           A_pos_shifted_by1_3_43_port, INPUT(213) => 
                           A_pos_shifted_by1_3_42_port, INPUT(214) => 
                           A_pos_shifted_by1_3_41_port, INPUT(215) => 
                           A_pos_shifted_by1_3_40_port, INPUT(216) => 
                           A_pos_shifted_by1_3_39_port, INPUT(217) => 
                           A_pos_shifted_by1_3_38_port, INPUT(218) => 
                           A_pos_shifted_by1_3_37_port, INPUT(219) => 
                           A_pos_shifted_by1_3_36_port, INPUT(220) => 
                           A_pos_shifted_by1_3_35_port, INPUT(221) => 
                           A_pos_shifted_by1_3_34_port, INPUT(222) => 
                           A_pos_shifted_by1_3_33_port, INPUT(223) => 
                           A_pos_shifted_by1_3_32_port, INPUT(224) => 
                           A_pos_shifted_by1_3_31_port, INPUT(225) => 
                           A_pos_shifted_by1_3_30_port, INPUT(226) => 
                           A_pos_shifted_by1_3_29_port, INPUT(227) => 
                           A_pos_shifted_by1_3_28_port, INPUT(228) => 
                           A_pos_shifted_by1_3_27_port, INPUT(229) => 
                           A_pos_shifted_by1_3_26_port, INPUT(230) => 
                           A_pos_shifted_by1_3_25_port, INPUT(231) => 
                           A_pos_shifted_by1_3_24_port, INPUT(232) => 
                           A_pos_shifted_by1_3_23_port, INPUT(233) => 
                           A_pos_shifted_by1_3_22_port, INPUT(234) => 
                           A_pos_shifted_by1_3_21_port, INPUT(235) => 
                           A_pos_shifted_by1_3_20_port, INPUT(236) => 
                           A_pos_shifted_by1_3_19_port, INPUT(237) => 
                           A_pos_shifted_by1_3_18_port, INPUT(238) => 
                           A_pos_shifted_by1_3_17_port, INPUT(239) => 
                           A_pos_shifted_by1_3_16_port, INPUT(240) => 
                           A_pos_shifted_by1_3_15_port, INPUT(241) => 
                           A_pos_shifted_by1_3_14_port, INPUT(242) => 
                           A_pos_shifted_by1_3_13_port, INPUT(243) => 
                           A_pos_shifted_by1_3_12_port, INPUT(244) => 
                           A_pos_shifted_by1_3_11_port, INPUT(245) => 
                           A_pos_shifted_by1_3_10_port, INPUT(246) => 
                           A_pos_shifted_by1_3_9_port, INPUT(247) => 
                           A_pos_shifted_by1_3_8_port, INPUT(248) => 
                           A_pos_shifted_by1_3_7_port, INPUT(249) => 
                           A_pos_shifted_by1_3_6_port, INPUT(250) => 
                           A_pos_shifted_by1_3_5_port, INPUT(251) => 
                           A_pos_shifted_by1_3_4_port, INPUT(252) => 
                           A_pos_shifted_by1_3_3_port, INPUT(253) => 
                           A_pos_shifted_by1_3_2_port, INPUT(254) => 
                           A_pos_shifted_by1_3_1_port, INPUT(255) => 
                           A_pos_shifted_by1_3_0_port, INPUT(256) => 
                           A_neg_shifted_by1_3_63_port, INPUT(257) => 
                           A_neg_shifted_by1_3_62_port, INPUT(258) => 
                           A_neg_shifted_by1_3_61_port, INPUT(259) => 
                           A_neg_shifted_by1_3_60_port, INPUT(260) => 
                           A_neg_shifted_by1_3_59_port, INPUT(261) => 
                           A_neg_shifted_by1_3_58_port, INPUT(262) => 
                           A_neg_shifted_by1_3_57_port, INPUT(263) => 
                           A_neg_shifted_by1_3_56_port, INPUT(264) => 
                           A_neg_shifted_by1_3_55_port, INPUT(265) => 
                           A_neg_shifted_by1_3_54_port, INPUT(266) => 
                           A_neg_shifted_by1_3_53_port, INPUT(267) => 
                           A_neg_shifted_by1_3_52_port, INPUT(268) => 
                           A_neg_shifted_by1_3_51_port, INPUT(269) => 
                           A_neg_shifted_by1_3_50_port, INPUT(270) => 
                           A_neg_shifted_by1_3_49_port, INPUT(271) => 
                           A_neg_shifted_by1_3_48_port, INPUT(272) => 
                           A_neg_shifted_by1_3_47_port, INPUT(273) => 
                           A_neg_shifted_by1_3_46_port, INPUT(274) => 
                           A_neg_shifted_by1_3_45_port, INPUT(275) => 
                           A_neg_shifted_by1_3_44_port, INPUT(276) => 
                           A_neg_shifted_by1_3_43_port, INPUT(277) => 
                           A_neg_shifted_by1_3_42_port, INPUT(278) => 
                           A_neg_shifted_by1_3_41_port, INPUT(279) => 
                           A_neg_shifted_by1_3_40_port, INPUT(280) => 
                           A_neg_shifted_by1_3_39_port, INPUT(281) => 
                           A_neg_shifted_by1_3_38_port, INPUT(282) => 
                           A_neg_shifted_by1_3_37_port, INPUT(283) => 
                           A_neg_shifted_by1_3_36_port, INPUT(284) => 
                           A_neg_shifted_by1_3_35_port, INPUT(285) => 
                           A_neg_shifted_by1_3_34_port, INPUT(286) => 
                           A_neg_shifted_by1_3_33_port, INPUT(287) => 
                           A_neg_shifted_by1_3_32_port, INPUT(288) => 
                           A_neg_shifted_by1_3_31_port, INPUT(289) => 
                           A_neg_shifted_by1_3_30_port, INPUT(290) => 
                           A_neg_shifted_by1_3_29_port, INPUT(291) => 
                           A_neg_shifted_by1_3_28_port, INPUT(292) => 
                           A_neg_shifted_by1_3_27_port, INPUT(293) => 
                           A_neg_shifted_by1_3_26_port, INPUT(294) => 
                           A_neg_shifted_by1_3_25_port, INPUT(295) => 
                           A_neg_shifted_by1_3_24_port, INPUT(296) => 
                           A_neg_shifted_by1_3_23_port, INPUT(297) => 
                           A_neg_shifted_by1_3_22_port, INPUT(298) => 
                           A_neg_shifted_by1_3_21_port, INPUT(299) => 
                           A_neg_shifted_by1_3_20_port, INPUT(300) => 
                           A_neg_shifted_by1_3_19_port, INPUT(301) => 
                           A_neg_shifted_by1_3_18_port, INPUT(302) => 
                           A_neg_shifted_by1_3_17_port, INPUT(303) => 
                           A_neg_shifted_by1_3_16_port, INPUT(304) => 
                           A_neg_shifted_by1_3_15_port, INPUT(305) => 
                           A_neg_shifted_by1_3_14_port, INPUT(306) => 
                           A_neg_shifted_by1_3_13_port, INPUT(307) => 
                           A_neg_shifted_by1_3_12_port, INPUT(308) => 
                           A_neg_shifted_by1_3_11_port, INPUT(309) => 
                           A_neg_shifted_by1_3_10_port, INPUT(310) => 
                           A_neg_shifted_by1_3_9_port, INPUT(311) => 
                           A_neg_shifted_by1_3_8_port, INPUT(312) => 
                           A_neg_shifted_by1_3_7_port, INPUT(313) => 
                           A_neg_shifted_by1_3_6_port, INPUT(314) => 
                           A_neg_shifted_by1_3_5_port, INPUT(315) => 
                           A_neg_shifted_by1_3_4_port, INPUT(316) => 
                           A_neg_shifted_by1_3_3_port, INPUT(317) => 
                           A_neg_shifted_by1_3_2_port, INPUT(318) => 
                           A_neg_shifted_by1_3_1_port, INPUT(319) => 
                           A_neg_shifted_by1_3_0_port, SEL(0) => 
                           selection_signal_3_2_port, SEL(1) => 
                           selection_signal_3_1_port, SEL(2) => 
                           selection_signal_3_0_port, Y(0) => OUT_MUX_3_63_port
                           , Y(1) => OUT_MUX_3_62_port, Y(2) => 
                           OUT_MUX_3_61_port, Y(3) => OUT_MUX_3_60_port, Y(4) 
                           => OUT_MUX_3_59_port, Y(5) => OUT_MUX_3_58_port, 
                           Y(6) => OUT_MUX_3_57_port, Y(7) => OUT_MUX_3_56_port
                           , Y(8) => OUT_MUX_3_55_port, Y(9) => 
                           OUT_MUX_3_54_port, Y(10) => OUT_MUX_3_53_port, Y(11)
                           => OUT_MUX_3_52_port, Y(12) => OUT_MUX_3_51_port, 
                           Y(13) => OUT_MUX_3_50_port, Y(14) => 
                           OUT_MUX_3_49_port, Y(15) => OUT_MUX_3_48_port, Y(16)
                           => OUT_MUX_3_47_port, Y(17) => OUT_MUX_3_46_port, 
                           Y(18) => OUT_MUX_3_45_port, Y(19) => 
                           OUT_MUX_3_44_port, Y(20) => OUT_MUX_3_43_port, Y(21)
                           => OUT_MUX_3_42_port, Y(22) => OUT_MUX_3_41_port, 
                           Y(23) => OUT_MUX_3_40_port, Y(24) => 
                           OUT_MUX_3_39_port, Y(25) => OUT_MUX_3_38_port, Y(26)
                           => OUT_MUX_3_37_port, Y(27) => OUT_MUX_3_36_port, 
                           Y(28) => OUT_MUX_3_35_port, Y(29) => 
                           OUT_MUX_3_34_port, Y(30) => OUT_MUX_3_33_port, Y(31)
                           => OUT_MUX_3_32_port, Y(32) => OUT_MUX_3_31_port, 
                           Y(33) => OUT_MUX_3_30_port, Y(34) => 
                           OUT_MUX_3_29_port, Y(35) => OUT_MUX_3_28_port, Y(36)
                           => OUT_MUX_3_27_port, Y(37) => OUT_MUX_3_26_port, 
                           Y(38) => OUT_MUX_3_25_port, Y(39) => 
                           OUT_MUX_3_24_port, Y(40) => OUT_MUX_3_23_port, Y(41)
                           => OUT_MUX_3_22_port, Y(42) => OUT_MUX_3_21_port, 
                           Y(43) => OUT_MUX_3_20_port, Y(44) => 
                           OUT_MUX_3_19_port, Y(45) => OUT_MUX_3_18_port, Y(46)
                           => OUT_MUX_3_17_port, Y(47) => OUT_MUX_3_16_port, 
                           Y(48) => OUT_MUX_3_15_port, Y(49) => 
                           OUT_MUX_3_14_port, Y(50) => OUT_MUX_3_13_port, Y(51)
                           => OUT_MUX_3_12_port, Y(52) => OUT_MUX_3_11_port, 
                           Y(53) => OUT_MUX_3_10_port, Y(54) => 
                           OUT_MUX_3_9_port, Y(55) => OUT_MUX_3_8_port, Y(56) 
                           => OUT_MUX_3_7_port, Y(57) => OUT_MUX_3_6_port, 
                           Y(58) => OUT_MUX_3_5_port, Y(59) => OUT_MUX_3_4_port
                           , Y(60) => OUT_MUX_3_3_port, Y(61) => 
                           OUT_MUX_3_2_port, Y(62) => OUT_MUX_3_1_port, Y(63) 
                           => OUT_MUX_3_0_port);
   MUXi_4 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_12 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_3_63_port, INPUT(65) => 
                           A_pos_shifted_by2_3_62_port, INPUT(66) => 
                           A_pos_shifted_by2_3_61_port, INPUT(67) => 
                           A_pos_shifted_by2_3_60_port, INPUT(68) => 
                           A_pos_shifted_by2_3_59_port, INPUT(69) => 
                           A_pos_shifted_by2_3_58_port, INPUT(70) => 
                           A_pos_shifted_by2_3_57_port, INPUT(71) => 
                           A_pos_shifted_by2_3_56_port, INPUT(72) => 
                           A_pos_shifted_by2_3_55_port, INPUT(73) => 
                           A_pos_shifted_by2_3_54_port, INPUT(74) => 
                           A_pos_shifted_by2_3_53_port, INPUT(75) => 
                           A_pos_shifted_by2_3_52_port, INPUT(76) => 
                           A_pos_shifted_by2_3_51_port, INPUT(77) => 
                           A_pos_shifted_by2_3_50_port, INPUT(78) => 
                           A_pos_shifted_by2_3_49_port, INPUT(79) => 
                           A_pos_shifted_by2_3_48_port, INPUT(80) => n239, 
                           INPUT(81) => A_pos_shifted_by2_3_46_port, INPUT(82) 
                           => A_pos_shifted_by2_3_45_port, INPUT(83) => 
                           A_pos_shifted_by2_3_44_port, INPUT(84) => 
                           A_pos_shifted_by2_3_43_port, INPUT(85) => 
                           A_pos_shifted_by2_3_42_port, INPUT(86) => 
                           A_pos_shifted_by2_3_41_port, INPUT(87) => 
                           A_pos_shifted_by2_3_40_port, INPUT(88) => 
                           A_pos_shifted_by2_3_39_port, INPUT(89) => 
                           A_pos_shifted_by2_3_38_port, INPUT(90) => 
                           A_pos_shifted_by2_3_37_port, INPUT(91) => 
                           A_pos_shifted_by2_3_36_port, INPUT(92) => 
                           A_pos_shifted_by2_3_35_port, INPUT(93) => 
                           A_pos_shifted_by2_3_34_port, INPUT(94) => 
                           A_pos_shifted_by2_3_33_port, INPUT(95) => 
                           A_pos_shifted_by2_3_32_port, INPUT(96) => 
                           A_pos_shifted_by2_3_31_port, INPUT(97) => 
                           A_pos_shifted_by2_3_30_port, INPUT(98) => 
                           A_pos_shifted_by2_3_29_port, INPUT(99) => 
                           A_pos_shifted_by2_3_28_port, INPUT(100) => 
                           A_pos_shifted_by2_3_27_port, INPUT(101) => 
                           A_pos_shifted_by2_3_26_port, INPUT(102) => 
                           A_pos_shifted_by2_3_25_port, INPUT(103) => 
                           A_pos_shifted_by2_3_24_port, INPUT(104) => 
                           A_pos_shifted_by2_3_23_port, INPUT(105) => 
                           A_pos_shifted_by2_3_22_port, INPUT(106) => 
                           A_pos_shifted_by2_3_21_port, INPUT(107) => 
                           A_pos_shifted_by2_3_20_port, INPUT(108) => 
                           A_pos_shifted_by2_3_19_port, INPUT(109) => 
                           A_pos_shifted_by2_3_18_port, INPUT(110) => 
                           A_pos_shifted_by2_3_17_port, INPUT(111) => 
                           A_pos_shifted_by2_3_16_port, INPUT(112) => 
                           A_pos_shifted_by2_3_15_port, INPUT(113) => 
                           A_pos_shifted_by2_3_14_port, INPUT(114) => 
                           A_pos_shifted_by2_3_13_port, INPUT(115) => 
                           A_pos_shifted_by2_3_12_port, INPUT(116) => 
                           A_pos_shifted_by2_3_11_port, INPUT(117) => 
                           A_pos_shifted_by2_3_10_port, INPUT(118) => 
                           A_pos_shifted_by2_3_9_port, INPUT(119) => 
                           A_pos_shifted_by2_3_8_port, INPUT(120) => 
                           A_pos_shifted_by2_3_7_port, INPUT(121) => 
                           A_pos_shifted_by2_3_6_port, INPUT(122) => 
                           A_pos_shifted_by2_3_5_port, INPUT(123) => 
                           A_pos_shifted_by2_3_4_port, INPUT(124) => 
                           A_pos_shifted_by2_3_3_port, INPUT(125) => 
                           A_pos_shifted_by2_3_2_port, INPUT(126) => 
                           A_pos_shifted_by2_3_1_port, INPUT(127) => 
                           A_pos_shifted_by2_3_0_port, INPUT(128) => 
                           A_neg_shifted_by2_3_63_port, INPUT(129) => 
                           A_neg_shifted_by2_3_62_port, INPUT(130) => 
                           A_neg_shifted_by2_3_61_port, INPUT(131) => 
                           A_neg_shifted_by2_3_60_port, INPUT(132) => 
                           A_neg_shifted_by2_3_59_port, INPUT(133) => 
                           A_neg_shifted_by2_3_58_port, INPUT(134) => 
                           A_neg_shifted_by2_3_57_port, INPUT(135) => 
                           A_neg_shifted_by2_3_56_port, INPUT(136) => 
                           A_neg_shifted_by2_3_55_port, INPUT(137) => 
                           A_neg_shifted_by2_3_54_port, INPUT(138) => 
                           A_neg_shifted_by2_3_53_port, INPUT(139) => 
                           A_neg_shifted_by2_3_52_port, INPUT(140) => 
                           A_neg_shifted_by2_3_51_port, INPUT(141) => 
                           A_neg_shifted_by2_3_50_port, INPUT(142) => 
                           A_neg_shifted_by2_3_49_port, INPUT(143) => 
                           A_neg_shifted_by2_3_48_port, INPUT(144) => n205, 
                           INPUT(145) => A_neg_shifted_by2_3_46_port, 
                           INPUT(146) => A_neg_shifted_by2_3_45_port, 
                           INPUT(147) => A_neg_shifted_by2_3_44_port, 
                           INPUT(148) => A_neg_shifted_by2_3_43_port, 
                           INPUT(149) => A_neg_shifted_by2_3_42_port, 
                           INPUT(150) => A_neg_shifted_by2_3_41_port, 
                           INPUT(151) => A_neg_shifted_by2_3_40_port, 
                           INPUT(152) => A_neg_shifted_by2_3_39_port, 
                           INPUT(153) => A_neg_shifted_by2_3_38_port, 
                           INPUT(154) => A_neg_shifted_by2_3_37_port, 
                           INPUT(155) => A_neg_shifted_by2_3_36_port, 
                           INPUT(156) => A_neg_shifted_by2_3_35_port, 
                           INPUT(157) => A_neg_shifted_by2_3_34_port, 
                           INPUT(158) => A_neg_shifted_by2_3_33_port, 
                           INPUT(159) => A_neg_shifted_by2_3_32_port, 
                           INPUT(160) => A_neg_shifted_by2_3_31_port, 
                           INPUT(161) => A_neg_shifted_by2_3_30_port, 
                           INPUT(162) => A_neg_shifted_by2_3_29_port, 
                           INPUT(163) => A_neg_shifted_by2_3_28_port, 
                           INPUT(164) => A_neg_shifted_by2_3_27_port, 
                           INPUT(165) => A_neg_shifted_by2_3_26_port, 
                           INPUT(166) => A_neg_shifted_by2_3_25_port, 
                           INPUT(167) => A_neg_shifted_by2_3_24_port, 
                           INPUT(168) => A_neg_shifted_by2_3_23_port, 
                           INPUT(169) => A_neg_shifted_by2_3_22_port, 
                           INPUT(170) => A_neg_shifted_by2_3_21_port, 
                           INPUT(171) => A_neg_shifted_by2_3_20_port, 
                           INPUT(172) => A_neg_shifted_by2_3_19_port, 
                           INPUT(173) => A_neg_shifted_by2_3_18_port, 
                           INPUT(174) => A_neg_shifted_by2_3_17_port, 
                           INPUT(175) => A_neg_shifted_by2_3_16_port, 
                           INPUT(176) => A_neg_shifted_by2_3_15_port, 
                           INPUT(177) => A_neg_shifted_by2_3_14_port, 
                           INPUT(178) => A_neg_shifted_by2_3_13_port, 
                           INPUT(179) => A_neg_shifted_by2_3_12_port, 
                           INPUT(180) => A_neg_shifted_by2_3_11_port, 
                           INPUT(181) => A_neg_shifted_by2_3_10_port, 
                           INPUT(182) => A_neg_shifted_by2_3_9_port, INPUT(183)
                           => A_neg_shifted_by2_3_8_port, INPUT(184) => 
                           A_neg_shifted_by2_3_7_port, INPUT(185) => 
                           A_neg_shifted_by2_3_6_port, INPUT(186) => 
                           A_neg_shifted_by2_3_5_port, INPUT(187) => 
                           A_neg_shifted_by2_3_4_port, INPUT(188) => 
                           A_neg_shifted_by2_3_3_port, INPUT(189) => 
                           A_neg_shifted_by2_3_2_port, INPUT(190) => 
                           A_neg_shifted_by2_3_1_port, INPUT(191) => 
                           A_neg_shifted_by2_3_0_port, INPUT(192) => 
                           A_pos_shifted_by1_4_63_port, INPUT(193) => 
                           A_pos_shifted_by1_4_62_port, INPUT(194) => 
                           A_pos_shifted_by1_4_61_port, INPUT(195) => 
                           A_pos_shifted_by1_4_60_port, INPUT(196) => 
                           A_pos_shifted_by1_4_59_port, INPUT(197) => 
                           A_pos_shifted_by1_4_58_port, INPUT(198) => 
                           A_pos_shifted_by1_4_57_port, INPUT(199) => 
                           A_pos_shifted_by1_4_56_port, INPUT(200) => 
                           A_pos_shifted_by1_4_55_port, INPUT(201) => 
                           A_pos_shifted_by1_4_54_port, INPUT(202) => 
                           A_pos_shifted_by1_4_53_port, INPUT(203) => 
                           A_pos_shifted_by1_4_52_port, INPUT(204) => 
                           A_pos_shifted_by1_4_51_port, INPUT(205) => 
                           A_pos_shifted_by1_4_50_port, INPUT(206) => 
                           A_pos_shifted_by1_4_49_port, INPUT(207) => 
                           A_pos_shifted_by1_4_48_port, INPUT(208) => 
                           A_pos_shifted_by1_4_47_port, INPUT(209) => 
                           A_pos_shifted_by1_4_46_port, INPUT(210) => 
                           A_pos_shifted_by1_4_45_port, INPUT(211) => 
                           A_pos_shifted_by1_4_44_port, INPUT(212) => 
                           A_pos_shifted_by1_4_43_port, INPUT(213) => 
                           A_pos_shifted_by1_4_42_port, INPUT(214) => 
                           A_pos_shifted_by1_4_41_port, INPUT(215) => 
                           A_pos_shifted_by1_4_40_port, INPUT(216) => 
                           A_pos_shifted_by1_4_39_port, INPUT(217) => 
                           A_pos_shifted_by1_4_38_port, INPUT(218) => 
                           A_pos_shifted_by1_4_37_port, INPUT(219) => 
                           A_pos_shifted_by1_4_36_port, INPUT(220) => 
                           A_pos_shifted_by1_4_35_port, INPUT(221) => 
                           A_pos_shifted_by1_4_34_port, INPUT(222) => 
                           A_pos_shifted_by1_4_33_port, INPUT(223) => 
                           A_pos_shifted_by1_4_32_port, INPUT(224) => 
                           A_pos_shifted_by1_4_31_port, INPUT(225) => 
                           A_pos_shifted_by1_4_30_port, INPUT(226) => 
                           A_pos_shifted_by1_4_29_port, INPUT(227) => 
                           A_pos_shifted_by1_4_28_port, INPUT(228) => 
                           A_pos_shifted_by1_4_27_port, INPUT(229) => 
                           A_pos_shifted_by1_4_26_port, INPUT(230) => 
                           A_pos_shifted_by1_4_25_port, INPUT(231) => 
                           A_pos_shifted_by1_4_24_port, INPUT(232) => 
                           A_pos_shifted_by1_4_23_port, INPUT(233) => 
                           A_pos_shifted_by1_4_22_port, INPUT(234) => 
                           A_pos_shifted_by1_4_21_port, INPUT(235) => 
                           A_pos_shifted_by1_4_20_port, INPUT(236) => 
                           A_pos_shifted_by1_4_19_port, INPUT(237) => 
                           A_pos_shifted_by1_4_18_port, INPUT(238) => 
                           A_pos_shifted_by1_4_17_port, INPUT(239) => 
                           A_pos_shifted_by1_4_16_port, INPUT(240) => 
                           A_pos_shifted_by1_4_15_port, INPUT(241) => 
                           A_pos_shifted_by1_4_14_port, INPUT(242) => 
                           A_pos_shifted_by1_4_13_port, INPUT(243) => 
                           A_pos_shifted_by1_4_12_port, INPUT(244) => 
                           A_pos_shifted_by1_4_11_port, INPUT(245) => 
                           A_pos_shifted_by1_4_10_port, INPUT(246) => 
                           A_pos_shifted_by1_4_9_port, INPUT(247) => 
                           A_pos_shifted_by1_4_8_port, INPUT(248) => 
                           A_pos_shifted_by1_4_7_port, INPUT(249) => 
                           A_pos_shifted_by1_4_6_port, INPUT(250) => 
                           A_pos_shifted_by1_4_5_port, INPUT(251) => 
                           A_pos_shifted_by1_4_4_port, INPUT(252) => 
                           A_pos_shifted_by1_4_3_port, INPUT(253) => 
                           A_pos_shifted_by1_4_2_port, INPUT(254) => 
                           A_pos_shifted_by1_4_1_port, INPUT(255) => 
                           A_pos_shifted_by1_4_0_port, INPUT(256) => 
                           A_neg_shifted_by1_4_63_port, INPUT(257) => 
                           A_neg_shifted_by1_4_62_port, INPUT(258) => 
                           A_neg_shifted_by1_4_61_port, INPUT(259) => 
                           A_neg_shifted_by1_4_60_port, INPUT(260) => 
                           A_neg_shifted_by1_4_59_port, INPUT(261) => 
                           A_neg_shifted_by1_4_58_port, INPUT(262) => 
                           A_neg_shifted_by1_4_57_port, INPUT(263) => 
                           A_neg_shifted_by1_4_56_port, INPUT(264) => 
                           A_neg_shifted_by1_4_55_port, INPUT(265) => 
                           A_neg_shifted_by1_4_54_port, INPUT(266) => 
                           A_neg_shifted_by1_4_53_port, INPUT(267) => 
                           A_neg_shifted_by1_4_52_port, INPUT(268) => 
                           A_neg_shifted_by1_4_51_port, INPUT(269) => 
                           A_neg_shifted_by1_4_50_port, INPUT(270) => 
                           A_neg_shifted_by1_4_49_port, INPUT(271) => 
                           A_neg_shifted_by1_4_48_port, INPUT(272) => 
                           A_neg_shifted_by1_4_47_port, INPUT(273) => 
                           A_neg_shifted_by1_4_46_port, INPUT(274) => 
                           A_neg_shifted_by1_4_45_port, INPUT(275) => 
                           A_neg_shifted_by1_4_44_port, INPUT(276) => 
                           A_neg_shifted_by1_4_43_port, INPUT(277) => 
                           A_neg_shifted_by1_4_42_port, INPUT(278) => 
                           A_neg_shifted_by1_4_41_port, INPUT(279) => 
                           A_neg_shifted_by1_4_40_port, INPUT(280) => 
                           A_neg_shifted_by1_4_39_port, INPUT(281) => 
                           A_neg_shifted_by1_4_38_port, INPUT(282) => 
                           A_neg_shifted_by1_4_37_port, INPUT(283) => 
                           A_neg_shifted_by1_4_36_port, INPUT(284) => 
                           A_neg_shifted_by1_4_35_port, INPUT(285) => 
                           A_neg_shifted_by1_4_34_port, INPUT(286) => 
                           A_neg_shifted_by1_4_33_port, INPUT(287) => 
                           A_neg_shifted_by1_4_32_port, INPUT(288) => 
                           A_neg_shifted_by1_4_31_port, INPUT(289) => 
                           A_neg_shifted_by1_4_30_port, INPUT(290) => 
                           A_neg_shifted_by1_4_29_port, INPUT(291) => 
                           A_neg_shifted_by1_4_28_port, INPUT(292) => 
                           A_neg_shifted_by1_4_27_port, INPUT(293) => 
                           A_neg_shifted_by1_4_26_port, INPUT(294) => 
                           A_neg_shifted_by1_4_25_port, INPUT(295) => 
                           A_neg_shifted_by1_4_24_port, INPUT(296) => 
                           A_neg_shifted_by1_4_23_port, INPUT(297) => 
                           A_neg_shifted_by1_4_22_port, INPUT(298) => 
                           A_neg_shifted_by1_4_21_port, INPUT(299) => 
                           A_neg_shifted_by1_4_20_port, INPUT(300) => 
                           A_neg_shifted_by1_4_19_port, INPUT(301) => 
                           A_neg_shifted_by1_4_18_port, INPUT(302) => 
                           A_neg_shifted_by1_4_17_port, INPUT(303) => 
                           A_neg_shifted_by1_4_16_port, INPUT(304) => 
                           A_neg_shifted_by1_4_15_port, INPUT(305) => 
                           A_neg_shifted_by1_4_14_port, INPUT(306) => 
                           A_neg_shifted_by1_4_13_port, INPUT(307) => 
                           A_neg_shifted_by1_4_12_port, INPUT(308) => 
                           A_neg_shifted_by1_4_11_port, INPUT(309) => 
                           A_neg_shifted_by1_4_10_port, INPUT(310) => 
                           A_neg_shifted_by1_4_9_port, INPUT(311) => 
                           A_neg_shifted_by1_4_8_port, INPUT(312) => 
                           A_neg_shifted_by1_4_7_port, INPUT(313) => 
                           A_neg_shifted_by1_4_6_port, INPUT(314) => 
                           A_neg_shifted_by1_4_5_port, INPUT(315) => 
                           A_neg_shifted_by1_4_4_port, INPUT(316) => 
                           A_neg_shifted_by1_4_3_port, INPUT(317) => 
                           A_neg_shifted_by1_4_2_port, INPUT(318) => 
                           A_neg_shifted_by1_4_1_port, INPUT(319) => 
                           A_neg_shifted_by1_4_0_port, SEL(0) => 
                           selection_signal_4_2_port, SEL(1) => 
                           selection_signal_4_1_port, SEL(2) => 
                           selection_signal_4_0_port, Y(0) => OUT_MUX_4_63_port
                           , Y(1) => OUT_MUX_4_62_port, Y(2) => 
                           OUT_MUX_4_61_port, Y(3) => OUT_MUX_4_60_port, Y(4) 
                           => OUT_MUX_4_59_port, Y(5) => OUT_MUX_4_58_port, 
                           Y(6) => OUT_MUX_4_57_port, Y(7) => OUT_MUX_4_56_port
                           , Y(8) => OUT_MUX_4_55_port, Y(9) => 
                           OUT_MUX_4_54_port, Y(10) => OUT_MUX_4_53_port, Y(11)
                           => OUT_MUX_4_52_port, Y(12) => OUT_MUX_4_51_port, 
                           Y(13) => OUT_MUX_4_50_port, Y(14) => 
                           OUT_MUX_4_49_port, Y(15) => OUT_MUX_4_48_port, Y(16)
                           => OUT_MUX_4_47_port, Y(17) => OUT_MUX_4_46_port, 
                           Y(18) => OUT_MUX_4_45_port, Y(19) => 
                           OUT_MUX_4_44_port, Y(20) => OUT_MUX_4_43_port, Y(21)
                           => OUT_MUX_4_42_port, Y(22) => OUT_MUX_4_41_port, 
                           Y(23) => OUT_MUX_4_40_port, Y(24) => 
                           OUT_MUX_4_39_port, Y(25) => OUT_MUX_4_38_port, Y(26)
                           => OUT_MUX_4_37_port, Y(27) => OUT_MUX_4_36_port, 
                           Y(28) => OUT_MUX_4_35_port, Y(29) => 
                           OUT_MUX_4_34_port, Y(30) => OUT_MUX_4_33_port, Y(31)
                           => OUT_MUX_4_32_port, Y(32) => OUT_MUX_4_31_port, 
                           Y(33) => OUT_MUX_4_30_port, Y(34) => 
                           OUT_MUX_4_29_port, Y(35) => OUT_MUX_4_28_port, Y(36)
                           => OUT_MUX_4_27_port, Y(37) => OUT_MUX_4_26_port, 
                           Y(38) => OUT_MUX_4_25_port, Y(39) => 
                           OUT_MUX_4_24_port, Y(40) => OUT_MUX_4_23_port, Y(41)
                           => OUT_MUX_4_22_port, Y(42) => OUT_MUX_4_21_port, 
                           Y(43) => OUT_MUX_4_20_port, Y(44) => 
                           OUT_MUX_4_19_port, Y(45) => OUT_MUX_4_18_port, Y(46)
                           => OUT_MUX_4_17_port, Y(47) => OUT_MUX_4_16_port, 
                           Y(48) => OUT_MUX_4_15_port, Y(49) => 
                           OUT_MUX_4_14_port, Y(50) => OUT_MUX_4_13_port, Y(51)
                           => OUT_MUX_4_12_port, Y(52) => OUT_MUX_4_11_port, 
                           Y(53) => OUT_MUX_4_10_port, Y(54) => 
                           OUT_MUX_4_9_port, Y(55) => OUT_MUX_4_8_port, Y(56) 
                           => OUT_MUX_4_7_port, Y(57) => OUT_MUX_4_6_port, 
                           Y(58) => OUT_MUX_4_5_port, Y(59) => OUT_MUX_4_4_port
                           , Y(60) => OUT_MUX_4_3_port, Y(61) => 
                           OUT_MUX_4_2_port, Y(62) => OUT_MUX_4_1_port, Y(63) 
                           => OUT_MUX_4_0_port);
   MUXi_5 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_11 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_4_63_port, INPUT(65) => 
                           A_pos_shifted_by2_4_62_port, INPUT(66) => 
                           A_pos_shifted_by2_4_61_port, INPUT(67) => 
                           A_pos_shifted_by2_4_60_port, INPUT(68) => 
                           A_pos_shifted_by2_4_59_port, INPUT(69) => 
                           A_pos_shifted_by2_4_58_port, INPUT(70) => 
                           A_pos_shifted_by2_4_57_port, INPUT(71) => 
                           A_pos_shifted_by2_4_56_port, INPUT(72) => 
                           A_pos_shifted_by2_4_55_port, INPUT(73) => 
                           A_pos_shifted_by2_4_54_port, INPUT(74) => 
                           A_pos_shifted_by2_4_53_port, INPUT(75) => 
                           A_pos_shifted_by2_4_52_port, INPUT(76) => 
                           A_pos_shifted_by2_4_51_port, INPUT(77) => 
                           A_pos_shifted_by2_4_50_port, INPUT(78) => 
                           A_pos_shifted_by2_4_49_port, INPUT(79) => 
                           A_pos_shifted_by2_4_48_port, INPUT(80) => n238, 
                           INPUT(81) => A_pos_shifted_by2_4_46_port, INPUT(82) 
                           => A_pos_shifted_by2_4_45_port, INPUT(83) => 
                           A_pos_shifted_by2_4_44_port, INPUT(84) => 
                           A_pos_shifted_by2_4_43_port, INPUT(85) => 
                           A_pos_shifted_by2_4_42_port, INPUT(86) => 
                           A_pos_shifted_by2_4_41_port, INPUT(87) => 
                           A_pos_shifted_by2_4_40_port, INPUT(88) => 
                           A_pos_shifted_by2_4_39_port, INPUT(89) => 
                           A_pos_shifted_by2_4_38_port, INPUT(90) => 
                           A_pos_shifted_by2_4_37_port, INPUT(91) => 
                           A_pos_shifted_by2_4_36_port, INPUT(92) => 
                           A_pos_shifted_by2_4_35_port, INPUT(93) => 
                           A_pos_shifted_by2_4_34_port, INPUT(94) => 
                           A_pos_shifted_by2_4_33_port, INPUT(95) => 
                           A_pos_shifted_by2_4_32_port, INPUT(96) => 
                           A_pos_shifted_by2_4_31_port, INPUT(97) => 
                           A_pos_shifted_by2_4_30_port, INPUT(98) => 
                           A_pos_shifted_by2_4_29_port, INPUT(99) => 
                           A_pos_shifted_by2_4_28_port, INPUT(100) => 
                           A_pos_shifted_by2_4_27_port, INPUT(101) => 
                           A_pos_shifted_by2_4_26_port, INPUT(102) => 
                           A_pos_shifted_by2_4_25_port, INPUT(103) => 
                           A_pos_shifted_by2_4_24_port, INPUT(104) => 
                           A_pos_shifted_by2_4_23_port, INPUT(105) => 
                           A_pos_shifted_by2_4_22_port, INPUT(106) => 
                           A_pos_shifted_by2_4_21_port, INPUT(107) => 
                           A_pos_shifted_by2_4_20_port, INPUT(108) => 
                           A_pos_shifted_by2_4_19_port, INPUT(109) => 
                           A_pos_shifted_by2_4_18_port, INPUT(110) => 
                           A_pos_shifted_by2_4_17_port, INPUT(111) => 
                           A_pos_shifted_by2_4_16_port, INPUT(112) => 
                           A_pos_shifted_by2_4_15_port, INPUT(113) => 
                           A_pos_shifted_by2_4_14_port, INPUT(114) => 
                           A_pos_shifted_by2_4_13_port, INPUT(115) => 
                           A_pos_shifted_by2_4_12_port, INPUT(116) => 
                           A_pos_shifted_by2_4_11_port, INPUT(117) => 
                           A_pos_shifted_by2_4_10_port, INPUT(118) => 
                           A_pos_shifted_by2_4_9_port, INPUT(119) => 
                           A_pos_shifted_by2_4_8_port, INPUT(120) => 
                           A_pos_shifted_by2_4_7_port, INPUT(121) => 
                           A_pos_shifted_by2_4_6_port, INPUT(122) => 
                           A_pos_shifted_by2_4_5_port, INPUT(123) => 
                           A_pos_shifted_by2_4_4_port, INPUT(124) => 
                           A_pos_shifted_by2_4_3_port, INPUT(125) => 
                           A_pos_shifted_by2_4_2_port, INPUT(126) => 
                           A_pos_shifted_by2_4_1_port, INPUT(127) => 
                           A_pos_shifted_by2_4_0_port, INPUT(128) => 
                           A_neg_shifted_by2_4_63_port, INPUT(129) => 
                           A_neg_shifted_by2_4_62_port, INPUT(130) => 
                           A_neg_shifted_by2_4_61_port, INPUT(131) => 
                           A_neg_shifted_by2_4_60_port, INPUT(132) => 
                           A_neg_shifted_by2_4_59_port, INPUT(133) => 
                           A_neg_shifted_by2_4_58_port, INPUT(134) => 
                           A_neg_shifted_by2_4_57_port, INPUT(135) => 
                           A_neg_shifted_by2_4_56_port, INPUT(136) => 
                           A_neg_shifted_by2_4_55_port, INPUT(137) => 
                           A_neg_shifted_by2_4_54_port, INPUT(138) => 
                           A_neg_shifted_by2_4_53_port, INPUT(139) => 
                           A_neg_shifted_by2_4_52_port, INPUT(140) => 
                           A_neg_shifted_by2_4_51_port, INPUT(141) => 
                           A_neg_shifted_by2_4_50_port, INPUT(142) => 
                           A_neg_shifted_by2_4_49_port, INPUT(143) => 
                           A_neg_shifted_by2_4_48_port, INPUT(144) => n204, 
                           INPUT(145) => A_neg_shifted_by2_4_46_port, 
                           INPUT(146) => A_neg_shifted_by2_4_45_port, 
                           INPUT(147) => A_neg_shifted_by2_4_44_port, 
                           INPUT(148) => A_neg_shifted_by2_4_43_port, 
                           INPUT(149) => A_neg_shifted_by2_4_42_port, 
                           INPUT(150) => A_neg_shifted_by2_4_41_port, 
                           INPUT(151) => A_neg_shifted_by2_4_40_port, 
                           INPUT(152) => A_neg_shifted_by2_4_39_port, 
                           INPUT(153) => A_neg_shifted_by2_4_38_port, 
                           INPUT(154) => A_neg_shifted_by2_4_37_port, 
                           INPUT(155) => A_neg_shifted_by2_4_36_port, 
                           INPUT(156) => A_neg_shifted_by2_4_35_port, 
                           INPUT(157) => A_neg_shifted_by2_4_34_port, 
                           INPUT(158) => A_neg_shifted_by2_4_33_port, 
                           INPUT(159) => A_neg_shifted_by2_4_32_port, 
                           INPUT(160) => A_neg_shifted_by2_4_31_port, 
                           INPUT(161) => A_neg_shifted_by2_4_30_port, 
                           INPUT(162) => A_neg_shifted_by2_4_29_port, 
                           INPUT(163) => A_neg_shifted_by2_4_28_port, 
                           INPUT(164) => A_neg_shifted_by2_4_27_port, 
                           INPUT(165) => A_neg_shifted_by2_4_26_port, 
                           INPUT(166) => A_neg_shifted_by2_4_25_port, 
                           INPUT(167) => A_neg_shifted_by2_4_24_port, 
                           INPUT(168) => A_neg_shifted_by2_4_23_port, 
                           INPUT(169) => A_neg_shifted_by2_4_22_port, 
                           INPUT(170) => A_neg_shifted_by2_4_21_port, 
                           INPUT(171) => A_neg_shifted_by2_4_20_port, 
                           INPUT(172) => A_neg_shifted_by2_4_19_port, 
                           INPUT(173) => A_neg_shifted_by2_4_18_port, 
                           INPUT(174) => A_neg_shifted_by2_4_17_port, 
                           INPUT(175) => A_neg_shifted_by2_4_16_port, 
                           INPUT(176) => A_neg_shifted_by2_4_15_port, 
                           INPUT(177) => A_neg_shifted_by2_4_14_port, 
                           INPUT(178) => A_neg_shifted_by2_4_13_port, 
                           INPUT(179) => A_neg_shifted_by2_4_12_port, 
                           INPUT(180) => A_neg_shifted_by2_4_11_port, 
                           INPUT(181) => A_neg_shifted_by2_4_10_port, 
                           INPUT(182) => A_neg_shifted_by2_4_9_port, INPUT(183)
                           => A_neg_shifted_by2_4_8_port, INPUT(184) => 
                           A_neg_shifted_by2_4_7_port, INPUT(185) => 
                           A_neg_shifted_by2_4_6_port, INPUT(186) => 
                           A_neg_shifted_by2_4_5_port, INPUT(187) => 
                           A_neg_shifted_by2_4_4_port, INPUT(188) => 
                           A_neg_shifted_by2_4_3_port, INPUT(189) => 
                           A_neg_shifted_by2_4_2_port, INPUT(190) => 
                           A_neg_shifted_by2_4_1_port, INPUT(191) => 
                           A_neg_shifted_by2_4_0_port, INPUT(192) => 
                           A_pos_shifted_by1_5_63_port, INPUT(193) => 
                           A_pos_shifted_by1_5_62_port, INPUT(194) => 
                           A_pos_shifted_by1_5_61_port, INPUT(195) => 
                           A_pos_shifted_by1_5_60_port, INPUT(196) => 
                           A_pos_shifted_by1_5_59_port, INPUT(197) => 
                           A_pos_shifted_by1_5_58_port, INPUT(198) => 
                           A_pos_shifted_by1_5_57_port, INPUT(199) => 
                           A_pos_shifted_by1_5_56_port, INPUT(200) => 
                           A_pos_shifted_by1_5_55_port, INPUT(201) => 
                           A_pos_shifted_by1_5_54_port, INPUT(202) => 
                           A_pos_shifted_by1_5_53_port, INPUT(203) => 
                           A_pos_shifted_by1_5_52_port, INPUT(204) => 
                           A_pos_shifted_by1_5_51_port, INPUT(205) => 
                           A_pos_shifted_by1_5_50_port, INPUT(206) => 
                           A_pos_shifted_by1_5_49_port, INPUT(207) => 
                           A_pos_shifted_by1_5_48_port, INPUT(208) => 
                           A_pos_shifted_by1_5_47_port, INPUT(209) => 
                           A_pos_shifted_by1_5_46_port, INPUT(210) => 
                           A_pos_shifted_by1_5_45_port, INPUT(211) => 
                           A_pos_shifted_by1_5_44_port, INPUT(212) => 
                           A_pos_shifted_by1_5_43_port, INPUT(213) => 
                           A_pos_shifted_by1_5_42_port, INPUT(214) => 
                           A_pos_shifted_by1_5_41_port, INPUT(215) => 
                           A_pos_shifted_by1_5_40_port, INPUT(216) => 
                           A_pos_shifted_by1_5_39_port, INPUT(217) => 
                           A_pos_shifted_by1_5_38_port, INPUT(218) => 
                           A_pos_shifted_by1_5_37_port, INPUT(219) => 
                           A_pos_shifted_by1_5_36_port, INPUT(220) => 
                           A_pos_shifted_by1_5_35_port, INPUT(221) => 
                           A_pos_shifted_by1_5_34_port, INPUT(222) => 
                           A_pos_shifted_by1_5_33_port, INPUT(223) => 
                           A_pos_shifted_by1_5_32_port, INPUT(224) => 
                           A_pos_shifted_by1_5_31_port, INPUT(225) => 
                           A_pos_shifted_by1_5_30_port, INPUT(226) => 
                           A_pos_shifted_by1_5_29_port, INPUT(227) => 
                           A_pos_shifted_by1_5_28_port, INPUT(228) => 
                           A_pos_shifted_by1_5_27_port, INPUT(229) => 
                           A_pos_shifted_by1_5_26_port, INPUT(230) => 
                           A_pos_shifted_by1_5_25_port, INPUT(231) => 
                           A_pos_shifted_by1_5_24_port, INPUT(232) => 
                           A_pos_shifted_by1_5_23_port, INPUT(233) => 
                           A_pos_shifted_by1_5_22_port, INPUT(234) => 
                           A_pos_shifted_by1_5_21_port, INPUT(235) => 
                           A_pos_shifted_by1_5_20_port, INPUT(236) => 
                           A_pos_shifted_by1_5_19_port, INPUT(237) => 
                           A_pos_shifted_by1_5_18_port, INPUT(238) => 
                           A_pos_shifted_by1_5_17_port, INPUT(239) => 
                           A_pos_shifted_by1_5_16_port, INPUT(240) => 
                           A_pos_shifted_by1_5_15_port, INPUT(241) => 
                           A_pos_shifted_by1_5_14_port, INPUT(242) => 
                           A_pos_shifted_by1_5_13_port, INPUT(243) => 
                           A_pos_shifted_by1_5_12_port, INPUT(244) => 
                           A_pos_shifted_by1_5_11_port, INPUT(245) => 
                           A_pos_shifted_by1_5_10_port, INPUT(246) => 
                           A_pos_shifted_by1_5_9_port, INPUT(247) => 
                           A_pos_shifted_by1_5_8_port, INPUT(248) => 
                           A_pos_shifted_by1_5_7_port, INPUT(249) => 
                           A_pos_shifted_by1_5_6_port, INPUT(250) => 
                           A_pos_shifted_by1_5_5_port, INPUT(251) => 
                           A_pos_shifted_by1_5_4_port, INPUT(252) => 
                           A_pos_shifted_by1_5_3_port, INPUT(253) => 
                           A_pos_shifted_by1_5_2_port, INPUT(254) => 
                           A_pos_shifted_by1_5_1_port, INPUT(255) => 
                           A_pos_shifted_by1_5_0_port, INPUT(256) => 
                           A_neg_shifted_by1_5_63_port, INPUT(257) => 
                           A_neg_shifted_by1_5_62_port, INPUT(258) => 
                           A_neg_shifted_by1_5_61_port, INPUT(259) => 
                           A_neg_shifted_by1_5_60_port, INPUT(260) => 
                           A_neg_shifted_by1_5_59_port, INPUT(261) => 
                           A_neg_shifted_by1_5_58_port, INPUT(262) => 
                           A_neg_shifted_by1_5_57_port, INPUT(263) => 
                           A_neg_shifted_by1_5_56_port, INPUT(264) => 
                           A_neg_shifted_by1_5_55_port, INPUT(265) => 
                           A_neg_shifted_by1_5_54_port, INPUT(266) => 
                           A_neg_shifted_by1_5_53_port, INPUT(267) => 
                           A_neg_shifted_by1_5_52_port, INPUT(268) => 
                           A_neg_shifted_by1_5_51_port, INPUT(269) => 
                           A_neg_shifted_by1_5_50_port, INPUT(270) => 
                           A_neg_shifted_by1_5_49_port, INPUT(271) => 
                           A_neg_shifted_by1_5_48_port, INPUT(272) => 
                           A_neg_shifted_by1_5_47_port, INPUT(273) => 
                           A_neg_shifted_by1_5_46_port, INPUT(274) => 
                           A_neg_shifted_by1_5_45_port, INPUT(275) => 
                           A_neg_shifted_by1_5_44_port, INPUT(276) => 
                           A_neg_shifted_by1_5_43_port, INPUT(277) => 
                           A_neg_shifted_by1_5_42_port, INPUT(278) => 
                           A_neg_shifted_by1_5_41_port, INPUT(279) => 
                           A_neg_shifted_by1_5_40_port, INPUT(280) => 
                           A_neg_shifted_by1_5_39_port, INPUT(281) => 
                           A_neg_shifted_by1_5_38_port, INPUT(282) => 
                           A_neg_shifted_by1_5_37_port, INPUT(283) => 
                           A_neg_shifted_by1_5_36_port, INPUT(284) => 
                           A_neg_shifted_by1_5_35_port, INPUT(285) => 
                           A_neg_shifted_by1_5_34_port, INPUT(286) => 
                           A_neg_shifted_by1_5_33_port, INPUT(287) => 
                           A_neg_shifted_by1_5_32_port, INPUT(288) => 
                           A_neg_shifted_by1_5_31_port, INPUT(289) => 
                           A_neg_shifted_by1_5_30_port, INPUT(290) => 
                           A_neg_shifted_by1_5_29_port, INPUT(291) => 
                           A_neg_shifted_by1_5_28_port, INPUT(292) => 
                           A_neg_shifted_by1_5_27_port, INPUT(293) => 
                           A_neg_shifted_by1_5_26_port, INPUT(294) => 
                           A_neg_shifted_by1_5_25_port, INPUT(295) => 
                           A_neg_shifted_by1_5_24_port, INPUT(296) => 
                           A_neg_shifted_by1_5_23_port, INPUT(297) => 
                           A_neg_shifted_by1_5_22_port, INPUT(298) => 
                           A_neg_shifted_by1_5_21_port, INPUT(299) => 
                           A_neg_shifted_by1_5_20_port, INPUT(300) => 
                           A_neg_shifted_by1_5_19_port, INPUT(301) => 
                           A_neg_shifted_by1_5_18_port, INPUT(302) => 
                           A_neg_shifted_by1_5_17_port, INPUT(303) => 
                           A_neg_shifted_by1_5_16_port, INPUT(304) => 
                           A_neg_shifted_by1_5_15_port, INPUT(305) => 
                           A_neg_shifted_by1_5_14_port, INPUT(306) => 
                           A_neg_shifted_by1_5_13_port, INPUT(307) => 
                           A_neg_shifted_by1_5_12_port, INPUT(308) => 
                           A_neg_shifted_by1_5_11_port, INPUT(309) => 
                           A_neg_shifted_by1_5_10_port, INPUT(310) => 
                           A_neg_shifted_by1_5_9_port, INPUT(311) => 
                           A_neg_shifted_by1_5_8_port, INPUT(312) => 
                           A_neg_shifted_by1_5_7_port, INPUT(313) => 
                           A_neg_shifted_by1_5_6_port, INPUT(314) => 
                           A_neg_shifted_by1_5_5_port, INPUT(315) => 
                           A_neg_shifted_by1_5_4_port, INPUT(316) => 
                           A_neg_shifted_by1_5_3_port, INPUT(317) => 
                           A_neg_shifted_by1_5_2_port, INPUT(318) => 
                           A_neg_shifted_by1_5_1_port, INPUT(319) => 
                           A_neg_shifted_by1_5_0_port, SEL(0) => 
                           selection_signal_5_2_port, SEL(1) => 
                           selection_signal_5_1_port, SEL(2) => 
                           selection_signal_5_0_port, Y(0) => OUT_MUX_5_63_port
                           , Y(1) => OUT_MUX_5_62_port, Y(2) => 
                           OUT_MUX_5_61_port, Y(3) => OUT_MUX_5_60_port, Y(4) 
                           => OUT_MUX_5_59_port, Y(5) => OUT_MUX_5_58_port, 
                           Y(6) => OUT_MUX_5_57_port, Y(7) => OUT_MUX_5_56_port
                           , Y(8) => OUT_MUX_5_55_port, Y(9) => 
                           OUT_MUX_5_54_port, Y(10) => OUT_MUX_5_53_port, Y(11)
                           => OUT_MUX_5_52_port, Y(12) => OUT_MUX_5_51_port, 
                           Y(13) => OUT_MUX_5_50_port, Y(14) => 
                           OUT_MUX_5_49_port, Y(15) => OUT_MUX_5_48_port, Y(16)
                           => OUT_MUX_5_47_port, Y(17) => OUT_MUX_5_46_port, 
                           Y(18) => OUT_MUX_5_45_port, Y(19) => 
                           OUT_MUX_5_44_port, Y(20) => OUT_MUX_5_43_port, Y(21)
                           => OUT_MUX_5_42_port, Y(22) => OUT_MUX_5_41_port, 
                           Y(23) => OUT_MUX_5_40_port, Y(24) => 
                           OUT_MUX_5_39_port, Y(25) => OUT_MUX_5_38_port, Y(26)
                           => OUT_MUX_5_37_port, Y(27) => OUT_MUX_5_36_port, 
                           Y(28) => OUT_MUX_5_35_port, Y(29) => 
                           OUT_MUX_5_34_port, Y(30) => OUT_MUX_5_33_port, Y(31)
                           => OUT_MUX_5_32_port, Y(32) => OUT_MUX_5_31_port, 
                           Y(33) => OUT_MUX_5_30_port, Y(34) => 
                           OUT_MUX_5_29_port, Y(35) => OUT_MUX_5_28_port, Y(36)
                           => OUT_MUX_5_27_port, Y(37) => OUT_MUX_5_26_port, 
                           Y(38) => OUT_MUX_5_25_port, Y(39) => 
                           OUT_MUX_5_24_port, Y(40) => OUT_MUX_5_23_port, Y(41)
                           => OUT_MUX_5_22_port, Y(42) => OUT_MUX_5_21_port, 
                           Y(43) => OUT_MUX_5_20_port, Y(44) => 
                           OUT_MUX_5_19_port, Y(45) => OUT_MUX_5_18_port, Y(46)
                           => OUT_MUX_5_17_port, Y(47) => OUT_MUX_5_16_port, 
                           Y(48) => OUT_MUX_5_15_port, Y(49) => 
                           OUT_MUX_5_14_port, Y(50) => OUT_MUX_5_13_port, Y(51)
                           => OUT_MUX_5_12_port, Y(52) => OUT_MUX_5_11_port, 
                           Y(53) => OUT_MUX_5_10_port, Y(54) => 
                           OUT_MUX_5_9_port, Y(55) => OUT_MUX_5_8_port, Y(56) 
                           => OUT_MUX_5_7_port, Y(57) => OUT_MUX_5_6_port, 
                           Y(58) => OUT_MUX_5_5_port, Y(59) => OUT_MUX_5_4_port
                           , Y(60) => OUT_MUX_5_3_port, Y(61) => 
                           OUT_MUX_5_2_port, Y(62) => OUT_MUX_5_1_port, Y(63) 
                           => OUT_MUX_5_0_port);
   MUXi_6 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_10 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_5_63_port, INPUT(65) => 
                           A_pos_shifted_by2_5_62_port, INPUT(66) => 
                           A_pos_shifted_by2_5_61_port, INPUT(67) => 
                           A_pos_shifted_by2_5_60_port, INPUT(68) => 
                           A_pos_shifted_by2_5_59_port, INPUT(69) => 
                           A_pos_shifted_by2_5_58_port, INPUT(70) => 
                           A_pos_shifted_by2_5_57_port, INPUT(71) => 
                           A_pos_shifted_by2_5_56_port, INPUT(72) => 
                           A_pos_shifted_by2_5_55_port, INPUT(73) => 
                           A_pos_shifted_by2_5_54_port, INPUT(74) => 
                           A_pos_shifted_by2_5_53_port, INPUT(75) => 
                           A_pos_shifted_by2_5_52_port, INPUT(76) => 
                           A_pos_shifted_by2_5_51_port, INPUT(77) => 
                           A_pos_shifted_by2_5_50_port, INPUT(78) => 
                           A_pos_shifted_by2_5_49_port, INPUT(79) => 
                           A_pos_shifted_by2_5_48_port, INPUT(80) => n237, 
                           INPUT(81) => A_pos_shifted_by2_5_46_port, INPUT(82) 
                           => A_pos_shifted_by2_5_45_port, INPUT(83) => 
                           A_pos_shifted_by2_5_44_port, INPUT(84) => 
                           A_pos_shifted_by2_5_43_port, INPUT(85) => 
                           A_pos_shifted_by2_5_42_port, INPUT(86) => 
                           A_pos_shifted_by2_5_41_port, INPUT(87) => 
                           A_pos_shifted_by2_5_40_port, INPUT(88) => 
                           A_pos_shifted_by2_5_39_port, INPUT(89) => 
                           A_pos_shifted_by2_5_38_port, INPUT(90) => 
                           A_pos_shifted_by2_5_37_port, INPUT(91) => 
                           A_pos_shifted_by2_5_36_port, INPUT(92) => 
                           A_pos_shifted_by2_5_35_port, INPUT(93) => 
                           A_pos_shifted_by2_5_34_port, INPUT(94) => 
                           A_pos_shifted_by2_5_33_port, INPUT(95) => 
                           A_pos_shifted_by2_5_32_port, INPUT(96) => 
                           A_pos_shifted_by2_5_31_port, INPUT(97) => 
                           A_pos_shifted_by2_5_30_port, INPUT(98) => 
                           A_pos_shifted_by2_5_29_port, INPUT(99) => 
                           A_pos_shifted_by2_5_28_port, INPUT(100) => 
                           A_pos_shifted_by2_5_27_port, INPUT(101) => 
                           A_pos_shifted_by2_5_26_port, INPUT(102) => 
                           A_pos_shifted_by2_5_25_port, INPUT(103) => 
                           A_pos_shifted_by2_5_24_port, INPUT(104) => 
                           A_pos_shifted_by2_5_23_port, INPUT(105) => 
                           A_pos_shifted_by2_5_22_port, INPUT(106) => 
                           A_pos_shifted_by2_5_21_port, INPUT(107) => 
                           A_pos_shifted_by2_5_20_port, INPUT(108) => 
                           A_pos_shifted_by2_5_19_port, INPUT(109) => 
                           A_pos_shifted_by2_5_18_port, INPUT(110) => 
                           A_pos_shifted_by2_5_17_port, INPUT(111) => 
                           A_pos_shifted_by2_5_16_port, INPUT(112) => 
                           A_pos_shifted_by2_5_15_port, INPUT(113) => 
                           A_pos_shifted_by2_5_14_port, INPUT(114) => 
                           A_pos_shifted_by2_5_13_port, INPUT(115) => 
                           A_pos_shifted_by2_5_12_port, INPUT(116) => 
                           A_pos_shifted_by2_5_11_port, INPUT(117) => 
                           A_pos_shifted_by2_5_10_port, INPUT(118) => 
                           A_pos_shifted_by2_5_9_port, INPUT(119) => 
                           A_pos_shifted_by2_5_8_port, INPUT(120) => 
                           A_pos_shifted_by2_5_7_port, INPUT(121) => 
                           A_pos_shifted_by2_5_6_port, INPUT(122) => 
                           A_pos_shifted_by2_5_5_port, INPUT(123) => 
                           A_pos_shifted_by2_5_4_port, INPUT(124) => 
                           A_pos_shifted_by2_5_3_port, INPUT(125) => 
                           A_pos_shifted_by2_5_2_port, INPUT(126) => 
                           A_pos_shifted_by2_5_1_port, INPUT(127) => 
                           A_pos_shifted_by2_5_0_port, INPUT(128) => 
                           A_neg_shifted_by2_5_63_port, INPUT(129) => 
                           A_neg_shifted_by2_5_62_port, INPUT(130) => 
                           A_neg_shifted_by2_5_61_port, INPUT(131) => 
                           A_neg_shifted_by2_5_60_port, INPUT(132) => 
                           A_neg_shifted_by2_5_59_port, INPUT(133) => 
                           A_neg_shifted_by2_5_58_port, INPUT(134) => 
                           A_neg_shifted_by2_5_57_port, INPUT(135) => 
                           A_neg_shifted_by2_5_56_port, INPUT(136) => 
                           A_neg_shifted_by2_5_55_port, INPUT(137) => 
                           A_neg_shifted_by2_5_54_port, INPUT(138) => 
                           A_neg_shifted_by2_5_53_port, INPUT(139) => 
                           A_neg_shifted_by2_5_52_port, INPUT(140) => 
                           A_neg_shifted_by2_5_51_port, INPUT(141) => 
                           A_neg_shifted_by2_5_50_port, INPUT(142) => 
                           A_neg_shifted_by2_5_49_port, INPUT(143) => 
                           A_neg_shifted_by2_5_48_port, INPUT(144) => n203, 
                           INPUT(145) => A_neg_shifted_by2_5_46_port, 
                           INPUT(146) => A_neg_shifted_by2_5_45_port, 
                           INPUT(147) => A_neg_shifted_by2_5_44_port, 
                           INPUT(148) => A_neg_shifted_by2_5_43_port, 
                           INPUT(149) => A_neg_shifted_by2_5_42_port, 
                           INPUT(150) => A_neg_shifted_by2_5_41_port, 
                           INPUT(151) => A_neg_shifted_by2_5_40_port, 
                           INPUT(152) => A_neg_shifted_by2_5_39_port, 
                           INPUT(153) => A_neg_shifted_by2_5_38_port, 
                           INPUT(154) => A_neg_shifted_by2_5_37_port, 
                           INPUT(155) => A_neg_shifted_by2_5_36_port, 
                           INPUT(156) => A_neg_shifted_by2_5_35_port, 
                           INPUT(157) => A_neg_shifted_by2_5_34_port, 
                           INPUT(158) => A_neg_shifted_by2_5_33_port, 
                           INPUT(159) => A_neg_shifted_by2_5_32_port, 
                           INPUT(160) => A_neg_shifted_by2_5_31_port, 
                           INPUT(161) => A_neg_shifted_by2_5_30_port, 
                           INPUT(162) => A_neg_shifted_by2_5_29_port, 
                           INPUT(163) => A_neg_shifted_by2_5_28_port, 
                           INPUT(164) => A_neg_shifted_by2_5_27_port, 
                           INPUT(165) => A_neg_shifted_by2_5_26_port, 
                           INPUT(166) => A_neg_shifted_by2_5_25_port, 
                           INPUT(167) => A_neg_shifted_by2_5_24_port, 
                           INPUT(168) => A_neg_shifted_by2_5_23_port, 
                           INPUT(169) => A_neg_shifted_by2_5_22_port, 
                           INPUT(170) => A_neg_shifted_by2_5_21_port, 
                           INPUT(171) => A_neg_shifted_by2_5_20_port, 
                           INPUT(172) => A_neg_shifted_by2_5_19_port, 
                           INPUT(173) => A_neg_shifted_by2_5_18_port, 
                           INPUT(174) => A_neg_shifted_by2_5_17_port, 
                           INPUT(175) => A_neg_shifted_by2_5_16_port, 
                           INPUT(176) => A_neg_shifted_by2_5_15_port, 
                           INPUT(177) => A_neg_shifted_by2_5_14_port, 
                           INPUT(178) => A_neg_shifted_by2_5_13_port, 
                           INPUT(179) => A_neg_shifted_by2_5_12_port, 
                           INPUT(180) => A_neg_shifted_by2_5_11_port, 
                           INPUT(181) => A_neg_shifted_by2_5_10_port, 
                           INPUT(182) => A_neg_shifted_by2_5_9_port, INPUT(183)
                           => A_neg_shifted_by2_5_8_port, INPUT(184) => 
                           A_neg_shifted_by2_5_7_port, INPUT(185) => 
                           A_neg_shifted_by2_5_6_port, INPUT(186) => 
                           A_neg_shifted_by2_5_5_port, INPUT(187) => 
                           A_neg_shifted_by2_5_4_port, INPUT(188) => 
                           A_neg_shifted_by2_5_3_port, INPUT(189) => 
                           A_neg_shifted_by2_5_2_port, INPUT(190) => 
                           A_neg_shifted_by2_5_1_port, INPUT(191) => 
                           A_neg_shifted_by2_5_0_port, INPUT(192) => 
                           A_pos_shifted_by1_6_63_port, INPUT(193) => 
                           A_pos_shifted_by1_6_62_port, INPUT(194) => 
                           A_pos_shifted_by1_6_61_port, INPUT(195) => 
                           A_pos_shifted_by1_6_60_port, INPUT(196) => 
                           A_pos_shifted_by1_6_59_port, INPUT(197) => 
                           A_pos_shifted_by1_6_58_port, INPUT(198) => 
                           A_pos_shifted_by1_6_57_port, INPUT(199) => 
                           A_pos_shifted_by1_6_56_port, INPUT(200) => 
                           A_pos_shifted_by1_6_55_port, INPUT(201) => 
                           A_pos_shifted_by1_6_54_port, INPUT(202) => 
                           A_pos_shifted_by1_6_53_port, INPUT(203) => 
                           A_pos_shifted_by1_6_52_port, INPUT(204) => 
                           A_pos_shifted_by1_6_51_port, INPUT(205) => 
                           A_pos_shifted_by1_6_50_port, INPUT(206) => 
                           A_pos_shifted_by1_6_49_port, INPUT(207) => 
                           A_pos_shifted_by1_6_48_port, INPUT(208) => 
                           A_pos_shifted_by1_6_47_port, INPUT(209) => 
                           A_pos_shifted_by1_6_46_port, INPUT(210) => 
                           A_pos_shifted_by1_6_45_port, INPUT(211) => 
                           A_pos_shifted_by1_6_44_port, INPUT(212) => 
                           A_pos_shifted_by1_6_43_port, INPUT(213) => 
                           A_pos_shifted_by1_6_42_port, INPUT(214) => 
                           A_pos_shifted_by1_6_41_port, INPUT(215) => 
                           A_pos_shifted_by1_6_40_port, INPUT(216) => 
                           A_pos_shifted_by1_6_39_port, INPUT(217) => 
                           A_pos_shifted_by1_6_38_port, INPUT(218) => 
                           A_pos_shifted_by1_6_37_port, INPUT(219) => 
                           A_pos_shifted_by1_6_36_port, INPUT(220) => 
                           A_pos_shifted_by1_6_35_port, INPUT(221) => 
                           A_pos_shifted_by1_6_34_port, INPUT(222) => 
                           A_pos_shifted_by1_6_33_port, INPUT(223) => 
                           A_pos_shifted_by1_6_32_port, INPUT(224) => 
                           A_pos_shifted_by1_6_31_port, INPUT(225) => 
                           A_pos_shifted_by1_6_30_port, INPUT(226) => 
                           A_pos_shifted_by1_6_29_port, INPUT(227) => 
                           A_pos_shifted_by1_6_28_port, INPUT(228) => 
                           A_pos_shifted_by1_6_27_port, INPUT(229) => 
                           A_pos_shifted_by1_6_26_port, INPUT(230) => 
                           A_pos_shifted_by1_6_25_port, INPUT(231) => 
                           A_pos_shifted_by1_6_24_port, INPUT(232) => 
                           A_pos_shifted_by1_6_23_port, INPUT(233) => 
                           A_pos_shifted_by1_6_22_port, INPUT(234) => 
                           A_pos_shifted_by1_6_21_port, INPUT(235) => 
                           A_pos_shifted_by1_6_20_port, INPUT(236) => 
                           A_pos_shifted_by1_6_19_port, INPUT(237) => 
                           A_pos_shifted_by1_6_18_port, INPUT(238) => 
                           A_pos_shifted_by1_6_17_port, INPUT(239) => 
                           A_pos_shifted_by1_6_16_port, INPUT(240) => 
                           A_pos_shifted_by1_6_15_port, INPUT(241) => 
                           A_pos_shifted_by1_6_14_port, INPUT(242) => 
                           A_pos_shifted_by1_6_13_port, INPUT(243) => 
                           A_pos_shifted_by1_6_12_port, INPUT(244) => 
                           A_pos_shifted_by1_6_11_port, INPUT(245) => 
                           A_pos_shifted_by1_6_10_port, INPUT(246) => 
                           A_pos_shifted_by1_6_9_port, INPUT(247) => 
                           A_pos_shifted_by1_6_8_port, INPUT(248) => 
                           A_pos_shifted_by1_6_7_port, INPUT(249) => 
                           A_pos_shifted_by1_6_6_port, INPUT(250) => 
                           A_pos_shifted_by1_6_5_port, INPUT(251) => 
                           A_pos_shifted_by1_6_4_port, INPUT(252) => 
                           A_pos_shifted_by1_6_3_port, INPUT(253) => 
                           A_pos_shifted_by1_6_2_port, INPUT(254) => 
                           A_pos_shifted_by1_6_1_port, INPUT(255) => 
                           A_pos_shifted_by1_6_0_port, INPUT(256) => 
                           A_neg_shifted_by1_6_63_port, INPUT(257) => 
                           A_neg_shifted_by1_6_62_port, INPUT(258) => 
                           A_neg_shifted_by1_6_61_port, INPUT(259) => 
                           A_neg_shifted_by1_6_60_port, INPUT(260) => 
                           A_neg_shifted_by1_6_59_port, INPUT(261) => 
                           A_neg_shifted_by1_6_58_port, INPUT(262) => 
                           A_neg_shifted_by1_6_57_port, INPUT(263) => 
                           A_neg_shifted_by1_6_56_port, INPUT(264) => 
                           A_neg_shifted_by1_6_55_port, INPUT(265) => 
                           A_neg_shifted_by1_6_54_port, INPUT(266) => 
                           A_neg_shifted_by1_6_53_port, INPUT(267) => 
                           A_neg_shifted_by1_6_52_port, INPUT(268) => 
                           A_neg_shifted_by1_6_51_port, INPUT(269) => 
                           A_neg_shifted_by1_6_50_port, INPUT(270) => 
                           A_neg_shifted_by1_6_49_port, INPUT(271) => 
                           A_neg_shifted_by1_6_48_port, INPUT(272) => 
                           A_neg_shifted_by1_6_47_port, INPUT(273) => 
                           A_neg_shifted_by1_6_46_port, INPUT(274) => 
                           A_neg_shifted_by1_6_45_port, INPUT(275) => 
                           A_neg_shifted_by1_6_44_port, INPUT(276) => 
                           A_neg_shifted_by1_6_43_port, INPUT(277) => 
                           A_neg_shifted_by1_6_42_port, INPUT(278) => 
                           A_neg_shifted_by1_6_41_port, INPUT(279) => 
                           A_neg_shifted_by1_6_40_port, INPUT(280) => 
                           A_neg_shifted_by1_6_39_port, INPUT(281) => 
                           A_neg_shifted_by1_6_38_port, INPUT(282) => 
                           A_neg_shifted_by1_6_37_port, INPUT(283) => 
                           A_neg_shifted_by1_6_36_port, INPUT(284) => 
                           A_neg_shifted_by1_6_35_port, INPUT(285) => 
                           A_neg_shifted_by1_6_34_port, INPUT(286) => 
                           A_neg_shifted_by1_6_33_port, INPUT(287) => 
                           A_neg_shifted_by1_6_32_port, INPUT(288) => 
                           A_neg_shifted_by1_6_31_port, INPUT(289) => 
                           A_neg_shifted_by1_6_30_port, INPUT(290) => 
                           A_neg_shifted_by1_6_29_port, INPUT(291) => 
                           A_neg_shifted_by1_6_28_port, INPUT(292) => 
                           A_neg_shifted_by1_6_27_port, INPUT(293) => 
                           A_neg_shifted_by1_6_26_port, INPUT(294) => 
                           A_neg_shifted_by1_6_25_port, INPUT(295) => 
                           A_neg_shifted_by1_6_24_port, INPUT(296) => 
                           A_neg_shifted_by1_6_23_port, INPUT(297) => 
                           A_neg_shifted_by1_6_22_port, INPUT(298) => 
                           A_neg_shifted_by1_6_21_port, INPUT(299) => 
                           A_neg_shifted_by1_6_20_port, INPUT(300) => 
                           A_neg_shifted_by1_6_19_port, INPUT(301) => 
                           A_neg_shifted_by1_6_18_port, INPUT(302) => 
                           A_neg_shifted_by1_6_17_port, INPUT(303) => 
                           A_neg_shifted_by1_6_16_port, INPUT(304) => 
                           A_neg_shifted_by1_6_15_port, INPUT(305) => 
                           A_neg_shifted_by1_6_14_port, INPUT(306) => 
                           A_neg_shifted_by1_6_13_port, INPUT(307) => 
                           A_neg_shifted_by1_6_12_port, INPUT(308) => 
                           A_neg_shifted_by1_6_11_port, INPUT(309) => 
                           A_neg_shifted_by1_6_10_port, INPUT(310) => 
                           A_neg_shifted_by1_6_9_port, INPUT(311) => 
                           A_neg_shifted_by1_6_8_port, INPUT(312) => 
                           A_neg_shifted_by1_6_7_port, INPUT(313) => 
                           A_neg_shifted_by1_6_6_port, INPUT(314) => 
                           A_neg_shifted_by1_6_5_port, INPUT(315) => 
                           A_neg_shifted_by1_6_4_port, INPUT(316) => 
                           A_neg_shifted_by1_6_3_port, INPUT(317) => 
                           A_neg_shifted_by1_6_2_port, INPUT(318) => 
                           A_neg_shifted_by1_6_1_port, INPUT(319) => 
                           A_neg_shifted_by1_6_0_port, SEL(0) => 
                           selection_signal_6_2_port, SEL(1) => 
                           selection_signal_6_1_port, SEL(2) => 
                           selection_signal_6_0_port, Y(0) => OUT_MUX_6_63_port
                           , Y(1) => OUT_MUX_6_62_port, Y(2) => 
                           OUT_MUX_6_61_port, Y(3) => OUT_MUX_6_60_port, Y(4) 
                           => OUT_MUX_6_59_port, Y(5) => OUT_MUX_6_58_port, 
                           Y(6) => OUT_MUX_6_57_port, Y(7) => OUT_MUX_6_56_port
                           , Y(8) => OUT_MUX_6_55_port, Y(9) => 
                           OUT_MUX_6_54_port, Y(10) => OUT_MUX_6_53_port, Y(11)
                           => OUT_MUX_6_52_port, Y(12) => OUT_MUX_6_51_port, 
                           Y(13) => OUT_MUX_6_50_port, Y(14) => 
                           OUT_MUX_6_49_port, Y(15) => OUT_MUX_6_48_port, Y(16)
                           => OUT_MUX_6_47_port, Y(17) => OUT_MUX_6_46_port, 
                           Y(18) => OUT_MUX_6_45_port, Y(19) => 
                           OUT_MUX_6_44_port, Y(20) => OUT_MUX_6_43_port, Y(21)
                           => OUT_MUX_6_42_port, Y(22) => OUT_MUX_6_41_port, 
                           Y(23) => OUT_MUX_6_40_port, Y(24) => 
                           OUT_MUX_6_39_port, Y(25) => OUT_MUX_6_38_port, Y(26)
                           => OUT_MUX_6_37_port, Y(27) => OUT_MUX_6_36_port, 
                           Y(28) => OUT_MUX_6_35_port, Y(29) => 
                           OUT_MUX_6_34_port, Y(30) => OUT_MUX_6_33_port, Y(31)
                           => OUT_MUX_6_32_port, Y(32) => OUT_MUX_6_31_port, 
                           Y(33) => OUT_MUX_6_30_port, Y(34) => 
                           OUT_MUX_6_29_port, Y(35) => OUT_MUX_6_28_port, Y(36)
                           => OUT_MUX_6_27_port, Y(37) => OUT_MUX_6_26_port, 
                           Y(38) => OUT_MUX_6_25_port, Y(39) => 
                           OUT_MUX_6_24_port, Y(40) => OUT_MUX_6_23_port, Y(41)
                           => OUT_MUX_6_22_port, Y(42) => OUT_MUX_6_21_port, 
                           Y(43) => OUT_MUX_6_20_port, Y(44) => 
                           OUT_MUX_6_19_port, Y(45) => OUT_MUX_6_18_port, Y(46)
                           => OUT_MUX_6_17_port, Y(47) => OUT_MUX_6_16_port, 
                           Y(48) => OUT_MUX_6_15_port, Y(49) => 
                           OUT_MUX_6_14_port, Y(50) => OUT_MUX_6_13_port, Y(51)
                           => OUT_MUX_6_12_port, Y(52) => OUT_MUX_6_11_port, 
                           Y(53) => OUT_MUX_6_10_port, Y(54) => 
                           OUT_MUX_6_9_port, Y(55) => OUT_MUX_6_8_port, Y(56) 
                           => OUT_MUX_6_7_port, Y(57) => OUT_MUX_6_6_port, 
                           Y(58) => OUT_MUX_6_5_port, Y(59) => OUT_MUX_6_4_port
                           , Y(60) => OUT_MUX_6_3_port, Y(61) => 
                           OUT_MUX_6_2_port, Y(62) => OUT_MUX_6_1_port, Y(63) 
                           => OUT_MUX_6_0_port);
   MUXi_7 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_9 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_6_63_port, INPUT(65) => 
                           A_pos_shifted_by2_6_62_port, INPUT(66) => 
                           A_pos_shifted_by2_6_61_port, INPUT(67) => 
                           A_pos_shifted_by2_6_60_port, INPUT(68) => 
                           A_pos_shifted_by2_6_59_port, INPUT(69) => 
                           A_pos_shifted_by2_6_58_port, INPUT(70) => 
                           A_pos_shifted_by2_6_57_port, INPUT(71) => 
                           A_pos_shifted_by2_6_56_port, INPUT(72) => 
                           A_pos_shifted_by2_6_55_port, INPUT(73) => 
                           A_pos_shifted_by2_6_54_port, INPUT(74) => 
                           A_pos_shifted_by2_6_53_port, INPUT(75) => 
                           A_pos_shifted_by2_6_52_port, INPUT(76) => 
                           A_pos_shifted_by2_6_51_port, INPUT(77) => 
                           A_pos_shifted_by2_6_50_port, INPUT(78) => 
                           A_pos_shifted_by2_6_49_port, INPUT(79) => 
                           A_pos_shifted_by2_6_48_port, INPUT(80) => n236, 
                           INPUT(81) => A_pos_shifted_by2_6_46_port, INPUT(82) 
                           => A_pos_shifted_by2_6_45_port, INPUT(83) => 
                           A_pos_shifted_by2_6_44_port, INPUT(84) => 
                           A_pos_shifted_by2_6_43_port, INPUT(85) => 
                           A_pos_shifted_by2_6_42_port, INPUT(86) => 
                           A_pos_shifted_by2_6_41_port, INPUT(87) => 
                           A_pos_shifted_by2_6_40_port, INPUT(88) => 
                           A_pos_shifted_by2_6_39_port, INPUT(89) => 
                           A_pos_shifted_by2_6_38_port, INPUT(90) => 
                           A_pos_shifted_by2_6_37_port, INPUT(91) => 
                           A_pos_shifted_by2_6_36_port, INPUT(92) => 
                           A_pos_shifted_by2_6_35_port, INPUT(93) => 
                           A_pos_shifted_by2_6_34_port, INPUT(94) => 
                           A_pos_shifted_by2_6_33_port, INPUT(95) => 
                           A_pos_shifted_by2_6_32_port, INPUT(96) => 
                           A_pos_shifted_by2_6_31_port, INPUT(97) => 
                           A_pos_shifted_by2_6_30_port, INPUT(98) => 
                           A_pos_shifted_by2_6_29_port, INPUT(99) => 
                           A_pos_shifted_by2_6_28_port, INPUT(100) => 
                           A_pos_shifted_by2_6_27_port, INPUT(101) => 
                           A_pos_shifted_by2_6_26_port, INPUT(102) => 
                           A_pos_shifted_by2_6_25_port, INPUT(103) => 
                           A_pos_shifted_by2_6_24_port, INPUT(104) => 
                           A_pos_shifted_by2_6_23_port, INPUT(105) => 
                           A_pos_shifted_by2_6_22_port, INPUT(106) => 
                           A_pos_shifted_by2_6_21_port, INPUT(107) => 
                           A_pos_shifted_by2_6_20_port, INPUT(108) => 
                           A_pos_shifted_by2_6_19_port, INPUT(109) => 
                           A_pos_shifted_by2_6_18_port, INPUT(110) => 
                           A_pos_shifted_by2_6_17_port, INPUT(111) => 
                           A_pos_shifted_by2_6_16_port, INPUT(112) => 
                           A_pos_shifted_by2_6_15_port, INPUT(113) => 
                           A_pos_shifted_by2_6_14_port, INPUT(114) => 
                           A_pos_shifted_by2_6_13_port, INPUT(115) => 
                           A_pos_shifted_by2_6_12_port, INPUT(116) => 
                           A_pos_shifted_by2_6_11_port, INPUT(117) => 
                           A_pos_shifted_by2_6_10_port, INPUT(118) => 
                           A_pos_shifted_by2_6_9_port, INPUT(119) => 
                           A_pos_shifted_by2_6_8_port, INPUT(120) => 
                           A_pos_shifted_by2_6_7_port, INPUT(121) => 
                           A_pos_shifted_by2_6_6_port, INPUT(122) => 
                           A_pos_shifted_by2_6_5_port, INPUT(123) => 
                           A_pos_shifted_by2_6_4_port, INPUT(124) => 
                           A_pos_shifted_by2_6_3_port, INPUT(125) => 
                           A_pos_shifted_by2_6_2_port, INPUT(126) => 
                           A_pos_shifted_by2_6_1_port, INPUT(127) => 
                           A_pos_shifted_by2_6_0_port, INPUT(128) => 
                           A_neg_shifted_by2_6_63_port, INPUT(129) => 
                           A_neg_shifted_by2_6_62_port, INPUT(130) => 
                           A_neg_shifted_by2_6_61_port, INPUT(131) => 
                           A_neg_shifted_by2_6_60_port, INPUT(132) => 
                           A_neg_shifted_by2_6_59_port, INPUT(133) => 
                           A_neg_shifted_by2_6_58_port, INPUT(134) => 
                           A_neg_shifted_by2_6_57_port, INPUT(135) => 
                           A_neg_shifted_by2_6_56_port, INPUT(136) => 
                           A_neg_shifted_by2_6_55_port, INPUT(137) => 
                           A_neg_shifted_by2_6_54_port, INPUT(138) => 
                           A_neg_shifted_by2_6_53_port, INPUT(139) => 
                           A_neg_shifted_by2_6_52_port, INPUT(140) => 
                           A_neg_shifted_by2_6_51_port, INPUT(141) => 
                           A_neg_shifted_by2_6_50_port, INPUT(142) => 
                           A_neg_shifted_by2_6_49_port, INPUT(143) => 
                           A_neg_shifted_by2_6_48_port, INPUT(144) => n202, 
                           INPUT(145) => A_neg_shifted_by2_6_46_port, 
                           INPUT(146) => A_neg_shifted_by2_6_45_port, 
                           INPUT(147) => A_neg_shifted_by2_6_44_port, 
                           INPUT(148) => A_neg_shifted_by2_6_43_port, 
                           INPUT(149) => A_neg_shifted_by2_6_42_port, 
                           INPUT(150) => A_neg_shifted_by2_6_41_port, 
                           INPUT(151) => A_neg_shifted_by2_6_40_port, 
                           INPUT(152) => A_neg_shifted_by2_6_39_port, 
                           INPUT(153) => A_neg_shifted_by2_6_38_port, 
                           INPUT(154) => A_neg_shifted_by2_6_37_port, 
                           INPUT(155) => A_neg_shifted_by2_6_36_port, 
                           INPUT(156) => A_neg_shifted_by2_6_35_port, 
                           INPUT(157) => A_neg_shifted_by2_6_34_port, 
                           INPUT(158) => A_neg_shifted_by2_6_33_port, 
                           INPUT(159) => A_neg_shifted_by2_6_32_port, 
                           INPUT(160) => A_neg_shifted_by2_6_31_port, 
                           INPUT(161) => A_neg_shifted_by2_6_30_port, 
                           INPUT(162) => A_neg_shifted_by2_6_29_port, 
                           INPUT(163) => A_neg_shifted_by2_6_28_port, 
                           INPUT(164) => A_neg_shifted_by2_6_27_port, 
                           INPUT(165) => A_neg_shifted_by2_6_26_port, 
                           INPUT(166) => A_neg_shifted_by2_6_25_port, 
                           INPUT(167) => A_neg_shifted_by2_6_24_port, 
                           INPUT(168) => A_neg_shifted_by2_6_23_port, 
                           INPUT(169) => A_neg_shifted_by2_6_22_port, 
                           INPUT(170) => A_neg_shifted_by2_6_21_port, 
                           INPUT(171) => A_neg_shifted_by2_6_20_port, 
                           INPUT(172) => A_neg_shifted_by2_6_19_port, 
                           INPUT(173) => A_neg_shifted_by2_6_18_port, 
                           INPUT(174) => A_neg_shifted_by2_6_17_port, 
                           INPUT(175) => A_neg_shifted_by2_6_16_port, 
                           INPUT(176) => A_neg_shifted_by2_6_15_port, 
                           INPUT(177) => A_neg_shifted_by2_6_14_port, 
                           INPUT(178) => A_neg_shifted_by2_6_13_port, 
                           INPUT(179) => A_neg_shifted_by2_6_12_port, 
                           INPUT(180) => A_neg_shifted_by2_6_11_port, 
                           INPUT(181) => A_neg_shifted_by2_6_10_port, 
                           INPUT(182) => A_neg_shifted_by2_6_9_port, INPUT(183)
                           => A_neg_shifted_by2_6_8_port, INPUT(184) => 
                           A_neg_shifted_by2_6_7_port, INPUT(185) => 
                           A_neg_shifted_by2_6_6_port, INPUT(186) => 
                           A_neg_shifted_by2_6_5_port, INPUT(187) => 
                           A_neg_shifted_by2_6_4_port, INPUT(188) => 
                           A_neg_shifted_by2_6_3_port, INPUT(189) => 
                           A_neg_shifted_by2_6_2_port, INPUT(190) => 
                           A_neg_shifted_by2_6_1_port, INPUT(191) => 
                           A_neg_shifted_by2_6_0_port, INPUT(192) => 
                           A_pos_shifted_by1_7_63_port, INPUT(193) => 
                           A_pos_shifted_by1_7_62_port, INPUT(194) => 
                           A_pos_shifted_by1_7_61_port, INPUT(195) => 
                           A_pos_shifted_by1_7_60_port, INPUT(196) => 
                           A_pos_shifted_by1_7_59_port, INPUT(197) => 
                           A_pos_shifted_by1_7_58_port, INPUT(198) => 
                           A_pos_shifted_by1_7_57_port, INPUT(199) => 
                           A_pos_shifted_by1_7_56_port, INPUT(200) => 
                           A_pos_shifted_by1_7_55_port, INPUT(201) => 
                           A_pos_shifted_by1_7_54_port, INPUT(202) => 
                           A_pos_shifted_by1_7_53_port, INPUT(203) => 
                           A_pos_shifted_by1_7_52_port, INPUT(204) => 
                           A_pos_shifted_by1_7_51_port, INPUT(205) => 
                           A_pos_shifted_by1_7_50_port, INPUT(206) => 
                           A_pos_shifted_by1_7_49_port, INPUT(207) => 
                           A_pos_shifted_by1_7_48_port, INPUT(208) => 
                           A_pos_shifted_by1_7_47_port, INPUT(209) => 
                           A_pos_shifted_by1_7_46_port, INPUT(210) => 
                           A_pos_shifted_by1_7_45_port, INPUT(211) => 
                           A_pos_shifted_by1_7_44_port, INPUT(212) => 
                           A_pos_shifted_by1_7_43_port, INPUT(213) => 
                           A_pos_shifted_by1_7_42_port, INPUT(214) => 
                           A_pos_shifted_by1_7_41_port, INPUT(215) => 
                           A_pos_shifted_by1_7_40_port, INPUT(216) => 
                           A_pos_shifted_by1_7_39_port, INPUT(217) => 
                           A_pos_shifted_by1_7_38_port, INPUT(218) => 
                           A_pos_shifted_by1_7_37_port, INPUT(219) => 
                           A_pos_shifted_by1_7_36_port, INPUT(220) => 
                           A_pos_shifted_by1_7_35_port, INPUT(221) => 
                           A_pos_shifted_by1_7_34_port, INPUT(222) => 
                           A_pos_shifted_by1_7_33_port, INPUT(223) => 
                           A_pos_shifted_by1_7_32_port, INPUT(224) => 
                           A_pos_shifted_by1_7_31_port, INPUT(225) => 
                           A_pos_shifted_by1_7_30_port, INPUT(226) => 
                           A_pos_shifted_by1_7_29_port, INPUT(227) => 
                           A_pos_shifted_by1_7_28_port, INPUT(228) => 
                           A_pos_shifted_by1_7_27_port, INPUT(229) => 
                           A_pos_shifted_by1_7_26_port, INPUT(230) => 
                           A_pos_shifted_by1_7_25_port, INPUT(231) => 
                           A_pos_shifted_by1_7_24_port, INPUT(232) => 
                           A_pos_shifted_by1_7_23_port, INPUT(233) => 
                           A_pos_shifted_by1_7_22_port, INPUT(234) => 
                           A_pos_shifted_by1_7_21_port, INPUT(235) => 
                           A_pos_shifted_by1_7_20_port, INPUT(236) => 
                           A_pos_shifted_by1_7_19_port, INPUT(237) => 
                           A_pos_shifted_by1_7_18_port, INPUT(238) => 
                           A_pos_shifted_by1_7_17_port, INPUT(239) => 
                           A_pos_shifted_by1_7_16_port, INPUT(240) => 
                           A_pos_shifted_by1_7_15_port, INPUT(241) => 
                           A_pos_shifted_by1_7_14_port, INPUT(242) => 
                           A_pos_shifted_by1_7_13_port, INPUT(243) => 
                           A_pos_shifted_by1_7_12_port, INPUT(244) => 
                           A_pos_shifted_by1_7_11_port, INPUT(245) => 
                           A_pos_shifted_by1_7_10_port, INPUT(246) => 
                           A_pos_shifted_by1_7_9_port, INPUT(247) => 
                           A_pos_shifted_by1_7_8_port, INPUT(248) => 
                           A_pos_shifted_by1_7_7_port, INPUT(249) => 
                           A_pos_shifted_by1_7_6_port, INPUT(250) => 
                           A_pos_shifted_by1_7_5_port, INPUT(251) => 
                           A_pos_shifted_by1_7_4_port, INPUT(252) => 
                           A_pos_shifted_by1_7_3_port, INPUT(253) => 
                           A_pos_shifted_by1_7_2_port, INPUT(254) => 
                           A_pos_shifted_by1_7_1_port, INPUT(255) => 
                           A_pos_shifted_by1_7_0_port, INPUT(256) => 
                           A_neg_shifted_by1_7_63_port, INPUT(257) => 
                           A_neg_shifted_by1_7_62_port, INPUT(258) => 
                           A_neg_shifted_by1_7_61_port, INPUT(259) => 
                           A_neg_shifted_by1_7_60_port, INPUT(260) => 
                           A_neg_shifted_by1_7_59_port, INPUT(261) => 
                           A_neg_shifted_by1_7_58_port, INPUT(262) => 
                           A_neg_shifted_by1_7_57_port, INPUT(263) => 
                           A_neg_shifted_by1_7_56_port, INPUT(264) => 
                           A_neg_shifted_by1_7_55_port, INPUT(265) => 
                           A_neg_shifted_by1_7_54_port, INPUT(266) => 
                           A_neg_shifted_by1_7_53_port, INPUT(267) => 
                           A_neg_shifted_by1_7_52_port, INPUT(268) => 
                           A_neg_shifted_by1_7_51_port, INPUT(269) => 
                           A_neg_shifted_by1_7_50_port, INPUT(270) => 
                           A_neg_shifted_by1_7_49_port, INPUT(271) => 
                           A_neg_shifted_by1_7_48_port, INPUT(272) => 
                           A_neg_shifted_by1_7_47_port, INPUT(273) => 
                           A_neg_shifted_by1_7_46_port, INPUT(274) => 
                           A_neg_shifted_by1_7_45_port, INPUT(275) => 
                           A_neg_shifted_by1_7_44_port, INPUT(276) => 
                           A_neg_shifted_by1_7_43_port, INPUT(277) => 
                           A_neg_shifted_by1_7_42_port, INPUT(278) => 
                           A_neg_shifted_by1_7_41_port, INPUT(279) => 
                           A_neg_shifted_by1_7_40_port, INPUT(280) => 
                           A_neg_shifted_by1_7_39_port, INPUT(281) => 
                           A_neg_shifted_by1_7_38_port, INPUT(282) => 
                           A_neg_shifted_by1_7_37_port, INPUT(283) => 
                           A_neg_shifted_by1_7_36_port, INPUT(284) => 
                           A_neg_shifted_by1_7_35_port, INPUT(285) => 
                           A_neg_shifted_by1_7_34_port, INPUT(286) => 
                           A_neg_shifted_by1_7_33_port, INPUT(287) => 
                           A_neg_shifted_by1_7_32_port, INPUT(288) => 
                           A_neg_shifted_by1_7_31_port, INPUT(289) => 
                           A_neg_shifted_by1_7_30_port, INPUT(290) => 
                           A_neg_shifted_by1_7_29_port, INPUT(291) => 
                           A_neg_shifted_by1_7_28_port, INPUT(292) => 
                           A_neg_shifted_by1_7_27_port, INPUT(293) => 
                           A_neg_shifted_by1_7_26_port, INPUT(294) => 
                           A_neg_shifted_by1_7_25_port, INPUT(295) => 
                           A_neg_shifted_by1_7_24_port, INPUT(296) => 
                           A_neg_shifted_by1_7_23_port, INPUT(297) => 
                           A_neg_shifted_by1_7_22_port, INPUT(298) => 
                           A_neg_shifted_by1_7_21_port, INPUT(299) => 
                           A_neg_shifted_by1_7_20_port, INPUT(300) => 
                           A_neg_shifted_by1_7_19_port, INPUT(301) => 
                           A_neg_shifted_by1_7_18_port, INPUT(302) => 
                           A_neg_shifted_by1_7_17_port, INPUT(303) => 
                           A_neg_shifted_by1_7_16_port, INPUT(304) => 
                           A_neg_shifted_by1_7_15_port, INPUT(305) => 
                           A_neg_shifted_by1_7_14_port, INPUT(306) => 
                           A_neg_shifted_by1_7_13_port, INPUT(307) => 
                           A_neg_shifted_by1_7_12_port, INPUT(308) => 
                           A_neg_shifted_by1_7_11_port, INPUT(309) => 
                           A_neg_shifted_by1_7_10_port, INPUT(310) => 
                           A_neg_shifted_by1_7_9_port, INPUT(311) => 
                           A_neg_shifted_by1_7_8_port, INPUT(312) => 
                           A_neg_shifted_by1_7_7_port, INPUT(313) => 
                           A_neg_shifted_by1_7_6_port, INPUT(314) => 
                           A_neg_shifted_by1_7_5_port, INPUT(315) => 
                           A_neg_shifted_by1_7_4_port, INPUT(316) => 
                           A_neg_shifted_by1_7_3_port, INPUT(317) => 
                           A_neg_shifted_by1_7_2_port, INPUT(318) => 
                           A_neg_shifted_by1_7_1_port, INPUT(319) => 
                           A_neg_shifted_by1_7_0_port, SEL(0) => 
                           selection_signal_7_2_port, SEL(1) => 
                           selection_signal_7_1_port, SEL(2) => 
                           selection_signal_7_0_port, Y(0) => OUT_MUX_7_63_port
                           , Y(1) => OUT_MUX_7_62_port, Y(2) => 
                           OUT_MUX_7_61_port, Y(3) => OUT_MUX_7_60_port, Y(4) 
                           => OUT_MUX_7_59_port, Y(5) => OUT_MUX_7_58_port, 
                           Y(6) => OUT_MUX_7_57_port, Y(7) => OUT_MUX_7_56_port
                           , Y(8) => OUT_MUX_7_55_port, Y(9) => 
                           OUT_MUX_7_54_port, Y(10) => OUT_MUX_7_53_port, Y(11)
                           => OUT_MUX_7_52_port, Y(12) => OUT_MUX_7_51_port, 
                           Y(13) => OUT_MUX_7_50_port, Y(14) => 
                           OUT_MUX_7_49_port, Y(15) => OUT_MUX_7_48_port, Y(16)
                           => OUT_MUX_7_47_port, Y(17) => OUT_MUX_7_46_port, 
                           Y(18) => OUT_MUX_7_45_port, Y(19) => 
                           OUT_MUX_7_44_port, Y(20) => OUT_MUX_7_43_port, Y(21)
                           => OUT_MUX_7_42_port, Y(22) => OUT_MUX_7_41_port, 
                           Y(23) => OUT_MUX_7_40_port, Y(24) => 
                           OUT_MUX_7_39_port, Y(25) => OUT_MUX_7_38_port, Y(26)
                           => OUT_MUX_7_37_port, Y(27) => OUT_MUX_7_36_port, 
                           Y(28) => OUT_MUX_7_35_port, Y(29) => 
                           OUT_MUX_7_34_port, Y(30) => OUT_MUX_7_33_port, Y(31)
                           => OUT_MUX_7_32_port, Y(32) => OUT_MUX_7_31_port, 
                           Y(33) => OUT_MUX_7_30_port, Y(34) => 
                           OUT_MUX_7_29_port, Y(35) => OUT_MUX_7_28_port, Y(36)
                           => OUT_MUX_7_27_port, Y(37) => OUT_MUX_7_26_port, 
                           Y(38) => OUT_MUX_7_25_port, Y(39) => 
                           OUT_MUX_7_24_port, Y(40) => OUT_MUX_7_23_port, Y(41)
                           => OUT_MUX_7_22_port, Y(42) => OUT_MUX_7_21_port, 
                           Y(43) => OUT_MUX_7_20_port, Y(44) => 
                           OUT_MUX_7_19_port, Y(45) => OUT_MUX_7_18_port, Y(46)
                           => OUT_MUX_7_17_port, Y(47) => OUT_MUX_7_16_port, 
                           Y(48) => OUT_MUX_7_15_port, Y(49) => 
                           OUT_MUX_7_14_port, Y(50) => OUT_MUX_7_13_port, Y(51)
                           => OUT_MUX_7_12_port, Y(52) => OUT_MUX_7_11_port, 
                           Y(53) => OUT_MUX_7_10_port, Y(54) => 
                           OUT_MUX_7_9_port, Y(55) => OUT_MUX_7_8_port, Y(56) 
                           => OUT_MUX_7_7_port, Y(57) => OUT_MUX_7_6_port, 
                           Y(58) => OUT_MUX_7_5_port, Y(59) => OUT_MUX_7_4_port
                           , Y(60) => OUT_MUX_7_3_port, Y(61) => 
                           OUT_MUX_7_2_port, Y(62) => OUT_MUX_7_1_port, Y(63) 
                           => OUT_MUX_7_0_port);
   MUXi_8 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_8 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_7_63_port, INPUT(65) => 
                           A_pos_shifted_by2_7_62_port, INPUT(66) => 
                           A_pos_shifted_by2_7_61_port, INPUT(67) => 
                           A_pos_shifted_by2_7_60_port, INPUT(68) => 
                           A_pos_shifted_by2_7_59_port, INPUT(69) => 
                           A_pos_shifted_by2_7_58_port, INPUT(70) => 
                           A_pos_shifted_by2_7_57_port, INPUT(71) => 
                           A_pos_shifted_by2_7_56_port, INPUT(72) => 
                           A_pos_shifted_by2_7_55_port, INPUT(73) => 
                           A_pos_shifted_by2_7_54_port, INPUT(74) => 
                           A_pos_shifted_by2_7_53_port, INPUT(75) => 
                           A_pos_shifted_by2_7_52_port, INPUT(76) => 
                           A_pos_shifted_by2_7_51_port, INPUT(77) => 
                           A_pos_shifted_by2_7_50_port, INPUT(78) => 
                           A_pos_shifted_by2_7_49_port, INPUT(79) => 
                           A_pos_shifted_by2_7_48_port, INPUT(80) => 
                           A_pos_shifted_by2_7_47_port, INPUT(81) => 
                           A_pos_shifted_by2_7_46_port, INPUT(82) => 
                           A_pos_shifted_by2_7_45_port, INPUT(83) => 
                           A_pos_shifted_by2_7_44_port, INPUT(84) => 
                           A_pos_shifted_by2_7_43_port, INPUT(85) => 
                           A_pos_shifted_by2_7_42_port, INPUT(86) => 
                           A_pos_shifted_by2_7_41_port, INPUT(87) => 
                           A_pos_shifted_by2_7_40_port, INPUT(88) => 
                           A_pos_shifted_by2_7_39_port, INPUT(89) => 
                           A_pos_shifted_by2_7_38_port, INPUT(90) => 
                           A_pos_shifted_by2_7_37_port, INPUT(91) => 
                           A_pos_shifted_by2_7_36_port, INPUT(92) => 
                           A_pos_shifted_by2_7_35_port, INPUT(93) => 
                           A_pos_shifted_by2_7_34_port, INPUT(94) => 
                           A_pos_shifted_by2_7_33_port, INPUT(95) => 
                           A_pos_shifted_by2_7_32_port, INPUT(96) => 
                           A_pos_shifted_by2_7_31_port, INPUT(97) => 
                           A_pos_shifted_by2_7_30_port, INPUT(98) => 
                           A_pos_shifted_by2_7_29_port, INPUT(99) => 
                           A_pos_shifted_by2_7_28_port, INPUT(100) => 
                           A_pos_shifted_by2_7_27_port, INPUT(101) => 
                           A_pos_shifted_by2_7_26_port, INPUT(102) => 
                           A_pos_shifted_by2_7_25_port, INPUT(103) => 
                           A_pos_shifted_by2_7_24_port, INPUT(104) => 
                           A_pos_shifted_by2_7_23_port, INPUT(105) => 
                           A_pos_shifted_by2_7_22_port, INPUT(106) => 
                           A_pos_shifted_by2_7_21_port, INPUT(107) => 
                           A_pos_shifted_by2_7_20_port, INPUT(108) => 
                           A_pos_shifted_by2_7_19_port, INPUT(109) => 
                           A_pos_shifted_by2_7_18_port, INPUT(110) => 
                           A_pos_shifted_by2_7_17_port, INPUT(111) => 
                           A_pos_shifted_by2_7_16_port, INPUT(112) => 
                           A_pos_shifted_by2_7_15_port, INPUT(113) => 
                           A_pos_shifted_by2_7_14_port, INPUT(114) => 
                           A_pos_shifted_by2_7_13_port, INPUT(115) => 
                           A_pos_shifted_by2_7_12_port, INPUT(116) => 
                           A_pos_shifted_by2_7_11_port, INPUT(117) => 
                           A_pos_shifted_by2_7_10_port, INPUT(118) => 
                           A_pos_shifted_by2_7_9_port, INPUT(119) => 
                           A_pos_shifted_by2_7_8_port, INPUT(120) => 
                           A_pos_shifted_by2_7_7_port, INPUT(121) => 
                           A_pos_shifted_by2_7_6_port, INPUT(122) => 
                           A_pos_shifted_by2_7_5_port, INPUT(123) => 
                           A_pos_shifted_by2_7_4_port, INPUT(124) => 
                           A_pos_shifted_by2_7_3_port, INPUT(125) => 
                           A_pos_shifted_by2_7_2_port, INPUT(126) => 
                           A_pos_shifted_by2_7_1_port, INPUT(127) => 
                           A_pos_shifted_by2_7_0_port, INPUT(128) => 
                           A_neg_shifted_by2_7_63_port, INPUT(129) => 
                           A_neg_shifted_by2_7_62_port, INPUT(130) => 
                           A_neg_shifted_by2_7_61_port, INPUT(131) => 
                           A_neg_shifted_by2_7_60_port, INPUT(132) => 
                           A_neg_shifted_by2_7_59_port, INPUT(133) => 
                           A_neg_shifted_by2_7_58_port, INPUT(134) => 
                           A_neg_shifted_by2_7_57_port, INPUT(135) => 
                           A_neg_shifted_by2_7_56_port, INPUT(136) => 
                           A_neg_shifted_by2_7_55_port, INPUT(137) => 
                           A_neg_shifted_by2_7_54_port, INPUT(138) => 
                           A_neg_shifted_by2_7_53_port, INPUT(139) => 
                           A_neg_shifted_by2_7_52_port, INPUT(140) => 
                           A_neg_shifted_by2_7_51_port, INPUT(141) => 
                           A_neg_shifted_by2_7_50_port, INPUT(142) => 
                           A_neg_shifted_by2_7_49_port, INPUT(143) => 
                           A_neg_shifted_by2_7_48_port, INPUT(144) => 
                           A_neg_shifted_by2_7_47_port, INPUT(145) => 
                           A_neg_shifted_by2_7_46_port, INPUT(146) => 
                           A_neg_shifted_by2_7_45_port, INPUT(147) => 
                           A_neg_shifted_by2_7_44_port, INPUT(148) => 
                           A_neg_shifted_by2_7_43_port, INPUT(149) => 
                           A_neg_shifted_by2_7_42_port, INPUT(150) => 
                           A_neg_shifted_by2_7_41_port, INPUT(151) => 
                           A_neg_shifted_by2_7_40_port, INPUT(152) => 
                           A_neg_shifted_by2_7_39_port, INPUT(153) => 
                           A_neg_shifted_by2_7_38_port, INPUT(154) => 
                           A_neg_shifted_by2_7_37_port, INPUT(155) => 
                           A_neg_shifted_by2_7_36_port, INPUT(156) => 
                           A_neg_shifted_by2_7_35_port, INPUT(157) => 
                           A_neg_shifted_by2_7_34_port, INPUT(158) => 
                           A_neg_shifted_by2_7_33_port, INPUT(159) => 
                           A_neg_shifted_by2_7_32_port, INPUT(160) => 
                           A_neg_shifted_by2_7_31_port, INPUT(161) => 
                           A_neg_shifted_by2_7_30_port, INPUT(162) => 
                           A_neg_shifted_by2_7_29_port, INPUT(163) => 
                           A_neg_shifted_by2_7_28_port, INPUT(164) => 
                           A_neg_shifted_by2_7_27_port, INPUT(165) => 
                           A_neg_shifted_by2_7_26_port, INPUT(166) => 
                           A_neg_shifted_by2_7_25_port, INPUT(167) => 
                           A_neg_shifted_by2_7_24_port, INPUT(168) => 
                           A_neg_shifted_by2_7_23_port, INPUT(169) => 
                           A_neg_shifted_by2_7_22_port, INPUT(170) => 
                           A_neg_shifted_by2_7_21_port, INPUT(171) => 
                           A_neg_shifted_by2_7_20_port, INPUT(172) => 
                           A_neg_shifted_by2_7_19_port, INPUT(173) => 
                           A_neg_shifted_by2_7_18_port, INPUT(174) => 
                           A_neg_shifted_by2_7_17_port, INPUT(175) => 
                           A_neg_shifted_by2_7_16_port, INPUT(176) => 
                           A_neg_shifted_by2_7_15_port, INPUT(177) => 
                           A_neg_shifted_by2_7_14_port, INPUT(178) => 
                           A_neg_shifted_by2_7_13_port, INPUT(179) => 
                           A_neg_shifted_by2_7_12_port, INPUT(180) => 
                           A_neg_shifted_by2_7_11_port, INPUT(181) => 
                           A_neg_shifted_by2_7_10_port, INPUT(182) => 
                           A_neg_shifted_by2_7_9_port, INPUT(183) => 
                           A_neg_shifted_by2_7_8_port, INPUT(184) => 
                           A_neg_shifted_by2_7_7_port, INPUT(185) => 
                           A_neg_shifted_by2_7_6_port, INPUT(186) => 
                           A_neg_shifted_by2_7_5_port, INPUT(187) => 
                           A_neg_shifted_by2_7_4_port, INPUT(188) => 
                           A_neg_shifted_by2_7_3_port, INPUT(189) => 
                           A_neg_shifted_by2_7_2_port, INPUT(190) => 
                           A_neg_shifted_by2_7_1_port, INPUT(191) => 
                           A_neg_shifted_by2_7_0_port, INPUT(192) => 
                           A_pos_shifted_by1_8_63_port, INPUT(193) => 
                           A_pos_shifted_by1_8_62_port, INPUT(194) => 
                           A_pos_shifted_by1_8_61_port, INPUT(195) => 
                           A_pos_shifted_by1_8_60_port, INPUT(196) => 
                           A_pos_shifted_by1_8_59_port, INPUT(197) => 
                           A_pos_shifted_by1_8_58_port, INPUT(198) => 
                           A_pos_shifted_by1_8_57_port, INPUT(199) => 
                           A_pos_shifted_by1_8_56_port, INPUT(200) => 
                           A_pos_shifted_by1_8_55_port, INPUT(201) => 
                           A_pos_shifted_by1_8_54_port, INPUT(202) => 
                           A_pos_shifted_by1_8_53_port, INPUT(203) => 
                           A_pos_shifted_by1_8_52_port, INPUT(204) => 
                           A_pos_shifted_by1_8_51_port, INPUT(205) => 
                           A_pos_shifted_by1_8_50_port, INPUT(206) => 
                           A_pos_shifted_by1_8_49_port, INPUT(207) => 
                           A_pos_shifted_by1_8_48_port, INPUT(208) => 
                           A_pos_shifted_by1_8_47_port, INPUT(209) => 
                           A_pos_shifted_by1_8_46_port, INPUT(210) => 
                           A_pos_shifted_by1_8_45_port, INPUT(211) => 
                           A_pos_shifted_by1_8_44_port, INPUT(212) => 
                           A_pos_shifted_by1_8_43_port, INPUT(213) => 
                           A_pos_shifted_by1_8_42_port, INPUT(214) => 
                           A_pos_shifted_by1_8_41_port, INPUT(215) => 
                           A_pos_shifted_by1_8_40_port, INPUT(216) => 
                           A_pos_shifted_by1_8_39_port, INPUT(217) => 
                           A_pos_shifted_by1_8_38_port, INPUT(218) => 
                           A_pos_shifted_by1_8_37_port, INPUT(219) => 
                           A_pos_shifted_by1_8_36_port, INPUT(220) => 
                           A_pos_shifted_by1_8_35_port, INPUT(221) => 
                           A_pos_shifted_by1_8_34_port, INPUT(222) => 
                           A_pos_shifted_by1_8_33_port, INPUT(223) => 
                           A_pos_shifted_by1_8_32_port, INPUT(224) => 
                           A_pos_shifted_by1_8_31_port, INPUT(225) => 
                           A_pos_shifted_by1_8_30_port, INPUT(226) => 
                           A_pos_shifted_by1_8_29_port, INPUT(227) => 
                           A_pos_shifted_by1_8_28_port, INPUT(228) => 
                           A_pos_shifted_by1_8_27_port, INPUT(229) => 
                           A_pos_shifted_by1_8_26_port, INPUT(230) => 
                           A_pos_shifted_by1_8_25_port, INPUT(231) => 
                           A_pos_shifted_by1_8_24_port, INPUT(232) => 
                           A_pos_shifted_by1_8_23_port, INPUT(233) => 
                           A_pos_shifted_by1_8_22_port, INPUT(234) => 
                           A_pos_shifted_by1_8_21_port, INPUT(235) => 
                           A_pos_shifted_by1_8_20_port, INPUT(236) => 
                           A_pos_shifted_by1_8_19_port, INPUT(237) => 
                           A_pos_shifted_by1_8_18_port, INPUT(238) => 
                           A_pos_shifted_by1_8_17_port, INPUT(239) => 
                           A_pos_shifted_by1_8_16_port, INPUT(240) => 
                           A_pos_shifted_by1_8_15_port, INPUT(241) => 
                           A_pos_shifted_by1_8_14_port, INPUT(242) => 
                           A_pos_shifted_by1_8_13_port, INPUT(243) => 
                           A_pos_shifted_by1_8_12_port, INPUT(244) => 
                           A_pos_shifted_by1_8_11_port, INPUT(245) => 
                           A_pos_shifted_by1_8_10_port, INPUT(246) => 
                           A_pos_shifted_by1_8_9_port, INPUT(247) => 
                           A_pos_shifted_by1_8_8_port, INPUT(248) => 
                           A_pos_shifted_by1_8_7_port, INPUT(249) => 
                           A_pos_shifted_by1_8_6_port, INPUT(250) => 
                           A_pos_shifted_by1_8_5_port, INPUT(251) => 
                           A_pos_shifted_by1_8_4_port, INPUT(252) => 
                           A_pos_shifted_by1_8_3_port, INPUT(253) => 
                           A_pos_shifted_by1_8_2_port, INPUT(254) => 
                           A_pos_shifted_by1_8_1_port, INPUT(255) => 
                           A_pos_shifted_by1_8_0_port, INPUT(256) => 
                           A_neg_shifted_by1_8_63_port, INPUT(257) => 
                           A_neg_shifted_by1_8_62_port, INPUT(258) => 
                           A_neg_shifted_by1_8_61_port, INPUT(259) => 
                           A_neg_shifted_by1_8_60_port, INPUT(260) => 
                           A_neg_shifted_by1_8_59_port, INPUT(261) => 
                           A_neg_shifted_by1_8_58_port, INPUT(262) => 
                           A_neg_shifted_by1_8_57_port, INPUT(263) => 
                           A_neg_shifted_by1_8_56_port, INPUT(264) => 
                           A_neg_shifted_by1_8_55_port, INPUT(265) => 
                           A_neg_shifted_by1_8_54_port, INPUT(266) => 
                           A_neg_shifted_by1_8_53_port, INPUT(267) => 
                           A_neg_shifted_by1_8_52_port, INPUT(268) => 
                           A_neg_shifted_by1_8_51_port, INPUT(269) => 
                           A_neg_shifted_by1_8_50_port, INPUT(270) => 
                           A_neg_shifted_by1_8_49_port, INPUT(271) => 
                           A_neg_shifted_by1_8_48_port, INPUT(272) => 
                           A_neg_shifted_by1_8_47_port, INPUT(273) => 
                           A_neg_shifted_by1_8_46_port, INPUT(274) => 
                           A_neg_shifted_by1_8_45_port, INPUT(275) => 
                           A_neg_shifted_by1_8_44_port, INPUT(276) => 
                           A_neg_shifted_by1_8_43_port, INPUT(277) => 
                           A_neg_shifted_by1_8_42_port, INPUT(278) => 
                           A_neg_shifted_by1_8_41_port, INPUT(279) => 
                           A_neg_shifted_by1_8_40_port, INPUT(280) => 
                           A_neg_shifted_by1_8_39_port, INPUT(281) => 
                           A_neg_shifted_by1_8_38_port, INPUT(282) => 
                           A_neg_shifted_by1_8_37_port, INPUT(283) => 
                           A_neg_shifted_by1_8_36_port, INPUT(284) => 
                           A_neg_shifted_by1_8_35_port, INPUT(285) => 
                           A_neg_shifted_by1_8_34_port, INPUT(286) => 
                           A_neg_shifted_by1_8_33_port, INPUT(287) => 
                           A_neg_shifted_by1_8_32_port, INPUT(288) => 
                           A_neg_shifted_by1_8_31_port, INPUT(289) => 
                           A_neg_shifted_by1_8_30_port, INPUT(290) => 
                           A_neg_shifted_by1_8_29_port, INPUT(291) => 
                           A_neg_shifted_by1_8_28_port, INPUT(292) => 
                           A_neg_shifted_by1_8_27_port, INPUT(293) => 
                           A_neg_shifted_by1_8_26_port, INPUT(294) => 
                           A_neg_shifted_by1_8_25_port, INPUT(295) => 
                           A_neg_shifted_by1_8_24_port, INPUT(296) => 
                           A_neg_shifted_by1_8_23_port, INPUT(297) => 
                           A_neg_shifted_by1_8_22_port, INPUT(298) => 
                           A_neg_shifted_by1_8_21_port, INPUT(299) => 
                           A_neg_shifted_by1_8_20_port, INPUT(300) => 
                           A_neg_shifted_by1_8_19_port, INPUT(301) => 
                           A_neg_shifted_by1_8_18_port, INPUT(302) => 
                           A_neg_shifted_by1_8_17_port, INPUT(303) => 
                           A_neg_shifted_by1_8_16_port, INPUT(304) => 
                           A_neg_shifted_by1_8_15_port, INPUT(305) => 
                           A_neg_shifted_by1_8_14_port, INPUT(306) => 
                           A_neg_shifted_by1_8_13_port, INPUT(307) => 
                           A_neg_shifted_by1_8_12_port, INPUT(308) => 
                           A_neg_shifted_by1_8_11_port, INPUT(309) => 
                           A_neg_shifted_by1_8_10_port, INPUT(310) => 
                           A_neg_shifted_by1_8_9_port, INPUT(311) => 
                           A_neg_shifted_by1_8_8_port, INPUT(312) => 
                           A_neg_shifted_by1_8_7_port, INPUT(313) => 
                           A_neg_shifted_by1_8_6_port, INPUT(314) => 
                           A_neg_shifted_by1_8_5_port, INPUT(315) => 
                           A_neg_shifted_by1_8_4_port, INPUT(316) => 
                           A_neg_shifted_by1_8_3_port, INPUT(317) => 
                           A_neg_shifted_by1_8_2_port, INPUT(318) => 
                           A_neg_shifted_by1_8_1_port, INPUT(319) => 
                           A_neg_shifted_by1_8_0_port, SEL(0) => 
                           selection_signal_8_2_port, SEL(1) => 
                           selection_signal_8_1_port, SEL(2) => 
                           selection_signal_8_0_port, Y(0) => OUT_MUX_8_63_port
                           , Y(1) => OUT_MUX_8_62_port, Y(2) => 
                           OUT_MUX_8_61_port, Y(3) => OUT_MUX_8_60_port, Y(4) 
                           => OUT_MUX_8_59_port, Y(5) => OUT_MUX_8_58_port, 
                           Y(6) => OUT_MUX_8_57_port, Y(7) => OUT_MUX_8_56_port
                           , Y(8) => OUT_MUX_8_55_port, Y(9) => 
                           OUT_MUX_8_54_port, Y(10) => OUT_MUX_8_53_port, Y(11)
                           => OUT_MUX_8_52_port, Y(12) => OUT_MUX_8_51_port, 
                           Y(13) => OUT_MUX_8_50_port, Y(14) => 
                           OUT_MUX_8_49_port, Y(15) => OUT_MUX_8_48_port, Y(16)
                           => OUT_MUX_8_47_port, Y(17) => OUT_MUX_8_46_port, 
                           Y(18) => OUT_MUX_8_45_port, Y(19) => 
                           OUT_MUX_8_44_port, Y(20) => OUT_MUX_8_43_port, Y(21)
                           => OUT_MUX_8_42_port, Y(22) => OUT_MUX_8_41_port, 
                           Y(23) => OUT_MUX_8_40_port, Y(24) => 
                           OUT_MUX_8_39_port, Y(25) => OUT_MUX_8_38_port, Y(26)
                           => OUT_MUX_8_37_port, Y(27) => OUT_MUX_8_36_port, 
                           Y(28) => OUT_MUX_8_35_port, Y(29) => 
                           OUT_MUX_8_34_port, Y(30) => OUT_MUX_8_33_port, Y(31)
                           => OUT_MUX_8_32_port, Y(32) => OUT_MUX_8_31_port, 
                           Y(33) => OUT_MUX_8_30_port, Y(34) => 
                           OUT_MUX_8_29_port, Y(35) => OUT_MUX_8_28_port, Y(36)
                           => OUT_MUX_8_27_port, Y(37) => OUT_MUX_8_26_port, 
                           Y(38) => OUT_MUX_8_25_port, Y(39) => 
                           OUT_MUX_8_24_port, Y(40) => OUT_MUX_8_23_port, Y(41)
                           => OUT_MUX_8_22_port, Y(42) => OUT_MUX_8_21_port, 
                           Y(43) => OUT_MUX_8_20_port, Y(44) => 
                           OUT_MUX_8_19_port, Y(45) => OUT_MUX_8_18_port, Y(46)
                           => OUT_MUX_8_17_port, Y(47) => OUT_MUX_8_16_port, 
                           Y(48) => OUT_MUX_8_15_port, Y(49) => 
                           OUT_MUX_8_14_port, Y(50) => OUT_MUX_8_13_port, Y(51)
                           => OUT_MUX_8_12_port, Y(52) => OUT_MUX_8_11_port, 
                           Y(53) => OUT_MUX_8_10_port, Y(54) => 
                           OUT_MUX_8_9_port, Y(55) => OUT_MUX_8_8_port, Y(56) 
                           => OUT_MUX_8_7_port, Y(57) => OUT_MUX_8_6_port, 
                           Y(58) => OUT_MUX_8_5_port, Y(59) => OUT_MUX_8_4_port
                           , Y(60) => OUT_MUX_8_3_port, Y(61) => 
                           OUT_MUX_8_2_port, Y(62) => OUT_MUX_8_1_port, Y(63) 
                           => OUT_MUX_8_0_port);
   MUXi_9 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_7 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_8_63_port, INPUT(65) => 
                           A_pos_shifted_by2_8_62_port, INPUT(66) => 
                           A_pos_shifted_by2_8_61_port, INPUT(67) => 
                           A_pos_shifted_by2_8_60_port, INPUT(68) => 
                           A_pos_shifted_by2_8_59_port, INPUT(69) => 
                           A_pos_shifted_by2_8_58_port, INPUT(70) => 
                           A_pos_shifted_by2_8_57_port, INPUT(71) => 
                           A_pos_shifted_by2_8_56_port, INPUT(72) => 
                           A_pos_shifted_by2_8_55_port, INPUT(73) => 
                           A_pos_shifted_by2_8_54_port, INPUT(74) => 
                           A_pos_shifted_by2_8_53_port, INPUT(75) => 
                           A_pos_shifted_by2_8_52_port, INPUT(76) => 
                           A_pos_shifted_by2_8_51_port, INPUT(77) => 
                           A_pos_shifted_by2_8_50_port, INPUT(78) => 
                           A_pos_shifted_by2_8_49_port, INPUT(79) => 
                           A_pos_shifted_by2_8_48_port, INPUT(80) => 
                           A_pos_shifted_by2_8_47_port, INPUT(81) => 
                           A_pos_shifted_by2_8_46_port, INPUT(82) => 
                           A_pos_shifted_by2_8_45_port, INPUT(83) => 
                           A_pos_shifted_by2_8_44_port, INPUT(84) => 
                           A_pos_shifted_by2_8_43_port, INPUT(85) => 
                           A_pos_shifted_by2_8_42_port, INPUT(86) => 
                           A_pos_shifted_by2_8_41_port, INPUT(87) => 
                           A_pos_shifted_by2_8_40_port, INPUT(88) => 
                           A_pos_shifted_by2_8_39_port, INPUT(89) => 
                           A_pos_shifted_by2_8_38_port, INPUT(90) => 
                           A_pos_shifted_by2_8_37_port, INPUT(91) => 
                           A_pos_shifted_by2_8_36_port, INPUT(92) => 
                           A_pos_shifted_by2_8_35_port, INPUT(93) => 
                           A_pos_shifted_by2_8_34_port, INPUT(94) => 
                           A_pos_shifted_by2_8_33_port, INPUT(95) => 
                           A_pos_shifted_by2_8_32_port, INPUT(96) => 
                           A_pos_shifted_by2_8_31_port, INPUT(97) => 
                           A_pos_shifted_by2_8_30_port, INPUT(98) => 
                           A_pos_shifted_by2_8_29_port, INPUT(99) => 
                           A_pos_shifted_by2_8_28_port, INPUT(100) => 
                           A_pos_shifted_by2_8_27_port, INPUT(101) => 
                           A_pos_shifted_by2_8_26_port, INPUT(102) => 
                           A_pos_shifted_by2_8_25_port, INPUT(103) => 
                           A_pos_shifted_by2_8_24_port, INPUT(104) => 
                           A_pos_shifted_by2_8_23_port, INPUT(105) => 
                           A_pos_shifted_by2_8_22_port, INPUT(106) => 
                           A_pos_shifted_by2_8_21_port, INPUT(107) => 
                           A_pos_shifted_by2_8_20_port, INPUT(108) => 
                           A_pos_shifted_by2_8_19_port, INPUT(109) => 
                           A_pos_shifted_by2_8_18_port, INPUT(110) => 
                           A_pos_shifted_by2_8_17_port, INPUT(111) => 
                           A_pos_shifted_by2_8_16_port, INPUT(112) => 
                           A_pos_shifted_by2_8_15_port, INPUT(113) => 
                           A_pos_shifted_by2_8_14_port, INPUT(114) => 
                           A_pos_shifted_by2_8_13_port, INPUT(115) => 
                           A_pos_shifted_by2_8_12_port, INPUT(116) => 
                           A_pos_shifted_by2_8_11_port, INPUT(117) => 
                           A_pos_shifted_by2_8_10_port, INPUT(118) => 
                           A_pos_shifted_by2_8_9_port, INPUT(119) => 
                           A_pos_shifted_by2_8_8_port, INPUT(120) => 
                           A_pos_shifted_by2_8_7_port, INPUT(121) => 
                           A_pos_shifted_by2_8_6_port, INPUT(122) => 
                           A_pos_shifted_by2_8_5_port, INPUT(123) => 
                           A_pos_shifted_by2_8_4_port, INPUT(124) => 
                           A_pos_shifted_by2_8_3_port, INPUT(125) => 
                           A_pos_shifted_by2_8_2_port, INPUT(126) => 
                           A_pos_shifted_by2_8_1_port, INPUT(127) => 
                           A_pos_shifted_by2_8_0_port, INPUT(128) => 
                           A_neg_shifted_by2_8_63_port, INPUT(129) => 
                           A_neg_shifted_by2_8_62_port, INPUT(130) => 
                           A_neg_shifted_by2_8_61_port, INPUT(131) => 
                           A_neg_shifted_by2_8_60_port, INPUT(132) => 
                           A_neg_shifted_by2_8_59_port, INPUT(133) => 
                           A_neg_shifted_by2_8_58_port, INPUT(134) => 
                           A_neg_shifted_by2_8_57_port, INPUT(135) => 
                           A_neg_shifted_by2_8_56_port, INPUT(136) => 
                           A_neg_shifted_by2_8_55_port, INPUT(137) => 
                           A_neg_shifted_by2_8_54_port, INPUT(138) => 
                           A_neg_shifted_by2_8_53_port, INPUT(139) => 
                           A_neg_shifted_by2_8_52_port, INPUT(140) => 
                           A_neg_shifted_by2_8_51_port, INPUT(141) => 
                           A_neg_shifted_by2_8_50_port, INPUT(142) => 
                           A_neg_shifted_by2_8_49_port, INPUT(143) => 
                           A_neg_shifted_by2_8_48_port, INPUT(144) => 
                           A_neg_shifted_by2_8_47_port, INPUT(145) => 
                           A_neg_shifted_by2_8_46_port, INPUT(146) => 
                           A_neg_shifted_by2_8_45_port, INPUT(147) => 
                           A_neg_shifted_by2_8_44_port, INPUT(148) => 
                           A_neg_shifted_by2_8_43_port, INPUT(149) => 
                           A_neg_shifted_by2_8_42_port, INPUT(150) => 
                           A_neg_shifted_by2_8_41_port, INPUT(151) => 
                           A_neg_shifted_by2_8_40_port, INPUT(152) => 
                           A_neg_shifted_by2_8_39_port, INPUT(153) => 
                           A_neg_shifted_by2_8_38_port, INPUT(154) => 
                           A_neg_shifted_by2_8_37_port, INPUT(155) => 
                           A_neg_shifted_by2_8_36_port, INPUT(156) => 
                           A_neg_shifted_by2_8_35_port, INPUT(157) => 
                           A_neg_shifted_by2_8_34_port, INPUT(158) => 
                           A_neg_shifted_by2_8_33_port, INPUT(159) => 
                           A_neg_shifted_by2_8_32_port, INPUT(160) => 
                           A_neg_shifted_by2_8_31_port, INPUT(161) => 
                           A_neg_shifted_by2_8_30_port, INPUT(162) => 
                           A_neg_shifted_by2_8_29_port, INPUT(163) => 
                           A_neg_shifted_by2_8_28_port, INPUT(164) => 
                           A_neg_shifted_by2_8_27_port, INPUT(165) => 
                           A_neg_shifted_by2_8_26_port, INPUT(166) => 
                           A_neg_shifted_by2_8_25_port, INPUT(167) => 
                           A_neg_shifted_by2_8_24_port, INPUT(168) => 
                           A_neg_shifted_by2_8_23_port, INPUT(169) => 
                           A_neg_shifted_by2_8_22_port, INPUT(170) => 
                           A_neg_shifted_by2_8_21_port, INPUT(171) => 
                           A_neg_shifted_by2_8_20_port, INPUT(172) => 
                           A_neg_shifted_by2_8_19_port, INPUT(173) => 
                           A_neg_shifted_by2_8_18_port, INPUT(174) => 
                           A_neg_shifted_by2_8_17_port, INPUT(175) => 
                           A_neg_shifted_by2_8_16_port, INPUT(176) => 
                           A_neg_shifted_by2_8_15_port, INPUT(177) => 
                           A_neg_shifted_by2_8_14_port, INPUT(178) => 
                           A_neg_shifted_by2_8_13_port, INPUT(179) => 
                           A_neg_shifted_by2_8_12_port, INPUT(180) => 
                           A_neg_shifted_by2_8_11_port, INPUT(181) => 
                           A_neg_shifted_by2_8_10_port, INPUT(182) => 
                           A_neg_shifted_by2_8_9_port, INPUT(183) => 
                           A_neg_shifted_by2_8_8_port, INPUT(184) => 
                           A_neg_shifted_by2_8_7_port, INPUT(185) => 
                           A_neg_shifted_by2_8_6_port, INPUT(186) => 
                           A_neg_shifted_by2_8_5_port, INPUT(187) => 
                           A_neg_shifted_by2_8_4_port, INPUT(188) => 
                           A_neg_shifted_by2_8_3_port, INPUT(189) => 
                           A_neg_shifted_by2_8_2_port, INPUT(190) => 
                           A_neg_shifted_by2_8_1_port, INPUT(191) => 
                           A_neg_shifted_by2_8_0_port, INPUT(192) => 
                           A_pos_shifted_by1_9_63_port, INPUT(193) => 
                           A_pos_shifted_by1_9_62_port, INPUT(194) => 
                           A_pos_shifted_by1_9_61_port, INPUT(195) => 
                           A_pos_shifted_by1_9_60_port, INPUT(196) => 
                           A_pos_shifted_by1_9_59_port, INPUT(197) => 
                           A_pos_shifted_by1_9_58_port, INPUT(198) => 
                           A_pos_shifted_by1_9_57_port, INPUT(199) => 
                           A_pos_shifted_by1_9_56_port, INPUT(200) => 
                           A_pos_shifted_by1_9_55_port, INPUT(201) => 
                           A_pos_shifted_by1_9_54_port, INPUT(202) => 
                           A_pos_shifted_by1_9_53_port, INPUT(203) => 
                           A_pos_shifted_by1_9_52_port, INPUT(204) => 
                           A_pos_shifted_by1_9_51_port, INPUT(205) => 
                           A_pos_shifted_by1_9_50_port, INPUT(206) => 
                           A_pos_shifted_by1_9_49_port, INPUT(207) => 
                           A_pos_shifted_by1_9_48_port, INPUT(208) => 
                           A_pos_shifted_by1_9_47_port, INPUT(209) => 
                           A_pos_shifted_by1_9_46_port, INPUT(210) => 
                           A_pos_shifted_by1_9_45_port, INPUT(211) => 
                           A_pos_shifted_by1_9_44_port, INPUT(212) => 
                           A_pos_shifted_by1_9_43_port, INPUT(213) => 
                           A_pos_shifted_by1_9_42_port, INPUT(214) => 
                           A_pos_shifted_by1_9_41_port, INPUT(215) => 
                           A_pos_shifted_by1_9_40_port, INPUT(216) => 
                           A_pos_shifted_by1_9_39_port, INPUT(217) => 
                           A_pos_shifted_by1_9_38_port, INPUT(218) => 
                           A_pos_shifted_by1_9_37_port, INPUT(219) => 
                           A_pos_shifted_by1_9_36_port, INPUT(220) => 
                           A_pos_shifted_by1_9_35_port, INPUT(221) => 
                           A_pos_shifted_by1_9_34_port, INPUT(222) => 
                           A_pos_shifted_by1_9_33_port, INPUT(223) => 
                           A_pos_shifted_by1_9_32_port, INPUT(224) => 
                           A_pos_shifted_by1_9_31_port, INPUT(225) => 
                           A_pos_shifted_by1_9_30_port, INPUT(226) => 
                           A_pos_shifted_by1_9_29_port, INPUT(227) => 
                           A_pos_shifted_by1_9_28_port, INPUT(228) => 
                           A_pos_shifted_by1_9_27_port, INPUT(229) => 
                           A_pos_shifted_by1_9_26_port, INPUT(230) => 
                           A_pos_shifted_by1_9_25_port, INPUT(231) => 
                           A_pos_shifted_by1_9_24_port, INPUT(232) => 
                           A_pos_shifted_by1_9_23_port, INPUT(233) => 
                           A_pos_shifted_by1_9_22_port, INPUT(234) => 
                           A_pos_shifted_by1_9_21_port, INPUT(235) => 
                           A_pos_shifted_by1_9_20_port, INPUT(236) => 
                           A_pos_shifted_by1_9_19_port, INPUT(237) => 
                           A_pos_shifted_by1_9_18_port, INPUT(238) => 
                           A_pos_shifted_by1_9_17_port, INPUT(239) => 
                           A_pos_shifted_by1_9_16_port, INPUT(240) => 
                           A_pos_shifted_by1_9_15_port, INPUT(241) => 
                           A_pos_shifted_by1_9_14_port, INPUT(242) => 
                           A_pos_shifted_by1_9_13_port, INPUT(243) => 
                           A_pos_shifted_by1_9_12_port, INPUT(244) => 
                           A_pos_shifted_by1_9_11_port, INPUT(245) => 
                           A_pos_shifted_by1_9_10_port, INPUT(246) => 
                           A_pos_shifted_by1_9_9_port, INPUT(247) => 
                           A_pos_shifted_by1_9_8_port, INPUT(248) => 
                           A_pos_shifted_by1_9_7_port, INPUT(249) => 
                           A_pos_shifted_by1_9_6_port, INPUT(250) => 
                           A_pos_shifted_by1_9_5_port, INPUT(251) => 
                           A_pos_shifted_by1_9_4_port, INPUT(252) => 
                           A_pos_shifted_by1_9_3_port, INPUT(253) => 
                           A_pos_shifted_by1_9_2_port, INPUT(254) => 
                           A_pos_shifted_by1_9_1_port, INPUT(255) => 
                           A_pos_shifted_by1_9_0_port, INPUT(256) => 
                           A_neg_shifted_by1_9_63_port, INPUT(257) => 
                           A_neg_shifted_by1_9_62_port, INPUT(258) => 
                           A_neg_shifted_by1_9_61_port, INPUT(259) => 
                           A_neg_shifted_by1_9_60_port, INPUT(260) => 
                           A_neg_shifted_by1_9_59_port, INPUT(261) => 
                           A_neg_shifted_by1_9_58_port, INPUT(262) => 
                           A_neg_shifted_by1_9_57_port, INPUT(263) => 
                           A_neg_shifted_by1_9_56_port, INPUT(264) => 
                           A_neg_shifted_by1_9_55_port, INPUT(265) => 
                           A_neg_shifted_by1_9_54_port, INPUT(266) => 
                           A_neg_shifted_by1_9_53_port, INPUT(267) => 
                           A_neg_shifted_by1_9_52_port, INPUT(268) => 
                           A_neg_shifted_by1_9_51_port, INPUT(269) => 
                           A_neg_shifted_by1_9_50_port, INPUT(270) => 
                           A_neg_shifted_by1_9_49_port, INPUT(271) => 
                           A_neg_shifted_by1_9_48_port, INPUT(272) => 
                           A_neg_shifted_by1_9_47_port, INPUT(273) => 
                           A_neg_shifted_by1_9_46_port, INPUT(274) => 
                           A_neg_shifted_by1_9_45_port, INPUT(275) => 
                           A_neg_shifted_by1_9_44_port, INPUT(276) => 
                           A_neg_shifted_by1_9_43_port, INPUT(277) => 
                           A_neg_shifted_by1_9_42_port, INPUT(278) => 
                           A_neg_shifted_by1_9_41_port, INPUT(279) => 
                           A_neg_shifted_by1_9_40_port, INPUT(280) => 
                           A_neg_shifted_by1_9_39_port, INPUT(281) => 
                           A_neg_shifted_by1_9_38_port, INPUT(282) => 
                           A_neg_shifted_by1_9_37_port, INPUT(283) => 
                           A_neg_shifted_by1_9_36_port, INPUT(284) => 
                           A_neg_shifted_by1_9_35_port, INPUT(285) => 
                           A_neg_shifted_by1_9_34_port, INPUT(286) => 
                           A_neg_shifted_by1_9_33_port, INPUT(287) => 
                           A_neg_shifted_by1_9_32_port, INPUT(288) => 
                           A_neg_shifted_by1_9_31_port, INPUT(289) => 
                           A_neg_shifted_by1_9_30_port, INPUT(290) => 
                           A_neg_shifted_by1_9_29_port, INPUT(291) => 
                           A_neg_shifted_by1_9_28_port, INPUT(292) => 
                           A_neg_shifted_by1_9_27_port, INPUT(293) => 
                           A_neg_shifted_by1_9_26_port, INPUT(294) => 
                           A_neg_shifted_by1_9_25_port, INPUT(295) => 
                           A_neg_shifted_by1_9_24_port, INPUT(296) => 
                           A_neg_shifted_by1_9_23_port, INPUT(297) => 
                           A_neg_shifted_by1_9_22_port, INPUT(298) => 
                           A_neg_shifted_by1_9_21_port, INPUT(299) => 
                           A_neg_shifted_by1_9_20_port, INPUT(300) => 
                           A_neg_shifted_by1_9_19_port, INPUT(301) => 
                           A_neg_shifted_by1_9_18_port, INPUT(302) => 
                           A_neg_shifted_by1_9_17_port, INPUT(303) => 
                           A_neg_shifted_by1_9_16_port, INPUT(304) => 
                           A_neg_shifted_by1_9_15_port, INPUT(305) => 
                           A_neg_shifted_by1_9_14_port, INPUT(306) => 
                           A_neg_shifted_by1_9_13_port, INPUT(307) => 
                           A_neg_shifted_by1_9_12_port, INPUT(308) => 
                           A_neg_shifted_by1_9_11_port, INPUT(309) => 
                           A_neg_shifted_by1_9_10_port, INPUT(310) => 
                           A_neg_shifted_by1_9_9_port, INPUT(311) => 
                           A_neg_shifted_by1_9_8_port, INPUT(312) => 
                           A_neg_shifted_by1_9_7_port, INPUT(313) => 
                           A_neg_shifted_by1_9_6_port, INPUT(314) => 
                           A_neg_shifted_by1_9_5_port, INPUT(315) => 
                           A_neg_shifted_by1_9_4_port, INPUT(316) => 
                           A_neg_shifted_by1_9_3_port, INPUT(317) => 
                           A_neg_shifted_by1_9_2_port, INPUT(318) => 
                           A_neg_shifted_by1_9_1_port, INPUT(319) => 
                           A_neg_shifted_by1_9_0_port, SEL(0) => 
                           selection_signal_9_2_port, SEL(1) => 
                           selection_signal_9_1_port, SEL(2) => 
                           selection_signal_9_0_port, Y(0) => OUT_MUX_9_63_port
                           , Y(1) => OUT_MUX_9_62_port, Y(2) => 
                           OUT_MUX_9_61_port, Y(3) => OUT_MUX_9_60_port, Y(4) 
                           => OUT_MUX_9_59_port, Y(5) => OUT_MUX_9_58_port, 
                           Y(6) => OUT_MUX_9_57_port, Y(7) => OUT_MUX_9_56_port
                           , Y(8) => OUT_MUX_9_55_port, Y(9) => 
                           OUT_MUX_9_54_port, Y(10) => OUT_MUX_9_53_port, Y(11)
                           => OUT_MUX_9_52_port, Y(12) => OUT_MUX_9_51_port, 
                           Y(13) => OUT_MUX_9_50_port, Y(14) => 
                           OUT_MUX_9_49_port, Y(15) => OUT_MUX_9_48_port, Y(16)
                           => OUT_MUX_9_47_port, Y(17) => OUT_MUX_9_46_port, 
                           Y(18) => OUT_MUX_9_45_port, Y(19) => 
                           OUT_MUX_9_44_port, Y(20) => OUT_MUX_9_43_port, Y(21)
                           => OUT_MUX_9_42_port, Y(22) => OUT_MUX_9_41_port, 
                           Y(23) => OUT_MUX_9_40_port, Y(24) => 
                           OUT_MUX_9_39_port, Y(25) => OUT_MUX_9_38_port, Y(26)
                           => OUT_MUX_9_37_port, Y(27) => OUT_MUX_9_36_port, 
                           Y(28) => OUT_MUX_9_35_port, Y(29) => 
                           OUT_MUX_9_34_port, Y(30) => OUT_MUX_9_33_port, Y(31)
                           => OUT_MUX_9_32_port, Y(32) => OUT_MUX_9_31_port, 
                           Y(33) => OUT_MUX_9_30_port, Y(34) => 
                           OUT_MUX_9_29_port, Y(35) => OUT_MUX_9_28_port, Y(36)
                           => OUT_MUX_9_27_port, Y(37) => OUT_MUX_9_26_port, 
                           Y(38) => OUT_MUX_9_25_port, Y(39) => 
                           OUT_MUX_9_24_port, Y(40) => OUT_MUX_9_23_port, Y(41)
                           => OUT_MUX_9_22_port, Y(42) => OUT_MUX_9_21_port, 
                           Y(43) => OUT_MUX_9_20_port, Y(44) => 
                           OUT_MUX_9_19_port, Y(45) => OUT_MUX_9_18_port, Y(46)
                           => OUT_MUX_9_17_port, Y(47) => OUT_MUX_9_16_port, 
                           Y(48) => OUT_MUX_9_15_port, Y(49) => 
                           OUT_MUX_9_14_port, Y(50) => OUT_MUX_9_13_port, Y(51)
                           => OUT_MUX_9_12_port, Y(52) => OUT_MUX_9_11_port, 
                           Y(53) => OUT_MUX_9_10_port, Y(54) => 
                           OUT_MUX_9_9_port, Y(55) => OUT_MUX_9_8_port, Y(56) 
                           => OUT_MUX_9_7_port, Y(57) => OUT_MUX_9_6_port, 
                           Y(58) => OUT_MUX_9_5_port, Y(59) => OUT_MUX_9_4_port
                           , Y(60) => OUT_MUX_9_3_port, Y(61) => 
                           OUT_MUX_9_2_port, Y(62) => OUT_MUX_9_1_port, Y(63) 
                           => OUT_MUX_9_0_port);
   MUXi_10 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_6 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_9_63_port, INPUT(65) => 
                           A_pos_shifted_by2_9_62_port, INPUT(66) => 
                           A_pos_shifted_by2_9_61_port, INPUT(67) => 
                           A_pos_shifted_by2_9_60_port, INPUT(68) => 
                           A_pos_shifted_by2_9_59_port, INPUT(69) => 
                           A_pos_shifted_by2_9_58_port, INPUT(70) => 
                           A_pos_shifted_by2_9_57_port, INPUT(71) => 
                           A_pos_shifted_by2_9_56_port, INPUT(72) => 
                           A_pos_shifted_by2_9_55_port, INPUT(73) => 
                           A_pos_shifted_by2_9_54_port, INPUT(74) => 
                           A_pos_shifted_by2_9_53_port, INPUT(75) => 
                           A_pos_shifted_by2_9_52_port, INPUT(76) => 
                           A_pos_shifted_by2_9_51_port, INPUT(77) => 
                           A_pos_shifted_by2_9_50_port, INPUT(78) => 
                           A_pos_shifted_by2_9_49_port, INPUT(79) => 
                           A_pos_shifted_by2_9_48_port, INPUT(80) => 
                           A_pos_shifted_by2_9_47_port, INPUT(81) => 
                           A_pos_shifted_by2_9_46_port, INPUT(82) => 
                           A_pos_shifted_by2_9_45_port, INPUT(83) => 
                           A_pos_shifted_by2_9_44_port, INPUT(84) => 
                           A_pos_shifted_by2_9_43_port, INPUT(85) => 
                           A_pos_shifted_by2_9_42_port, INPUT(86) => 
                           A_pos_shifted_by2_9_41_port, INPUT(87) => 
                           A_pos_shifted_by2_9_40_port, INPUT(88) => 
                           A_pos_shifted_by2_9_39_port, INPUT(89) => 
                           A_pos_shifted_by2_9_38_port, INPUT(90) => 
                           A_pos_shifted_by2_9_37_port, INPUT(91) => 
                           A_pos_shifted_by2_9_36_port, INPUT(92) => 
                           A_pos_shifted_by2_9_35_port, INPUT(93) => 
                           A_pos_shifted_by2_9_34_port, INPUT(94) => 
                           A_pos_shifted_by2_9_33_port, INPUT(95) => 
                           A_pos_shifted_by2_9_32_port, INPUT(96) => 
                           A_pos_shifted_by2_9_31_port, INPUT(97) => 
                           A_pos_shifted_by2_9_30_port, INPUT(98) => 
                           A_pos_shifted_by2_9_29_port, INPUT(99) => 
                           A_pos_shifted_by2_9_28_port, INPUT(100) => 
                           A_pos_shifted_by2_9_27_port, INPUT(101) => 
                           A_pos_shifted_by2_9_26_port, INPUT(102) => 
                           A_pos_shifted_by2_9_25_port, INPUT(103) => 
                           A_pos_shifted_by2_9_24_port, INPUT(104) => 
                           A_pos_shifted_by2_9_23_port, INPUT(105) => 
                           A_pos_shifted_by2_9_22_port, INPUT(106) => 
                           A_pos_shifted_by2_9_21_port, INPUT(107) => 
                           A_pos_shifted_by2_9_20_port, INPUT(108) => 
                           A_pos_shifted_by2_9_19_port, INPUT(109) => 
                           A_pos_shifted_by2_9_18_port, INPUT(110) => 
                           A_pos_shifted_by2_9_17_port, INPUT(111) => 
                           A_pos_shifted_by2_9_16_port, INPUT(112) => 
                           A_pos_shifted_by2_9_15_port, INPUT(113) => 
                           A_pos_shifted_by2_9_14_port, INPUT(114) => 
                           A_pos_shifted_by2_9_13_port, INPUT(115) => 
                           A_pos_shifted_by2_9_12_port, INPUT(116) => 
                           A_pos_shifted_by2_9_11_port, INPUT(117) => 
                           A_pos_shifted_by2_9_10_port, INPUT(118) => 
                           A_pos_shifted_by2_9_9_port, INPUT(119) => 
                           A_pos_shifted_by2_9_8_port, INPUT(120) => 
                           A_pos_shifted_by2_9_7_port, INPUT(121) => 
                           A_pos_shifted_by2_9_6_port, INPUT(122) => 
                           A_pos_shifted_by2_9_5_port, INPUT(123) => 
                           A_pos_shifted_by2_9_4_port, INPUT(124) => 
                           A_pos_shifted_by2_9_3_port, INPUT(125) => 
                           A_pos_shifted_by2_9_2_port, INPUT(126) => 
                           A_pos_shifted_by2_9_1_port, INPUT(127) => 
                           A_pos_shifted_by2_9_0_port, INPUT(128) => 
                           A_neg_shifted_by2_9_63_port, INPUT(129) => 
                           A_neg_shifted_by2_9_62_port, INPUT(130) => 
                           A_neg_shifted_by2_9_61_port, INPUT(131) => 
                           A_neg_shifted_by2_9_60_port, INPUT(132) => 
                           A_neg_shifted_by2_9_59_port, INPUT(133) => 
                           A_neg_shifted_by2_9_58_port, INPUT(134) => 
                           A_neg_shifted_by2_9_57_port, INPUT(135) => 
                           A_neg_shifted_by2_9_56_port, INPUT(136) => 
                           A_neg_shifted_by2_9_55_port, INPUT(137) => 
                           A_neg_shifted_by2_9_54_port, INPUT(138) => 
                           A_neg_shifted_by2_9_53_port, INPUT(139) => 
                           A_neg_shifted_by2_9_52_port, INPUT(140) => 
                           A_neg_shifted_by2_9_51_port, INPUT(141) => 
                           A_neg_shifted_by2_9_50_port, INPUT(142) => 
                           A_neg_shifted_by2_9_49_port, INPUT(143) => 
                           A_neg_shifted_by2_9_48_port, INPUT(144) => 
                           A_neg_shifted_by2_9_47_port, INPUT(145) => 
                           A_neg_shifted_by2_9_46_port, INPUT(146) => 
                           A_neg_shifted_by2_9_45_port, INPUT(147) => 
                           A_neg_shifted_by2_9_44_port, INPUT(148) => 
                           A_neg_shifted_by2_9_43_port, INPUT(149) => 
                           A_neg_shifted_by2_9_42_port, INPUT(150) => 
                           A_neg_shifted_by2_9_41_port, INPUT(151) => 
                           A_neg_shifted_by2_9_40_port, INPUT(152) => 
                           A_neg_shifted_by2_9_39_port, INPUT(153) => 
                           A_neg_shifted_by2_9_38_port, INPUT(154) => 
                           A_neg_shifted_by2_9_37_port, INPUT(155) => 
                           A_neg_shifted_by2_9_36_port, INPUT(156) => 
                           A_neg_shifted_by2_9_35_port, INPUT(157) => 
                           A_neg_shifted_by2_9_34_port, INPUT(158) => 
                           A_neg_shifted_by2_9_33_port, INPUT(159) => 
                           A_neg_shifted_by2_9_32_port, INPUT(160) => 
                           A_neg_shifted_by2_9_31_port, INPUT(161) => 
                           A_neg_shifted_by2_9_30_port, INPUT(162) => 
                           A_neg_shifted_by2_9_29_port, INPUT(163) => 
                           A_neg_shifted_by2_9_28_port, INPUT(164) => 
                           A_neg_shifted_by2_9_27_port, INPUT(165) => 
                           A_neg_shifted_by2_9_26_port, INPUT(166) => 
                           A_neg_shifted_by2_9_25_port, INPUT(167) => 
                           A_neg_shifted_by2_9_24_port, INPUT(168) => 
                           A_neg_shifted_by2_9_23_port, INPUT(169) => 
                           A_neg_shifted_by2_9_22_port, INPUT(170) => 
                           A_neg_shifted_by2_9_21_port, INPUT(171) => 
                           A_neg_shifted_by2_9_20_port, INPUT(172) => 
                           A_neg_shifted_by2_9_19_port, INPUT(173) => 
                           A_neg_shifted_by2_9_18_port, INPUT(174) => 
                           A_neg_shifted_by2_9_17_port, INPUT(175) => 
                           A_neg_shifted_by2_9_16_port, INPUT(176) => 
                           A_neg_shifted_by2_9_15_port, INPUT(177) => 
                           A_neg_shifted_by2_9_14_port, INPUT(178) => 
                           A_neg_shifted_by2_9_13_port, INPUT(179) => 
                           A_neg_shifted_by2_9_12_port, INPUT(180) => 
                           A_neg_shifted_by2_9_11_port, INPUT(181) => 
                           A_neg_shifted_by2_9_10_port, INPUT(182) => 
                           A_neg_shifted_by2_9_9_port, INPUT(183) => 
                           A_neg_shifted_by2_9_8_port, INPUT(184) => 
                           A_neg_shifted_by2_9_7_port, INPUT(185) => 
                           A_neg_shifted_by2_9_6_port, INPUT(186) => 
                           A_neg_shifted_by2_9_5_port, INPUT(187) => 
                           A_neg_shifted_by2_9_4_port, INPUT(188) => 
                           A_neg_shifted_by2_9_3_port, INPUT(189) => 
                           A_neg_shifted_by2_9_2_port, INPUT(190) => 
                           A_neg_shifted_by2_9_1_port, INPUT(191) => 
                           A_neg_shifted_by2_9_0_port, INPUT(192) => 
                           A_pos_shifted_by1_10_63_port, INPUT(193) => 
                           A_pos_shifted_by1_10_62_port, INPUT(194) => 
                           A_pos_shifted_by1_10_61_port, INPUT(195) => 
                           A_pos_shifted_by1_10_60_port, INPUT(196) => 
                           A_pos_shifted_by1_10_59_port, INPUT(197) => 
                           A_pos_shifted_by1_10_58_port, INPUT(198) => 
                           A_pos_shifted_by1_10_57_port, INPUT(199) => 
                           A_pos_shifted_by1_10_56_port, INPUT(200) => 
                           A_pos_shifted_by1_10_55_port, INPUT(201) => 
                           A_pos_shifted_by1_10_54_port, INPUT(202) => 
                           A_pos_shifted_by1_10_53_port, INPUT(203) => 
                           A_pos_shifted_by1_10_52_port, INPUT(204) => 
                           A_pos_shifted_by1_10_51_port, INPUT(205) => 
                           A_pos_shifted_by1_10_50_port, INPUT(206) => 
                           A_pos_shifted_by1_10_49_port, INPUT(207) => 
                           A_pos_shifted_by1_10_48_port, INPUT(208) => 
                           A_pos_shifted_by1_10_47_port, INPUT(209) => 
                           A_pos_shifted_by1_10_46_port, INPUT(210) => 
                           A_pos_shifted_by1_10_45_port, INPUT(211) => 
                           A_pos_shifted_by1_10_44_port, INPUT(212) => 
                           A_pos_shifted_by1_10_43_port, INPUT(213) => 
                           A_pos_shifted_by1_10_42_port, INPUT(214) => 
                           A_pos_shifted_by1_10_41_port, INPUT(215) => 
                           A_pos_shifted_by1_10_40_port, INPUT(216) => 
                           A_pos_shifted_by1_10_39_port, INPUT(217) => 
                           A_pos_shifted_by1_10_38_port, INPUT(218) => 
                           A_pos_shifted_by1_10_37_port, INPUT(219) => 
                           A_pos_shifted_by1_10_36_port, INPUT(220) => 
                           A_pos_shifted_by1_10_35_port, INPUT(221) => 
                           A_pos_shifted_by1_10_34_port, INPUT(222) => 
                           A_pos_shifted_by1_10_33_port, INPUT(223) => 
                           A_pos_shifted_by1_10_32_port, INPUT(224) => 
                           A_pos_shifted_by1_10_31_port, INPUT(225) => 
                           A_pos_shifted_by1_10_30_port, INPUT(226) => 
                           A_pos_shifted_by1_10_29_port, INPUT(227) => 
                           A_pos_shifted_by1_10_28_port, INPUT(228) => 
                           A_pos_shifted_by1_10_27_port, INPUT(229) => 
                           A_pos_shifted_by1_10_26_port, INPUT(230) => 
                           A_pos_shifted_by1_10_25_port, INPUT(231) => 
                           A_pos_shifted_by1_10_24_port, INPUT(232) => 
                           A_pos_shifted_by1_10_23_port, INPUT(233) => 
                           A_pos_shifted_by1_10_22_port, INPUT(234) => 
                           A_pos_shifted_by1_10_21_port, INPUT(235) => 
                           A_pos_shifted_by1_10_20_port, INPUT(236) => 
                           A_pos_shifted_by1_10_19_port, INPUT(237) => 
                           A_pos_shifted_by1_10_18_port, INPUT(238) => 
                           A_pos_shifted_by1_10_17_port, INPUT(239) => 
                           A_pos_shifted_by1_10_16_port, INPUT(240) => 
                           A_pos_shifted_by1_10_15_port, INPUT(241) => 
                           A_pos_shifted_by1_10_14_port, INPUT(242) => 
                           A_pos_shifted_by1_10_13_port, INPUT(243) => 
                           A_pos_shifted_by1_10_12_port, INPUT(244) => 
                           A_pos_shifted_by1_10_11_port, INPUT(245) => 
                           A_pos_shifted_by1_10_10_port, INPUT(246) => 
                           A_pos_shifted_by1_10_9_port, INPUT(247) => 
                           A_pos_shifted_by1_10_8_port, INPUT(248) => 
                           A_pos_shifted_by1_10_7_port, INPUT(249) => 
                           A_pos_shifted_by1_10_6_port, INPUT(250) => 
                           A_pos_shifted_by1_10_5_port, INPUT(251) => 
                           A_pos_shifted_by1_10_4_port, INPUT(252) => 
                           A_pos_shifted_by1_10_3_port, INPUT(253) => 
                           A_pos_shifted_by1_10_2_port, INPUT(254) => 
                           A_pos_shifted_by1_10_1_port, INPUT(255) => 
                           A_pos_shifted_by1_10_0_port, INPUT(256) => 
                           A_neg_shifted_by1_10_63_port, INPUT(257) => 
                           A_neg_shifted_by1_10_62_port, INPUT(258) => 
                           A_neg_shifted_by1_10_61_port, INPUT(259) => 
                           A_neg_shifted_by1_10_60_port, INPUT(260) => 
                           A_neg_shifted_by1_10_59_port, INPUT(261) => 
                           A_neg_shifted_by1_10_58_port, INPUT(262) => 
                           A_neg_shifted_by1_10_57_port, INPUT(263) => 
                           A_neg_shifted_by1_10_56_port, INPUT(264) => 
                           A_neg_shifted_by1_10_55_port, INPUT(265) => 
                           A_neg_shifted_by1_10_54_port, INPUT(266) => 
                           A_neg_shifted_by1_10_53_port, INPUT(267) => 
                           A_neg_shifted_by1_10_52_port, INPUT(268) => 
                           A_neg_shifted_by1_10_51_port, INPUT(269) => 
                           A_neg_shifted_by1_10_50_port, INPUT(270) => 
                           A_neg_shifted_by1_10_49_port, INPUT(271) => 
                           A_neg_shifted_by1_10_48_port, INPUT(272) => 
                           A_neg_shifted_by1_10_47_port, INPUT(273) => 
                           A_neg_shifted_by1_10_46_port, INPUT(274) => 
                           A_neg_shifted_by1_10_45_port, INPUT(275) => 
                           A_neg_shifted_by1_10_44_port, INPUT(276) => 
                           A_neg_shifted_by1_10_43_port, INPUT(277) => 
                           A_neg_shifted_by1_10_42_port, INPUT(278) => 
                           A_neg_shifted_by1_10_41_port, INPUT(279) => 
                           A_neg_shifted_by1_10_40_port, INPUT(280) => 
                           A_neg_shifted_by1_10_39_port, INPUT(281) => 
                           A_neg_shifted_by1_10_38_port, INPUT(282) => 
                           A_neg_shifted_by1_10_37_port, INPUT(283) => 
                           A_neg_shifted_by1_10_36_port, INPUT(284) => 
                           A_neg_shifted_by1_10_35_port, INPUT(285) => 
                           A_neg_shifted_by1_10_34_port, INPUT(286) => 
                           A_neg_shifted_by1_10_33_port, INPUT(287) => 
                           A_neg_shifted_by1_10_32_port, INPUT(288) => 
                           A_neg_shifted_by1_10_31_port, INPUT(289) => 
                           A_neg_shifted_by1_10_30_port, INPUT(290) => 
                           A_neg_shifted_by1_10_29_port, INPUT(291) => 
                           A_neg_shifted_by1_10_28_port, INPUT(292) => 
                           A_neg_shifted_by1_10_27_port, INPUT(293) => 
                           A_neg_shifted_by1_10_26_port, INPUT(294) => 
                           A_neg_shifted_by1_10_25_port, INPUT(295) => 
                           A_neg_shifted_by1_10_24_port, INPUT(296) => 
                           A_neg_shifted_by1_10_23_port, INPUT(297) => 
                           A_neg_shifted_by1_10_22_port, INPUT(298) => 
                           A_neg_shifted_by1_10_21_port, INPUT(299) => 
                           A_neg_shifted_by1_10_20_port, INPUT(300) => 
                           A_neg_shifted_by1_10_19_port, INPUT(301) => 
                           A_neg_shifted_by1_10_18_port, INPUT(302) => 
                           A_neg_shifted_by1_10_17_port, INPUT(303) => 
                           A_neg_shifted_by1_10_16_port, INPUT(304) => 
                           A_neg_shifted_by1_10_15_port, INPUT(305) => 
                           A_neg_shifted_by1_10_14_port, INPUT(306) => 
                           A_neg_shifted_by1_10_13_port, INPUT(307) => 
                           A_neg_shifted_by1_10_12_port, INPUT(308) => 
                           A_neg_shifted_by1_10_11_port, INPUT(309) => 
                           A_neg_shifted_by1_10_10_port, INPUT(310) => 
                           A_neg_shifted_by1_10_9_port, INPUT(311) => 
                           A_neg_shifted_by1_10_8_port, INPUT(312) => 
                           A_neg_shifted_by1_10_7_port, INPUT(313) => 
                           A_neg_shifted_by1_10_6_port, INPUT(314) => 
                           A_neg_shifted_by1_10_5_port, INPUT(315) => 
                           A_neg_shifted_by1_10_4_port, INPUT(316) => 
                           A_neg_shifted_by1_10_3_port, INPUT(317) => 
                           A_neg_shifted_by1_10_2_port, INPUT(318) => 
                           A_neg_shifted_by1_10_1_port, INPUT(319) => 
                           A_neg_shifted_by1_10_0_port, SEL(0) => 
                           selection_signal_10_2_port, SEL(1) => 
                           selection_signal_10_1_port, SEL(2) => 
                           selection_signal_10_0_port, Y(0) => 
                           OUT_MUX_10_63_port, Y(1) => OUT_MUX_10_62_port, Y(2)
                           => OUT_MUX_10_61_port, Y(3) => OUT_MUX_10_60_port, 
                           Y(4) => OUT_MUX_10_59_port, Y(5) => 
                           OUT_MUX_10_58_port, Y(6) => OUT_MUX_10_57_port, Y(7)
                           => OUT_MUX_10_56_port, Y(8) => OUT_MUX_10_55_port, 
                           Y(9) => OUT_MUX_10_54_port, Y(10) => 
                           OUT_MUX_10_53_port, Y(11) => OUT_MUX_10_52_port, 
                           Y(12) => OUT_MUX_10_51_port, Y(13) => 
                           OUT_MUX_10_50_port, Y(14) => OUT_MUX_10_49_port, 
                           Y(15) => OUT_MUX_10_48_port, Y(16) => 
                           OUT_MUX_10_47_port, Y(17) => OUT_MUX_10_46_port, 
                           Y(18) => OUT_MUX_10_45_port, Y(19) => 
                           OUT_MUX_10_44_port, Y(20) => OUT_MUX_10_43_port, 
                           Y(21) => OUT_MUX_10_42_port, Y(22) => 
                           OUT_MUX_10_41_port, Y(23) => OUT_MUX_10_40_port, 
                           Y(24) => OUT_MUX_10_39_port, Y(25) => 
                           OUT_MUX_10_38_port, Y(26) => OUT_MUX_10_37_port, 
                           Y(27) => OUT_MUX_10_36_port, Y(28) => 
                           OUT_MUX_10_35_port, Y(29) => OUT_MUX_10_34_port, 
                           Y(30) => OUT_MUX_10_33_port, Y(31) => 
                           OUT_MUX_10_32_port, Y(32) => OUT_MUX_10_31_port, 
                           Y(33) => OUT_MUX_10_30_port, Y(34) => 
                           OUT_MUX_10_29_port, Y(35) => OUT_MUX_10_28_port, 
                           Y(36) => OUT_MUX_10_27_port, Y(37) => 
                           OUT_MUX_10_26_port, Y(38) => OUT_MUX_10_25_port, 
                           Y(39) => OUT_MUX_10_24_port, Y(40) => 
                           OUT_MUX_10_23_port, Y(41) => OUT_MUX_10_22_port, 
                           Y(42) => OUT_MUX_10_21_port, Y(43) => 
                           OUT_MUX_10_20_port, Y(44) => OUT_MUX_10_19_port, 
                           Y(45) => OUT_MUX_10_18_port, Y(46) => 
                           OUT_MUX_10_17_port, Y(47) => OUT_MUX_10_16_port, 
                           Y(48) => OUT_MUX_10_15_port, Y(49) => 
                           OUT_MUX_10_14_port, Y(50) => OUT_MUX_10_13_port, 
                           Y(51) => OUT_MUX_10_12_port, Y(52) => 
                           OUT_MUX_10_11_port, Y(53) => OUT_MUX_10_10_port, 
                           Y(54) => OUT_MUX_10_9_port, Y(55) => 
                           OUT_MUX_10_8_port, Y(56) => OUT_MUX_10_7_port, Y(57)
                           => OUT_MUX_10_6_port, Y(58) => OUT_MUX_10_5_port, 
                           Y(59) => OUT_MUX_10_4_port, Y(60) => 
                           OUT_MUX_10_3_port, Y(61) => OUT_MUX_10_2_port, Y(62)
                           => OUT_MUX_10_1_port, Y(63) => OUT_MUX_10_0_port);
   MUXi_11 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_5 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_10_63_port, INPUT(65) => 
                           A_pos_shifted_by2_10_62_port, INPUT(66) => 
                           A_pos_shifted_by2_10_61_port, INPUT(67) => 
                           A_pos_shifted_by2_10_60_port, INPUT(68) => 
                           A_pos_shifted_by2_10_59_port, INPUT(69) => 
                           A_pos_shifted_by2_10_58_port, INPUT(70) => 
                           A_pos_shifted_by2_10_57_port, INPUT(71) => 
                           A_pos_shifted_by2_10_56_port, INPUT(72) => 
                           A_pos_shifted_by2_10_55_port, INPUT(73) => 
                           A_pos_shifted_by2_10_54_port, INPUT(74) => 
                           A_pos_shifted_by2_10_53_port, INPUT(75) => 
                           A_pos_shifted_by2_10_52_port, INPUT(76) => 
                           A_pos_shifted_by2_10_51_port, INPUT(77) => 
                           A_pos_shifted_by2_10_50_port, INPUT(78) => 
                           A_pos_shifted_by2_10_49_port, INPUT(79) => 
                           A_pos_shifted_by2_10_48_port, INPUT(80) => 
                           A_pos_shifted_by2_10_47_port, INPUT(81) => 
                           A_pos_shifted_by2_10_46_port, INPUT(82) => 
                           A_pos_shifted_by2_10_45_port, INPUT(83) => 
                           A_pos_shifted_by2_10_44_port, INPUT(84) => 
                           A_pos_shifted_by2_10_43_port, INPUT(85) => 
                           A_pos_shifted_by2_10_42_port, INPUT(86) => 
                           A_pos_shifted_by2_10_41_port, INPUT(87) => 
                           A_pos_shifted_by2_10_40_port, INPUT(88) => 
                           A_pos_shifted_by2_10_39_port, INPUT(89) => 
                           A_pos_shifted_by2_10_38_port, INPUT(90) => 
                           A_pos_shifted_by2_10_37_port, INPUT(91) => 
                           A_pos_shifted_by2_10_36_port, INPUT(92) => 
                           A_pos_shifted_by2_10_35_port, INPUT(93) => 
                           A_pos_shifted_by2_10_34_port, INPUT(94) => 
                           A_pos_shifted_by2_10_33_port, INPUT(95) => 
                           A_pos_shifted_by2_10_32_port, INPUT(96) => 
                           A_pos_shifted_by2_10_31_port, INPUT(97) => 
                           A_pos_shifted_by2_10_30_port, INPUT(98) => 
                           A_pos_shifted_by2_10_29_port, INPUT(99) => 
                           A_pos_shifted_by2_10_28_port, INPUT(100) => 
                           A_pos_shifted_by2_10_27_port, INPUT(101) => 
                           A_pos_shifted_by2_10_26_port, INPUT(102) => 
                           A_pos_shifted_by2_10_25_port, INPUT(103) => 
                           A_pos_shifted_by2_10_24_port, INPUT(104) => 
                           A_pos_shifted_by2_10_23_port, INPUT(105) => 
                           A_pos_shifted_by2_10_22_port, INPUT(106) => 
                           A_pos_shifted_by2_10_21_port, INPUT(107) => 
                           A_pos_shifted_by2_10_20_port, INPUT(108) => 
                           A_pos_shifted_by2_10_19_port, INPUT(109) => 
                           A_pos_shifted_by2_10_18_port, INPUT(110) => 
                           A_pos_shifted_by2_10_17_port, INPUT(111) => 
                           A_pos_shifted_by2_10_16_port, INPUT(112) => 
                           A_pos_shifted_by2_10_15_port, INPUT(113) => 
                           A_pos_shifted_by2_10_14_port, INPUT(114) => 
                           A_pos_shifted_by2_10_13_port, INPUT(115) => 
                           A_pos_shifted_by2_10_12_port, INPUT(116) => 
                           A_pos_shifted_by2_10_11_port, INPUT(117) => 
                           A_pos_shifted_by2_10_10_port, INPUT(118) => 
                           A_pos_shifted_by2_10_9_port, INPUT(119) => 
                           A_pos_shifted_by2_10_8_port, INPUT(120) => 
                           A_pos_shifted_by2_10_7_port, INPUT(121) => 
                           A_pos_shifted_by2_10_6_port, INPUT(122) => 
                           A_pos_shifted_by2_10_5_port, INPUT(123) => 
                           A_pos_shifted_by2_10_4_port, INPUT(124) => 
                           A_pos_shifted_by2_10_3_port, INPUT(125) => 
                           A_pos_shifted_by2_10_2_port, INPUT(126) => 
                           A_pos_shifted_by2_10_1_port, INPUT(127) => 
                           A_pos_shifted_by2_10_0_port, INPUT(128) => 
                           A_neg_shifted_by2_10_63_port, INPUT(129) => 
                           A_neg_shifted_by2_10_62_port, INPUT(130) => 
                           A_neg_shifted_by2_10_61_port, INPUT(131) => 
                           A_neg_shifted_by2_10_60_port, INPUT(132) => 
                           A_neg_shifted_by2_10_59_port, INPUT(133) => 
                           A_neg_shifted_by2_10_58_port, INPUT(134) => 
                           A_neg_shifted_by2_10_57_port, INPUT(135) => 
                           A_neg_shifted_by2_10_56_port, INPUT(136) => 
                           A_neg_shifted_by2_10_55_port, INPUT(137) => 
                           A_neg_shifted_by2_10_54_port, INPUT(138) => 
                           A_neg_shifted_by2_10_53_port, INPUT(139) => 
                           A_neg_shifted_by2_10_52_port, INPUT(140) => 
                           A_neg_shifted_by2_10_51_port, INPUT(141) => 
                           A_neg_shifted_by2_10_50_port, INPUT(142) => 
                           A_neg_shifted_by2_10_49_port, INPUT(143) => 
                           A_neg_shifted_by2_10_48_port, INPUT(144) => 
                           A_neg_shifted_by2_10_47_port, INPUT(145) => 
                           A_neg_shifted_by2_10_46_port, INPUT(146) => 
                           A_neg_shifted_by2_10_45_port, INPUT(147) => 
                           A_neg_shifted_by2_10_44_port, INPUT(148) => 
                           A_neg_shifted_by2_10_43_port, INPUT(149) => 
                           A_neg_shifted_by2_10_42_port, INPUT(150) => 
                           A_neg_shifted_by2_10_41_port, INPUT(151) => 
                           A_neg_shifted_by2_10_40_port, INPUT(152) => 
                           A_neg_shifted_by2_10_39_port, INPUT(153) => 
                           A_neg_shifted_by2_10_38_port, INPUT(154) => 
                           A_neg_shifted_by2_10_37_port, INPUT(155) => 
                           A_neg_shifted_by2_10_36_port, INPUT(156) => 
                           A_neg_shifted_by2_10_35_port, INPUT(157) => 
                           A_neg_shifted_by2_10_34_port, INPUT(158) => 
                           A_neg_shifted_by2_10_33_port, INPUT(159) => 
                           A_neg_shifted_by2_10_32_port, INPUT(160) => 
                           A_neg_shifted_by2_10_31_port, INPUT(161) => 
                           A_neg_shifted_by2_10_30_port, INPUT(162) => 
                           A_neg_shifted_by2_10_29_port, INPUT(163) => 
                           A_neg_shifted_by2_10_28_port, INPUT(164) => 
                           A_neg_shifted_by2_10_27_port, INPUT(165) => 
                           A_neg_shifted_by2_10_26_port, INPUT(166) => 
                           A_neg_shifted_by2_10_25_port, INPUT(167) => 
                           A_neg_shifted_by2_10_24_port, INPUT(168) => 
                           A_neg_shifted_by2_10_23_port, INPUT(169) => 
                           A_neg_shifted_by2_10_22_port, INPUT(170) => 
                           A_neg_shifted_by2_10_21_port, INPUT(171) => 
                           A_neg_shifted_by2_10_20_port, INPUT(172) => 
                           A_neg_shifted_by2_10_19_port, INPUT(173) => 
                           A_neg_shifted_by2_10_18_port, INPUT(174) => 
                           A_neg_shifted_by2_10_17_port, INPUT(175) => 
                           A_neg_shifted_by2_10_16_port, INPUT(176) => 
                           A_neg_shifted_by2_10_15_port, INPUT(177) => 
                           A_neg_shifted_by2_10_14_port, INPUT(178) => 
                           A_neg_shifted_by2_10_13_port, INPUT(179) => 
                           A_neg_shifted_by2_10_12_port, INPUT(180) => 
                           A_neg_shifted_by2_10_11_port, INPUT(181) => 
                           A_neg_shifted_by2_10_10_port, INPUT(182) => 
                           A_neg_shifted_by2_10_9_port, INPUT(183) => 
                           A_neg_shifted_by2_10_8_port, INPUT(184) => 
                           A_neg_shifted_by2_10_7_port, INPUT(185) => 
                           A_neg_shifted_by2_10_6_port, INPUT(186) => 
                           A_neg_shifted_by2_10_5_port, INPUT(187) => 
                           A_neg_shifted_by2_10_4_port, INPUT(188) => 
                           A_neg_shifted_by2_10_3_port, INPUT(189) => 
                           A_neg_shifted_by2_10_2_port, INPUT(190) => 
                           A_neg_shifted_by2_10_1_port, INPUT(191) => 
                           A_neg_shifted_by2_10_0_port, INPUT(192) => 
                           A_pos_shifted_by1_11_63_port, INPUT(193) => 
                           A_pos_shifted_by1_11_62_port, INPUT(194) => 
                           A_pos_shifted_by1_11_61_port, INPUT(195) => 
                           A_pos_shifted_by1_11_60_port, INPUT(196) => 
                           A_pos_shifted_by1_11_59_port, INPUT(197) => 
                           A_pos_shifted_by1_11_58_port, INPUT(198) => 
                           A_pos_shifted_by1_11_57_port, INPUT(199) => 
                           A_pos_shifted_by1_11_56_port, INPUT(200) => 
                           A_pos_shifted_by1_11_55_port, INPUT(201) => 
                           A_pos_shifted_by1_11_54_port, INPUT(202) => 
                           A_pos_shifted_by1_11_53_port, INPUT(203) => 
                           A_pos_shifted_by1_11_52_port, INPUT(204) => 
                           A_pos_shifted_by1_11_51_port, INPUT(205) => 
                           A_pos_shifted_by1_11_50_port, INPUT(206) => 
                           A_pos_shifted_by1_11_49_port, INPUT(207) => 
                           A_pos_shifted_by1_11_48_port, INPUT(208) => 
                           A_pos_shifted_by1_11_47_port, INPUT(209) => 
                           A_pos_shifted_by1_11_46_port, INPUT(210) => 
                           A_pos_shifted_by1_11_45_port, INPUT(211) => 
                           A_pos_shifted_by1_11_44_port, INPUT(212) => 
                           A_pos_shifted_by1_11_43_port, INPUT(213) => 
                           A_pos_shifted_by1_11_42_port, INPUT(214) => 
                           A_pos_shifted_by1_11_41_port, INPUT(215) => 
                           A_pos_shifted_by1_11_40_port, INPUT(216) => 
                           A_pos_shifted_by1_11_39_port, INPUT(217) => 
                           A_pos_shifted_by1_11_38_port, INPUT(218) => 
                           A_pos_shifted_by1_11_37_port, INPUT(219) => 
                           A_pos_shifted_by1_11_36_port, INPUT(220) => 
                           A_pos_shifted_by1_11_35_port, INPUT(221) => 
                           A_pos_shifted_by1_11_34_port, INPUT(222) => 
                           A_pos_shifted_by1_11_33_port, INPUT(223) => 
                           A_pos_shifted_by1_11_32_port, INPUT(224) => 
                           A_pos_shifted_by1_11_31_port, INPUT(225) => 
                           A_pos_shifted_by1_11_30_port, INPUT(226) => 
                           A_pos_shifted_by1_11_29_port, INPUT(227) => 
                           A_pos_shifted_by1_11_28_port, INPUT(228) => 
                           A_pos_shifted_by1_11_27_port, INPUT(229) => 
                           A_pos_shifted_by1_11_26_port, INPUT(230) => 
                           A_pos_shifted_by1_11_25_port, INPUT(231) => 
                           A_pos_shifted_by1_11_24_port, INPUT(232) => 
                           A_pos_shifted_by1_11_23_port, INPUT(233) => 
                           A_pos_shifted_by1_11_22_port, INPUT(234) => 
                           A_pos_shifted_by1_11_21_port, INPUT(235) => 
                           A_pos_shifted_by1_11_20_port, INPUT(236) => 
                           A_pos_shifted_by1_11_19_port, INPUT(237) => 
                           A_pos_shifted_by1_11_18_port, INPUT(238) => 
                           A_pos_shifted_by1_11_17_port, INPUT(239) => 
                           A_pos_shifted_by1_11_16_port, INPUT(240) => 
                           A_pos_shifted_by1_11_15_port, INPUT(241) => 
                           A_pos_shifted_by1_11_14_port, INPUT(242) => 
                           A_pos_shifted_by1_11_13_port, INPUT(243) => 
                           A_pos_shifted_by1_11_12_port, INPUT(244) => 
                           A_pos_shifted_by1_11_11_port, INPUT(245) => 
                           A_pos_shifted_by1_11_10_port, INPUT(246) => 
                           A_pos_shifted_by1_11_9_port, INPUT(247) => 
                           A_pos_shifted_by1_11_8_port, INPUT(248) => 
                           A_pos_shifted_by1_11_7_port, INPUT(249) => 
                           A_pos_shifted_by1_11_6_port, INPUT(250) => 
                           A_pos_shifted_by1_11_5_port, INPUT(251) => 
                           A_pos_shifted_by1_11_4_port, INPUT(252) => 
                           A_pos_shifted_by1_11_3_port, INPUT(253) => 
                           A_pos_shifted_by1_11_2_port, INPUT(254) => 
                           A_pos_shifted_by1_11_1_port, INPUT(255) => 
                           A_pos_shifted_by1_11_0_port, INPUT(256) => 
                           A_neg_shifted_by1_11_63_port, INPUT(257) => 
                           A_neg_shifted_by1_11_62_port, INPUT(258) => 
                           A_neg_shifted_by1_11_61_port, INPUT(259) => 
                           A_neg_shifted_by1_11_60_port, INPUT(260) => 
                           A_neg_shifted_by1_11_59_port, INPUT(261) => 
                           A_neg_shifted_by1_11_58_port, INPUT(262) => 
                           A_neg_shifted_by1_11_57_port, INPUT(263) => 
                           A_neg_shifted_by1_11_56_port, INPUT(264) => 
                           A_neg_shifted_by1_11_55_port, INPUT(265) => 
                           A_neg_shifted_by1_11_54_port, INPUT(266) => 
                           A_neg_shifted_by1_11_53_port, INPUT(267) => 
                           A_neg_shifted_by1_11_52_port, INPUT(268) => 
                           A_neg_shifted_by1_11_51_port, INPUT(269) => 
                           A_neg_shifted_by1_11_50_port, INPUT(270) => 
                           A_neg_shifted_by1_11_49_port, INPUT(271) => 
                           A_neg_shifted_by1_11_48_port, INPUT(272) => 
                           A_neg_shifted_by1_11_47_port, INPUT(273) => 
                           A_neg_shifted_by1_11_46_port, INPUT(274) => 
                           A_neg_shifted_by1_11_45_port, INPUT(275) => 
                           A_neg_shifted_by1_11_44_port, INPUT(276) => 
                           A_neg_shifted_by1_11_43_port, INPUT(277) => 
                           A_neg_shifted_by1_11_42_port, INPUT(278) => 
                           A_neg_shifted_by1_11_41_port, INPUT(279) => 
                           A_neg_shifted_by1_11_40_port, INPUT(280) => 
                           A_neg_shifted_by1_11_39_port, INPUT(281) => 
                           A_neg_shifted_by1_11_38_port, INPUT(282) => 
                           A_neg_shifted_by1_11_37_port, INPUT(283) => 
                           A_neg_shifted_by1_11_36_port, INPUT(284) => 
                           A_neg_shifted_by1_11_35_port, INPUT(285) => 
                           A_neg_shifted_by1_11_34_port, INPUT(286) => 
                           A_neg_shifted_by1_11_33_port, INPUT(287) => 
                           A_neg_shifted_by1_11_32_port, INPUT(288) => 
                           A_neg_shifted_by1_11_31_port, INPUT(289) => 
                           A_neg_shifted_by1_11_30_port, INPUT(290) => 
                           A_neg_shifted_by1_11_29_port, INPUT(291) => 
                           A_neg_shifted_by1_11_28_port, INPUT(292) => 
                           A_neg_shifted_by1_11_27_port, INPUT(293) => 
                           A_neg_shifted_by1_11_26_port, INPUT(294) => 
                           A_neg_shifted_by1_11_25_port, INPUT(295) => 
                           A_neg_shifted_by1_11_24_port, INPUT(296) => 
                           A_neg_shifted_by1_11_23_port, INPUT(297) => 
                           A_neg_shifted_by1_11_22_port, INPUT(298) => 
                           A_neg_shifted_by1_11_21_port, INPUT(299) => 
                           A_neg_shifted_by1_11_20_port, INPUT(300) => 
                           A_neg_shifted_by1_11_19_port, INPUT(301) => 
                           A_neg_shifted_by1_11_18_port, INPUT(302) => 
                           A_neg_shifted_by1_11_17_port, INPUT(303) => 
                           A_neg_shifted_by1_11_16_port, INPUT(304) => 
                           A_neg_shifted_by1_11_15_port, INPUT(305) => 
                           A_neg_shifted_by1_11_14_port, INPUT(306) => 
                           A_neg_shifted_by1_11_13_port, INPUT(307) => 
                           A_neg_shifted_by1_11_12_port, INPUT(308) => 
                           A_neg_shifted_by1_11_11_port, INPUT(309) => 
                           A_neg_shifted_by1_11_10_port, INPUT(310) => 
                           A_neg_shifted_by1_11_9_port, INPUT(311) => 
                           A_neg_shifted_by1_11_8_port, INPUT(312) => 
                           A_neg_shifted_by1_11_7_port, INPUT(313) => 
                           A_neg_shifted_by1_11_6_port, INPUT(314) => 
                           A_neg_shifted_by1_11_5_port, INPUT(315) => 
                           A_neg_shifted_by1_11_4_port, INPUT(316) => 
                           A_neg_shifted_by1_11_3_port, INPUT(317) => 
                           A_neg_shifted_by1_11_2_port, INPUT(318) => 
                           A_neg_shifted_by1_11_1_port, INPUT(319) => 
                           A_neg_shifted_by1_11_0_port, SEL(0) => 
                           selection_signal_11_2_port, SEL(1) => 
                           selection_signal_11_1_port, SEL(2) => 
                           selection_signal_11_0_port, Y(0) => 
                           OUT_MUX_11_63_port, Y(1) => OUT_MUX_11_62_port, Y(2)
                           => OUT_MUX_11_61_port, Y(3) => OUT_MUX_11_60_port, 
                           Y(4) => OUT_MUX_11_59_port, Y(5) => 
                           OUT_MUX_11_58_port, Y(6) => OUT_MUX_11_57_port, Y(7)
                           => OUT_MUX_11_56_port, Y(8) => OUT_MUX_11_55_port, 
                           Y(9) => OUT_MUX_11_54_port, Y(10) => 
                           OUT_MUX_11_53_port, Y(11) => OUT_MUX_11_52_port, 
                           Y(12) => OUT_MUX_11_51_port, Y(13) => 
                           OUT_MUX_11_50_port, Y(14) => OUT_MUX_11_49_port, 
                           Y(15) => OUT_MUX_11_48_port, Y(16) => 
                           OUT_MUX_11_47_port, Y(17) => OUT_MUX_11_46_port, 
                           Y(18) => OUT_MUX_11_45_port, Y(19) => 
                           OUT_MUX_11_44_port, Y(20) => OUT_MUX_11_43_port, 
                           Y(21) => OUT_MUX_11_42_port, Y(22) => 
                           OUT_MUX_11_41_port, Y(23) => OUT_MUX_11_40_port, 
                           Y(24) => OUT_MUX_11_39_port, Y(25) => 
                           OUT_MUX_11_38_port, Y(26) => OUT_MUX_11_37_port, 
                           Y(27) => OUT_MUX_11_36_port, Y(28) => 
                           OUT_MUX_11_35_port, Y(29) => OUT_MUX_11_34_port, 
                           Y(30) => OUT_MUX_11_33_port, Y(31) => 
                           OUT_MUX_11_32_port, Y(32) => OUT_MUX_11_31_port, 
                           Y(33) => OUT_MUX_11_30_port, Y(34) => 
                           OUT_MUX_11_29_port, Y(35) => OUT_MUX_11_28_port, 
                           Y(36) => OUT_MUX_11_27_port, Y(37) => 
                           OUT_MUX_11_26_port, Y(38) => OUT_MUX_11_25_port, 
                           Y(39) => OUT_MUX_11_24_port, Y(40) => 
                           OUT_MUX_11_23_port, Y(41) => OUT_MUX_11_22_port, 
                           Y(42) => OUT_MUX_11_21_port, Y(43) => 
                           OUT_MUX_11_20_port, Y(44) => OUT_MUX_11_19_port, 
                           Y(45) => OUT_MUX_11_18_port, Y(46) => 
                           OUT_MUX_11_17_port, Y(47) => OUT_MUX_11_16_port, 
                           Y(48) => OUT_MUX_11_15_port, Y(49) => 
                           OUT_MUX_11_14_port, Y(50) => OUT_MUX_11_13_port, 
                           Y(51) => OUT_MUX_11_12_port, Y(52) => 
                           OUT_MUX_11_11_port, Y(53) => OUT_MUX_11_10_port, 
                           Y(54) => OUT_MUX_11_9_port, Y(55) => 
                           OUT_MUX_11_8_port, Y(56) => OUT_MUX_11_7_port, Y(57)
                           => OUT_MUX_11_6_port, Y(58) => OUT_MUX_11_5_port, 
                           Y(59) => OUT_MUX_11_4_port, Y(60) => 
                           OUT_MUX_11_3_port, Y(61) => OUT_MUX_11_2_port, Y(62)
                           => OUT_MUX_11_1_port, Y(63) => OUT_MUX_11_0_port);
   MUXi_12 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_4 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_11_63_port, INPUT(65) => 
                           A_pos_shifted_by2_11_62_port, INPUT(66) => 
                           A_pos_shifted_by2_11_61_port, INPUT(67) => 
                           A_pos_shifted_by2_11_60_port, INPUT(68) => 
                           A_pos_shifted_by2_11_59_port, INPUT(69) => 
                           A_pos_shifted_by2_11_58_port, INPUT(70) => 
                           A_pos_shifted_by2_11_57_port, INPUT(71) => 
                           A_pos_shifted_by2_11_56_port, INPUT(72) => 
                           A_pos_shifted_by2_11_55_port, INPUT(73) => 
                           A_pos_shifted_by2_11_54_port, INPUT(74) => 
                           A_pos_shifted_by2_11_53_port, INPUT(75) => 
                           A_pos_shifted_by2_11_52_port, INPUT(76) => 
                           A_pos_shifted_by2_11_51_port, INPUT(77) => 
                           A_pos_shifted_by2_11_50_port, INPUT(78) => 
                           A_pos_shifted_by2_11_49_port, INPUT(79) => 
                           A_pos_shifted_by2_11_48_port, INPUT(80) => 
                           A_pos_shifted_by2_11_47_port, INPUT(81) => 
                           A_pos_shifted_by2_11_46_port, INPUT(82) => 
                           A_pos_shifted_by2_11_45_port, INPUT(83) => 
                           A_pos_shifted_by2_11_44_port, INPUT(84) => 
                           A_pos_shifted_by2_11_43_port, INPUT(85) => 
                           A_pos_shifted_by2_11_42_port, INPUT(86) => 
                           A_pos_shifted_by2_11_41_port, INPUT(87) => 
                           A_pos_shifted_by2_11_40_port, INPUT(88) => 
                           A_pos_shifted_by2_11_39_port, INPUT(89) => 
                           A_pos_shifted_by2_11_38_port, INPUT(90) => 
                           A_pos_shifted_by2_11_37_port, INPUT(91) => 
                           A_pos_shifted_by2_11_36_port, INPUT(92) => 
                           A_pos_shifted_by2_11_35_port, INPUT(93) => 
                           A_pos_shifted_by2_11_34_port, INPUT(94) => 
                           A_pos_shifted_by2_11_33_port, INPUT(95) => 
                           A_pos_shifted_by2_11_32_port, INPUT(96) => 
                           A_pos_shifted_by2_11_31_port, INPUT(97) => 
                           A_pos_shifted_by2_11_30_port, INPUT(98) => 
                           A_pos_shifted_by2_11_29_port, INPUT(99) => 
                           A_pos_shifted_by2_11_28_port, INPUT(100) => 
                           A_pos_shifted_by2_11_27_port, INPUT(101) => 
                           A_pos_shifted_by2_11_26_port, INPUT(102) => 
                           A_pos_shifted_by2_11_25_port, INPUT(103) => 
                           A_pos_shifted_by2_11_24_port, INPUT(104) => 
                           A_pos_shifted_by2_11_23_port, INPUT(105) => 
                           A_pos_shifted_by2_11_22_port, INPUT(106) => 
                           A_pos_shifted_by2_11_21_port, INPUT(107) => 
                           A_pos_shifted_by2_11_20_port, INPUT(108) => 
                           A_pos_shifted_by2_11_19_port, INPUT(109) => 
                           A_pos_shifted_by2_11_18_port, INPUT(110) => 
                           A_pos_shifted_by2_11_17_port, INPUT(111) => 
                           A_pos_shifted_by2_11_16_port, INPUT(112) => 
                           A_pos_shifted_by2_11_15_port, INPUT(113) => 
                           A_pos_shifted_by2_11_14_port, INPUT(114) => 
                           A_pos_shifted_by2_11_13_port, INPUT(115) => 
                           A_pos_shifted_by2_11_12_port, INPUT(116) => 
                           A_pos_shifted_by2_11_11_port, INPUT(117) => 
                           A_pos_shifted_by2_11_10_port, INPUT(118) => 
                           A_pos_shifted_by2_11_9_port, INPUT(119) => 
                           A_pos_shifted_by2_11_8_port, INPUT(120) => 
                           A_pos_shifted_by2_11_7_port, INPUT(121) => 
                           A_pos_shifted_by2_11_6_port, INPUT(122) => 
                           A_pos_shifted_by2_11_5_port, INPUT(123) => 
                           A_pos_shifted_by2_11_4_port, INPUT(124) => 
                           A_pos_shifted_by2_11_3_port, INPUT(125) => 
                           A_pos_shifted_by2_11_2_port, INPUT(126) => 
                           A_pos_shifted_by2_11_1_port, INPUT(127) => 
                           A_pos_shifted_by2_11_0_port, INPUT(128) => 
                           A_neg_shifted_by2_11_63_port, INPUT(129) => 
                           A_neg_shifted_by2_11_62_port, INPUT(130) => 
                           A_neg_shifted_by2_11_61_port, INPUT(131) => 
                           A_neg_shifted_by2_11_60_port, INPUT(132) => 
                           A_neg_shifted_by2_11_59_port, INPUT(133) => 
                           A_neg_shifted_by2_11_58_port, INPUT(134) => 
                           A_neg_shifted_by2_11_57_port, INPUT(135) => 
                           A_neg_shifted_by2_11_56_port, INPUT(136) => 
                           A_neg_shifted_by2_11_55_port, INPUT(137) => 
                           A_neg_shifted_by2_11_54_port, INPUT(138) => 
                           A_neg_shifted_by2_11_53_port, INPUT(139) => 
                           A_neg_shifted_by2_11_52_port, INPUT(140) => 
                           A_neg_shifted_by2_11_51_port, INPUT(141) => 
                           A_neg_shifted_by2_11_50_port, INPUT(142) => 
                           A_neg_shifted_by2_11_49_port, INPUT(143) => 
                           A_neg_shifted_by2_11_48_port, INPUT(144) => 
                           A_neg_shifted_by2_11_47_port, INPUT(145) => 
                           A_neg_shifted_by2_11_46_port, INPUT(146) => 
                           A_neg_shifted_by2_11_45_port, INPUT(147) => 
                           A_neg_shifted_by2_11_44_port, INPUT(148) => 
                           A_neg_shifted_by2_11_43_port, INPUT(149) => 
                           A_neg_shifted_by2_11_42_port, INPUT(150) => 
                           A_neg_shifted_by2_11_41_port, INPUT(151) => 
                           A_neg_shifted_by2_11_40_port, INPUT(152) => 
                           A_neg_shifted_by2_11_39_port, INPUT(153) => 
                           A_neg_shifted_by2_11_38_port, INPUT(154) => 
                           A_neg_shifted_by2_11_37_port, INPUT(155) => 
                           A_neg_shifted_by2_11_36_port, INPUT(156) => 
                           A_neg_shifted_by2_11_35_port, INPUT(157) => 
                           A_neg_shifted_by2_11_34_port, INPUT(158) => 
                           A_neg_shifted_by2_11_33_port, INPUT(159) => 
                           A_neg_shifted_by2_11_32_port, INPUT(160) => 
                           A_neg_shifted_by2_11_31_port, INPUT(161) => 
                           A_neg_shifted_by2_11_30_port, INPUT(162) => 
                           A_neg_shifted_by2_11_29_port, INPUT(163) => 
                           A_neg_shifted_by2_11_28_port, INPUT(164) => 
                           A_neg_shifted_by2_11_27_port, INPUT(165) => 
                           A_neg_shifted_by2_11_26_port, INPUT(166) => 
                           A_neg_shifted_by2_11_25_port, INPUT(167) => 
                           A_neg_shifted_by2_11_24_port, INPUT(168) => 
                           A_neg_shifted_by2_11_23_port, INPUT(169) => 
                           A_neg_shifted_by2_11_22_port, INPUT(170) => 
                           A_neg_shifted_by2_11_21_port, INPUT(171) => 
                           A_neg_shifted_by2_11_20_port, INPUT(172) => 
                           A_neg_shifted_by2_11_19_port, INPUT(173) => 
                           A_neg_shifted_by2_11_18_port, INPUT(174) => 
                           A_neg_shifted_by2_11_17_port, INPUT(175) => 
                           A_neg_shifted_by2_11_16_port, INPUT(176) => 
                           A_neg_shifted_by2_11_15_port, INPUT(177) => 
                           A_neg_shifted_by2_11_14_port, INPUT(178) => 
                           A_neg_shifted_by2_11_13_port, INPUT(179) => 
                           A_neg_shifted_by2_11_12_port, INPUT(180) => 
                           A_neg_shifted_by2_11_11_port, INPUT(181) => 
                           A_neg_shifted_by2_11_10_port, INPUT(182) => 
                           A_neg_shifted_by2_11_9_port, INPUT(183) => 
                           A_neg_shifted_by2_11_8_port, INPUT(184) => 
                           A_neg_shifted_by2_11_7_port, INPUT(185) => 
                           A_neg_shifted_by2_11_6_port, INPUT(186) => 
                           A_neg_shifted_by2_11_5_port, INPUT(187) => 
                           A_neg_shifted_by2_11_4_port, INPUT(188) => 
                           A_neg_shifted_by2_11_3_port, INPUT(189) => 
                           A_neg_shifted_by2_11_2_port, INPUT(190) => 
                           A_neg_shifted_by2_11_1_port, INPUT(191) => 
                           A_neg_shifted_by2_11_0_port, INPUT(192) => 
                           A_pos_shifted_by1_12_63_port, INPUT(193) => 
                           A_pos_shifted_by1_12_62_port, INPUT(194) => 
                           A_pos_shifted_by1_12_61_port, INPUT(195) => 
                           A_pos_shifted_by1_12_60_port, INPUT(196) => 
                           A_pos_shifted_by1_12_59_port, INPUT(197) => 
                           A_pos_shifted_by1_12_58_port, INPUT(198) => 
                           A_pos_shifted_by1_12_57_port, INPUT(199) => 
                           A_pos_shifted_by1_12_56_port, INPUT(200) => 
                           A_pos_shifted_by1_12_55_port, INPUT(201) => 
                           A_pos_shifted_by1_12_54_port, INPUT(202) => 
                           A_pos_shifted_by1_12_53_port, INPUT(203) => 
                           A_pos_shifted_by1_12_52_port, INPUT(204) => 
                           A_pos_shifted_by1_12_51_port, INPUT(205) => 
                           A_pos_shifted_by1_12_50_port, INPUT(206) => 
                           A_pos_shifted_by1_12_49_port, INPUT(207) => 
                           A_pos_shifted_by1_12_48_port, INPUT(208) => 
                           A_pos_shifted_by1_12_47_port, INPUT(209) => 
                           A_pos_shifted_by1_12_46_port, INPUT(210) => 
                           A_pos_shifted_by1_12_45_port, INPUT(211) => 
                           A_pos_shifted_by1_12_44_port, INPUT(212) => 
                           A_pos_shifted_by1_12_43_port, INPUT(213) => 
                           A_pos_shifted_by1_12_42_port, INPUT(214) => 
                           A_pos_shifted_by1_12_41_port, INPUT(215) => 
                           A_pos_shifted_by1_12_40_port, INPUT(216) => 
                           A_pos_shifted_by1_12_39_port, INPUT(217) => 
                           A_pos_shifted_by1_12_38_port, INPUT(218) => 
                           A_pos_shifted_by1_12_37_port, INPUT(219) => 
                           A_pos_shifted_by1_12_36_port, INPUT(220) => 
                           A_pos_shifted_by1_12_35_port, INPUT(221) => 
                           A_pos_shifted_by1_12_34_port, INPUT(222) => 
                           A_pos_shifted_by1_12_33_port, INPUT(223) => 
                           A_pos_shifted_by1_12_32_port, INPUT(224) => 
                           A_pos_shifted_by1_12_31_port, INPUT(225) => 
                           A_pos_shifted_by1_12_30_port, INPUT(226) => 
                           A_pos_shifted_by1_12_29_port, INPUT(227) => 
                           A_pos_shifted_by1_12_28_port, INPUT(228) => 
                           A_pos_shifted_by1_12_27_port, INPUT(229) => 
                           A_pos_shifted_by1_12_26_port, INPUT(230) => 
                           A_pos_shifted_by1_12_25_port, INPUT(231) => 
                           A_pos_shifted_by1_12_24_port, INPUT(232) => 
                           A_pos_shifted_by1_12_23_port, INPUT(233) => 
                           A_pos_shifted_by1_12_22_port, INPUT(234) => 
                           A_pos_shifted_by1_12_21_port, INPUT(235) => 
                           A_pos_shifted_by1_12_20_port, INPUT(236) => 
                           A_pos_shifted_by1_12_19_port, INPUT(237) => 
                           A_pos_shifted_by1_12_18_port, INPUT(238) => 
                           A_pos_shifted_by1_12_17_port, INPUT(239) => 
                           A_pos_shifted_by1_12_16_port, INPUT(240) => 
                           A_pos_shifted_by1_12_15_port, INPUT(241) => 
                           A_pos_shifted_by1_12_14_port, INPUT(242) => 
                           A_pos_shifted_by1_12_13_port, INPUT(243) => 
                           A_pos_shifted_by1_12_12_port, INPUT(244) => 
                           A_pos_shifted_by1_12_11_port, INPUT(245) => 
                           A_pos_shifted_by1_12_10_port, INPUT(246) => 
                           A_pos_shifted_by1_12_9_port, INPUT(247) => 
                           A_pos_shifted_by1_12_8_port, INPUT(248) => 
                           A_pos_shifted_by1_12_7_port, INPUT(249) => 
                           A_pos_shifted_by1_12_6_port, INPUT(250) => 
                           A_pos_shifted_by1_12_5_port, INPUT(251) => 
                           A_pos_shifted_by1_12_4_port, INPUT(252) => 
                           A_pos_shifted_by1_12_3_port, INPUT(253) => 
                           A_pos_shifted_by1_12_2_port, INPUT(254) => 
                           A_pos_shifted_by1_12_1_port, INPUT(255) => 
                           A_pos_shifted_by1_12_0_port, INPUT(256) => 
                           A_neg_shifted_by1_12_63_port, INPUT(257) => 
                           A_neg_shifted_by1_12_62_port, INPUT(258) => 
                           A_neg_shifted_by1_12_61_port, INPUT(259) => 
                           A_neg_shifted_by1_12_60_port, INPUT(260) => 
                           A_neg_shifted_by1_12_59_port, INPUT(261) => 
                           A_neg_shifted_by1_12_58_port, INPUT(262) => 
                           A_neg_shifted_by1_12_57_port, INPUT(263) => 
                           A_neg_shifted_by1_12_56_port, INPUT(264) => 
                           A_neg_shifted_by1_12_55_port, INPUT(265) => 
                           A_neg_shifted_by1_12_54_port, INPUT(266) => 
                           A_neg_shifted_by1_12_53_port, INPUT(267) => 
                           A_neg_shifted_by1_12_52_port, INPUT(268) => 
                           A_neg_shifted_by1_12_51_port, INPUT(269) => 
                           A_neg_shifted_by1_12_50_port, INPUT(270) => 
                           A_neg_shifted_by1_12_49_port, INPUT(271) => 
                           A_neg_shifted_by1_12_48_port, INPUT(272) => 
                           A_neg_shifted_by1_12_47_port, INPUT(273) => 
                           A_neg_shifted_by1_12_46_port, INPUT(274) => 
                           A_neg_shifted_by1_12_45_port, INPUT(275) => 
                           A_neg_shifted_by1_12_44_port, INPUT(276) => 
                           A_neg_shifted_by1_12_43_port, INPUT(277) => 
                           A_neg_shifted_by1_12_42_port, INPUT(278) => 
                           A_neg_shifted_by1_12_41_port, INPUT(279) => 
                           A_neg_shifted_by1_12_40_port, INPUT(280) => 
                           A_neg_shifted_by1_12_39_port, INPUT(281) => 
                           A_neg_shifted_by1_12_38_port, INPUT(282) => 
                           A_neg_shifted_by1_12_37_port, INPUT(283) => 
                           A_neg_shifted_by1_12_36_port, INPUT(284) => 
                           A_neg_shifted_by1_12_35_port, INPUT(285) => 
                           A_neg_shifted_by1_12_34_port, INPUT(286) => 
                           A_neg_shifted_by1_12_33_port, INPUT(287) => 
                           A_neg_shifted_by1_12_32_port, INPUT(288) => 
                           A_neg_shifted_by1_12_31_port, INPUT(289) => 
                           A_neg_shifted_by1_12_30_port, INPUT(290) => 
                           A_neg_shifted_by1_12_29_port, INPUT(291) => 
                           A_neg_shifted_by1_12_28_port, INPUT(292) => 
                           A_neg_shifted_by1_12_27_port, INPUT(293) => 
                           A_neg_shifted_by1_12_26_port, INPUT(294) => 
                           A_neg_shifted_by1_12_25_port, INPUT(295) => 
                           A_neg_shifted_by1_12_24_port, INPUT(296) => 
                           A_neg_shifted_by1_12_23_port, INPUT(297) => 
                           A_neg_shifted_by1_12_22_port, INPUT(298) => 
                           A_neg_shifted_by1_12_21_port, INPUT(299) => 
                           A_neg_shifted_by1_12_20_port, INPUT(300) => 
                           A_neg_shifted_by1_12_19_port, INPUT(301) => 
                           A_neg_shifted_by1_12_18_port, INPUT(302) => 
                           A_neg_shifted_by1_12_17_port, INPUT(303) => 
                           A_neg_shifted_by1_12_16_port, INPUT(304) => 
                           A_neg_shifted_by1_12_15_port, INPUT(305) => 
                           A_neg_shifted_by1_12_14_port, INPUT(306) => 
                           A_neg_shifted_by1_12_13_port, INPUT(307) => 
                           A_neg_shifted_by1_12_12_port, INPUT(308) => 
                           A_neg_shifted_by1_12_11_port, INPUT(309) => 
                           A_neg_shifted_by1_12_10_port, INPUT(310) => 
                           A_neg_shifted_by1_12_9_port, INPUT(311) => 
                           A_neg_shifted_by1_12_8_port, INPUT(312) => 
                           A_neg_shifted_by1_12_7_port, INPUT(313) => 
                           A_neg_shifted_by1_12_6_port, INPUT(314) => 
                           A_neg_shifted_by1_12_5_port, INPUT(315) => 
                           A_neg_shifted_by1_12_4_port, INPUT(316) => 
                           A_neg_shifted_by1_12_3_port, INPUT(317) => 
                           A_neg_shifted_by1_12_2_port, INPUT(318) => 
                           A_neg_shifted_by1_12_1_port, INPUT(319) => 
                           A_neg_shifted_by1_12_0_port, SEL(0) => 
                           selection_signal_12_2_port, SEL(1) => 
                           selection_signal_12_1_port, SEL(2) => 
                           selection_signal_12_0_port, Y(0) => 
                           OUT_MUX_12_63_port, Y(1) => OUT_MUX_12_62_port, Y(2)
                           => OUT_MUX_12_61_port, Y(3) => OUT_MUX_12_60_port, 
                           Y(4) => OUT_MUX_12_59_port, Y(5) => 
                           OUT_MUX_12_58_port, Y(6) => OUT_MUX_12_57_port, Y(7)
                           => OUT_MUX_12_56_port, Y(8) => OUT_MUX_12_55_port, 
                           Y(9) => OUT_MUX_12_54_port, Y(10) => 
                           OUT_MUX_12_53_port, Y(11) => OUT_MUX_12_52_port, 
                           Y(12) => OUT_MUX_12_51_port, Y(13) => 
                           OUT_MUX_12_50_port, Y(14) => OUT_MUX_12_49_port, 
                           Y(15) => OUT_MUX_12_48_port, Y(16) => 
                           OUT_MUX_12_47_port, Y(17) => OUT_MUX_12_46_port, 
                           Y(18) => OUT_MUX_12_45_port, Y(19) => 
                           OUT_MUX_12_44_port, Y(20) => OUT_MUX_12_43_port, 
                           Y(21) => OUT_MUX_12_42_port, Y(22) => 
                           OUT_MUX_12_41_port, Y(23) => OUT_MUX_12_40_port, 
                           Y(24) => OUT_MUX_12_39_port, Y(25) => 
                           OUT_MUX_12_38_port, Y(26) => OUT_MUX_12_37_port, 
                           Y(27) => OUT_MUX_12_36_port, Y(28) => 
                           OUT_MUX_12_35_port, Y(29) => OUT_MUX_12_34_port, 
                           Y(30) => OUT_MUX_12_33_port, Y(31) => 
                           OUT_MUX_12_32_port, Y(32) => OUT_MUX_12_31_port, 
                           Y(33) => OUT_MUX_12_30_port, Y(34) => 
                           OUT_MUX_12_29_port, Y(35) => OUT_MUX_12_28_port, 
                           Y(36) => OUT_MUX_12_27_port, Y(37) => 
                           OUT_MUX_12_26_port, Y(38) => OUT_MUX_12_25_port, 
                           Y(39) => OUT_MUX_12_24_port, Y(40) => 
                           OUT_MUX_12_23_port, Y(41) => OUT_MUX_12_22_port, 
                           Y(42) => OUT_MUX_12_21_port, Y(43) => 
                           OUT_MUX_12_20_port, Y(44) => OUT_MUX_12_19_port, 
                           Y(45) => OUT_MUX_12_18_port, Y(46) => 
                           OUT_MUX_12_17_port, Y(47) => OUT_MUX_12_16_port, 
                           Y(48) => OUT_MUX_12_15_port, Y(49) => 
                           OUT_MUX_12_14_port, Y(50) => OUT_MUX_12_13_port, 
                           Y(51) => OUT_MUX_12_12_port, Y(52) => 
                           OUT_MUX_12_11_port, Y(53) => OUT_MUX_12_10_port, 
                           Y(54) => OUT_MUX_12_9_port, Y(55) => 
                           OUT_MUX_12_8_port, Y(56) => OUT_MUX_12_7_port, Y(57)
                           => OUT_MUX_12_6_port, Y(58) => OUT_MUX_12_5_port, 
                           Y(59) => OUT_MUX_12_4_port, Y(60) => 
                           OUT_MUX_12_3_port, Y(61) => OUT_MUX_12_2_port, Y(62)
                           => OUT_MUX_12_1_port, Y(63) => OUT_MUX_12_0_port);
   MUXi_13 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_3 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_12_63_port, INPUT(65) => 
                           A_pos_shifted_by2_12_62_port, INPUT(66) => 
                           A_pos_shifted_by2_12_61_port, INPUT(67) => 
                           A_pos_shifted_by2_12_60_port, INPUT(68) => 
                           A_pos_shifted_by2_12_59_port, INPUT(69) => 
                           A_pos_shifted_by2_12_58_port, INPUT(70) => 
                           A_pos_shifted_by2_12_57_port, INPUT(71) => 
                           A_pos_shifted_by2_12_56_port, INPUT(72) => 
                           A_pos_shifted_by2_12_55_port, INPUT(73) => 
                           A_pos_shifted_by2_12_54_port, INPUT(74) => 
                           A_pos_shifted_by2_12_53_port, INPUT(75) => 
                           A_pos_shifted_by2_12_52_port, INPUT(76) => 
                           A_pos_shifted_by2_12_51_port, INPUT(77) => 
                           A_pos_shifted_by2_12_50_port, INPUT(78) => 
                           A_pos_shifted_by2_12_49_port, INPUT(79) => 
                           A_pos_shifted_by2_12_48_port, INPUT(80) => 
                           A_pos_shifted_by2_12_47_port, INPUT(81) => 
                           A_pos_shifted_by2_12_46_port, INPUT(82) => 
                           A_pos_shifted_by2_12_45_port, INPUT(83) => 
                           A_pos_shifted_by2_12_44_port, INPUT(84) => 
                           A_pos_shifted_by2_12_43_port, INPUT(85) => 
                           A_pos_shifted_by2_12_42_port, INPUT(86) => 
                           A_pos_shifted_by2_12_41_port, INPUT(87) => 
                           A_pos_shifted_by2_12_40_port, INPUT(88) => 
                           A_pos_shifted_by2_12_39_port, INPUT(89) => 
                           A_pos_shifted_by2_12_38_port, INPUT(90) => 
                           A_pos_shifted_by2_12_37_port, INPUT(91) => 
                           A_pos_shifted_by2_12_36_port, INPUT(92) => 
                           A_pos_shifted_by2_12_35_port, INPUT(93) => 
                           A_pos_shifted_by2_12_34_port, INPUT(94) => 
                           A_pos_shifted_by2_12_33_port, INPUT(95) => 
                           A_pos_shifted_by2_12_32_port, INPUT(96) => 
                           A_pos_shifted_by2_12_31_port, INPUT(97) => 
                           A_pos_shifted_by2_12_30_port, INPUT(98) => 
                           A_pos_shifted_by2_12_29_port, INPUT(99) => 
                           A_pos_shifted_by2_12_28_port, INPUT(100) => 
                           A_pos_shifted_by2_12_27_port, INPUT(101) => 
                           A_pos_shifted_by2_12_26_port, INPUT(102) => 
                           A_pos_shifted_by2_12_25_port, INPUT(103) => 
                           A_pos_shifted_by2_12_24_port, INPUT(104) => 
                           A_pos_shifted_by2_12_23_port, INPUT(105) => 
                           A_pos_shifted_by2_12_22_port, INPUT(106) => 
                           A_pos_shifted_by2_12_21_port, INPUT(107) => 
                           A_pos_shifted_by2_12_20_port, INPUT(108) => 
                           A_pos_shifted_by2_12_19_port, INPUT(109) => 
                           A_pos_shifted_by2_12_18_port, INPUT(110) => 
                           A_pos_shifted_by2_12_17_port, INPUT(111) => 
                           A_pos_shifted_by2_12_16_port, INPUT(112) => 
                           A_pos_shifted_by2_12_15_port, INPUT(113) => 
                           A_pos_shifted_by2_12_14_port, INPUT(114) => 
                           A_pos_shifted_by2_12_13_port, INPUT(115) => 
                           A_pos_shifted_by2_12_12_port, INPUT(116) => 
                           A_pos_shifted_by2_12_11_port, INPUT(117) => 
                           A_pos_shifted_by2_12_10_port, INPUT(118) => 
                           A_pos_shifted_by2_12_9_port, INPUT(119) => 
                           A_pos_shifted_by2_12_8_port, INPUT(120) => 
                           A_pos_shifted_by2_12_7_port, INPUT(121) => 
                           A_pos_shifted_by2_12_6_port, INPUT(122) => 
                           A_pos_shifted_by2_12_5_port, INPUT(123) => 
                           A_pos_shifted_by2_12_4_port, INPUT(124) => 
                           A_pos_shifted_by2_12_3_port, INPUT(125) => 
                           A_pos_shifted_by2_12_2_port, INPUT(126) => 
                           A_pos_shifted_by2_12_1_port, INPUT(127) => 
                           A_pos_shifted_by2_12_0_port, INPUT(128) => 
                           A_neg_shifted_by2_12_63_port, INPUT(129) => 
                           A_neg_shifted_by2_12_62_port, INPUT(130) => 
                           A_neg_shifted_by2_12_61_port, INPUT(131) => 
                           A_neg_shifted_by2_12_60_port, INPUT(132) => 
                           A_neg_shifted_by2_12_59_port, INPUT(133) => 
                           A_neg_shifted_by2_12_58_port, INPUT(134) => 
                           A_neg_shifted_by2_12_57_port, INPUT(135) => 
                           A_neg_shifted_by2_12_56_port, INPUT(136) => 
                           A_neg_shifted_by2_12_55_port, INPUT(137) => 
                           A_neg_shifted_by2_12_54_port, INPUT(138) => 
                           A_neg_shifted_by2_12_53_port, INPUT(139) => 
                           A_neg_shifted_by2_12_52_port, INPUT(140) => 
                           A_neg_shifted_by2_12_51_port, INPUT(141) => 
                           A_neg_shifted_by2_12_50_port, INPUT(142) => 
                           A_neg_shifted_by2_12_49_port, INPUT(143) => 
                           A_neg_shifted_by2_12_48_port, INPUT(144) => 
                           A_neg_shifted_by2_12_47_port, INPUT(145) => 
                           A_neg_shifted_by2_12_46_port, INPUT(146) => 
                           A_neg_shifted_by2_12_45_port, INPUT(147) => 
                           A_neg_shifted_by2_12_44_port, INPUT(148) => 
                           A_neg_shifted_by2_12_43_port, INPUT(149) => 
                           A_neg_shifted_by2_12_42_port, INPUT(150) => 
                           A_neg_shifted_by2_12_41_port, INPUT(151) => 
                           A_neg_shifted_by2_12_40_port, INPUT(152) => 
                           A_neg_shifted_by2_12_39_port, INPUT(153) => 
                           A_neg_shifted_by2_12_38_port, INPUT(154) => 
                           A_neg_shifted_by2_12_37_port, INPUT(155) => 
                           A_neg_shifted_by2_12_36_port, INPUT(156) => 
                           A_neg_shifted_by2_12_35_port, INPUT(157) => 
                           A_neg_shifted_by2_12_34_port, INPUT(158) => 
                           A_neg_shifted_by2_12_33_port, INPUT(159) => 
                           A_neg_shifted_by2_12_32_port, INPUT(160) => 
                           A_neg_shifted_by2_12_31_port, INPUT(161) => 
                           A_neg_shifted_by2_12_30_port, INPUT(162) => 
                           A_neg_shifted_by2_12_29_port, INPUT(163) => 
                           A_neg_shifted_by2_12_28_port, INPUT(164) => 
                           A_neg_shifted_by2_12_27_port, INPUT(165) => 
                           A_neg_shifted_by2_12_26_port, INPUT(166) => 
                           A_neg_shifted_by2_12_25_port, INPUT(167) => 
                           A_neg_shifted_by2_12_24_port, INPUT(168) => 
                           A_neg_shifted_by2_12_23_port, INPUT(169) => 
                           A_neg_shifted_by2_12_22_port, INPUT(170) => 
                           A_neg_shifted_by2_12_21_port, INPUT(171) => 
                           A_neg_shifted_by2_12_20_port, INPUT(172) => 
                           A_neg_shifted_by2_12_19_port, INPUT(173) => 
                           A_neg_shifted_by2_12_18_port, INPUT(174) => 
                           A_neg_shifted_by2_12_17_port, INPUT(175) => 
                           A_neg_shifted_by2_12_16_port, INPUT(176) => 
                           A_neg_shifted_by2_12_15_port, INPUT(177) => 
                           A_neg_shifted_by2_12_14_port, INPUT(178) => 
                           A_neg_shifted_by2_12_13_port, INPUT(179) => 
                           A_neg_shifted_by2_12_12_port, INPUT(180) => 
                           A_neg_shifted_by2_12_11_port, INPUT(181) => 
                           A_neg_shifted_by2_12_10_port, INPUT(182) => 
                           A_neg_shifted_by2_12_9_port, INPUT(183) => 
                           A_neg_shifted_by2_12_8_port, INPUT(184) => 
                           A_neg_shifted_by2_12_7_port, INPUT(185) => 
                           A_neg_shifted_by2_12_6_port, INPUT(186) => 
                           A_neg_shifted_by2_12_5_port, INPUT(187) => 
                           A_neg_shifted_by2_12_4_port, INPUT(188) => 
                           A_neg_shifted_by2_12_3_port, INPUT(189) => 
                           A_neg_shifted_by2_12_2_port, INPUT(190) => 
                           A_neg_shifted_by2_12_1_port, INPUT(191) => 
                           A_neg_shifted_by2_12_0_port, INPUT(192) => 
                           A_pos_shifted_by1_13_63_port, INPUT(193) => 
                           A_pos_shifted_by1_13_62_port, INPUT(194) => 
                           A_pos_shifted_by1_13_61_port, INPUT(195) => 
                           A_pos_shifted_by1_13_60_port, INPUT(196) => 
                           A_pos_shifted_by1_13_59_port, INPUT(197) => 
                           A_pos_shifted_by1_13_58_port, INPUT(198) => 
                           A_pos_shifted_by1_13_57_port, INPUT(199) => 
                           A_pos_shifted_by1_13_56_port, INPUT(200) => 
                           A_pos_shifted_by1_13_55_port, INPUT(201) => 
                           A_pos_shifted_by1_13_54_port, INPUT(202) => 
                           A_pos_shifted_by1_13_53_port, INPUT(203) => 
                           A_pos_shifted_by1_13_52_port, INPUT(204) => 
                           A_pos_shifted_by1_13_51_port, INPUT(205) => 
                           A_pos_shifted_by1_13_50_port, INPUT(206) => 
                           A_pos_shifted_by1_13_49_port, INPUT(207) => 
                           A_pos_shifted_by1_13_48_port, INPUT(208) => 
                           A_pos_shifted_by1_13_47_port, INPUT(209) => 
                           A_pos_shifted_by1_13_46_port, INPUT(210) => 
                           A_pos_shifted_by1_13_45_port, INPUT(211) => 
                           A_pos_shifted_by1_13_44_port, INPUT(212) => 
                           A_pos_shifted_by1_13_43_port, INPUT(213) => 
                           A_pos_shifted_by1_13_42_port, INPUT(214) => 
                           A_pos_shifted_by1_13_41_port, INPUT(215) => 
                           A_pos_shifted_by1_13_40_port, INPUT(216) => 
                           A_pos_shifted_by1_13_39_port, INPUT(217) => 
                           A_pos_shifted_by1_13_38_port, INPUT(218) => 
                           A_pos_shifted_by1_13_37_port, INPUT(219) => 
                           A_pos_shifted_by1_13_36_port, INPUT(220) => 
                           A_pos_shifted_by1_13_35_port, INPUT(221) => 
                           A_pos_shifted_by1_13_34_port, INPUT(222) => 
                           A_pos_shifted_by1_13_33_port, INPUT(223) => 
                           A_pos_shifted_by1_13_32_port, INPUT(224) => 
                           A_pos_shifted_by1_13_31_port, INPUT(225) => 
                           A_pos_shifted_by1_13_30_port, INPUT(226) => 
                           A_pos_shifted_by1_13_29_port, INPUT(227) => 
                           A_pos_shifted_by1_13_28_port, INPUT(228) => 
                           A_pos_shifted_by1_13_27_port, INPUT(229) => 
                           A_pos_shifted_by1_13_26_port, INPUT(230) => 
                           A_pos_shifted_by1_13_25_port, INPUT(231) => 
                           A_pos_shifted_by1_13_24_port, INPUT(232) => 
                           A_pos_shifted_by1_13_23_port, INPUT(233) => 
                           A_pos_shifted_by1_13_22_port, INPUT(234) => 
                           A_pos_shifted_by1_13_21_port, INPUT(235) => 
                           A_pos_shifted_by1_13_20_port, INPUT(236) => 
                           A_pos_shifted_by1_13_19_port, INPUT(237) => 
                           A_pos_shifted_by1_13_18_port, INPUT(238) => 
                           A_pos_shifted_by1_13_17_port, INPUT(239) => 
                           A_pos_shifted_by1_13_16_port, INPUT(240) => 
                           A_pos_shifted_by1_13_15_port, INPUT(241) => 
                           A_pos_shifted_by1_13_14_port, INPUT(242) => 
                           A_pos_shifted_by1_13_13_port, INPUT(243) => 
                           A_pos_shifted_by1_13_12_port, INPUT(244) => 
                           A_pos_shifted_by1_13_11_port, INPUT(245) => 
                           A_pos_shifted_by1_13_10_port, INPUT(246) => 
                           A_pos_shifted_by1_13_9_port, INPUT(247) => 
                           A_pos_shifted_by1_13_8_port, INPUT(248) => 
                           A_pos_shifted_by1_13_7_port, INPUT(249) => 
                           A_pos_shifted_by1_13_6_port, INPUT(250) => 
                           A_pos_shifted_by1_13_5_port, INPUT(251) => 
                           A_pos_shifted_by1_13_4_port, INPUT(252) => 
                           A_pos_shifted_by1_13_3_port, INPUT(253) => 
                           A_pos_shifted_by1_13_2_port, INPUT(254) => 
                           A_pos_shifted_by1_13_1_port, INPUT(255) => 
                           A_pos_shifted_by1_13_0_port, INPUT(256) => 
                           A_neg_shifted_by1_13_63_port, INPUT(257) => 
                           A_neg_shifted_by1_13_62_port, INPUT(258) => 
                           A_neg_shifted_by1_13_61_port, INPUT(259) => 
                           A_neg_shifted_by1_13_60_port, INPUT(260) => 
                           A_neg_shifted_by1_13_59_port, INPUT(261) => 
                           A_neg_shifted_by1_13_58_port, INPUT(262) => 
                           A_neg_shifted_by1_13_57_port, INPUT(263) => 
                           A_neg_shifted_by1_13_56_port, INPUT(264) => 
                           A_neg_shifted_by1_13_55_port, INPUT(265) => 
                           A_neg_shifted_by1_13_54_port, INPUT(266) => 
                           A_neg_shifted_by1_13_53_port, INPUT(267) => 
                           A_neg_shifted_by1_13_52_port, INPUT(268) => 
                           A_neg_shifted_by1_13_51_port, INPUT(269) => 
                           A_neg_shifted_by1_13_50_port, INPUT(270) => 
                           A_neg_shifted_by1_13_49_port, INPUT(271) => 
                           A_neg_shifted_by1_13_48_port, INPUT(272) => 
                           A_neg_shifted_by1_13_47_port, INPUT(273) => 
                           A_neg_shifted_by1_13_46_port, INPUT(274) => 
                           A_neg_shifted_by1_13_45_port, INPUT(275) => 
                           A_neg_shifted_by1_13_44_port, INPUT(276) => 
                           A_neg_shifted_by1_13_43_port, INPUT(277) => 
                           A_neg_shifted_by1_13_42_port, INPUT(278) => 
                           A_neg_shifted_by1_13_41_port, INPUT(279) => 
                           A_neg_shifted_by1_13_40_port, INPUT(280) => 
                           A_neg_shifted_by1_13_39_port, INPUT(281) => 
                           A_neg_shifted_by1_13_38_port, INPUT(282) => 
                           A_neg_shifted_by1_13_37_port, INPUT(283) => 
                           A_neg_shifted_by1_13_36_port, INPUT(284) => 
                           A_neg_shifted_by1_13_35_port, INPUT(285) => 
                           A_neg_shifted_by1_13_34_port, INPUT(286) => 
                           A_neg_shifted_by1_13_33_port, INPUT(287) => 
                           A_neg_shifted_by1_13_32_port, INPUT(288) => 
                           A_neg_shifted_by1_13_31_port, INPUT(289) => 
                           A_neg_shifted_by1_13_30_port, INPUT(290) => 
                           A_neg_shifted_by1_13_29_port, INPUT(291) => 
                           A_neg_shifted_by1_13_28_port, INPUT(292) => 
                           A_neg_shifted_by1_13_27_port, INPUT(293) => 
                           A_neg_shifted_by1_13_26_port, INPUT(294) => 
                           A_neg_shifted_by1_13_25_port, INPUT(295) => 
                           A_neg_shifted_by1_13_24_port, INPUT(296) => 
                           A_neg_shifted_by1_13_23_port, INPUT(297) => 
                           A_neg_shifted_by1_13_22_port, INPUT(298) => 
                           A_neg_shifted_by1_13_21_port, INPUT(299) => 
                           A_neg_shifted_by1_13_20_port, INPUT(300) => 
                           A_neg_shifted_by1_13_19_port, INPUT(301) => 
                           A_neg_shifted_by1_13_18_port, INPUT(302) => 
                           A_neg_shifted_by1_13_17_port, INPUT(303) => 
                           A_neg_shifted_by1_13_16_port, INPUT(304) => 
                           A_neg_shifted_by1_13_15_port, INPUT(305) => 
                           A_neg_shifted_by1_13_14_port, INPUT(306) => 
                           A_neg_shifted_by1_13_13_port, INPUT(307) => 
                           A_neg_shifted_by1_13_12_port, INPUT(308) => 
                           A_neg_shifted_by1_13_11_port, INPUT(309) => 
                           A_neg_shifted_by1_13_10_port, INPUT(310) => 
                           A_neg_shifted_by1_13_9_port, INPUT(311) => 
                           A_neg_shifted_by1_13_8_port, INPUT(312) => 
                           A_neg_shifted_by1_13_7_port, INPUT(313) => 
                           A_neg_shifted_by1_13_6_port, INPUT(314) => 
                           A_neg_shifted_by1_13_5_port, INPUT(315) => 
                           A_neg_shifted_by1_13_4_port, INPUT(316) => 
                           A_neg_shifted_by1_13_3_port, INPUT(317) => 
                           A_neg_shifted_by1_13_2_port, INPUT(318) => 
                           A_neg_shifted_by1_13_1_port, INPUT(319) => 
                           A_neg_shifted_by1_13_0_port, SEL(0) => 
                           selection_signal_13_2_port, SEL(1) => 
                           selection_signal_13_1_port, SEL(2) => 
                           selection_signal_13_0_port, Y(0) => 
                           OUT_MUX_13_63_port, Y(1) => OUT_MUX_13_62_port, Y(2)
                           => OUT_MUX_13_61_port, Y(3) => OUT_MUX_13_60_port, 
                           Y(4) => OUT_MUX_13_59_port, Y(5) => 
                           OUT_MUX_13_58_port, Y(6) => OUT_MUX_13_57_port, Y(7)
                           => OUT_MUX_13_56_port, Y(8) => OUT_MUX_13_55_port, 
                           Y(9) => OUT_MUX_13_54_port, Y(10) => 
                           OUT_MUX_13_53_port, Y(11) => OUT_MUX_13_52_port, 
                           Y(12) => OUT_MUX_13_51_port, Y(13) => 
                           OUT_MUX_13_50_port, Y(14) => OUT_MUX_13_49_port, 
                           Y(15) => OUT_MUX_13_48_port, Y(16) => 
                           OUT_MUX_13_47_port, Y(17) => OUT_MUX_13_46_port, 
                           Y(18) => OUT_MUX_13_45_port, Y(19) => 
                           OUT_MUX_13_44_port, Y(20) => OUT_MUX_13_43_port, 
                           Y(21) => OUT_MUX_13_42_port, Y(22) => 
                           OUT_MUX_13_41_port, Y(23) => OUT_MUX_13_40_port, 
                           Y(24) => OUT_MUX_13_39_port, Y(25) => 
                           OUT_MUX_13_38_port, Y(26) => OUT_MUX_13_37_port, 
                           Y(27) => OUT_MUX_13_36_port, Y(28) => 
                           OUT_MUX_13_35_port, Y(29) => OUT_MUX_13_34_port, 
                           Y(30) => OUT_MUX_13_33_port, Y(31) => 
                           OUT_MUX_13_32_port, Y(32) => OUT_MUX_13_31_port, 
                           Y(33) => OUT_MUX_13_30_port, Y(34) => 
                           OUT_MUX_13_29_port, Y(35) => OUT_MUX_13_28_port, 
                           Y(36) => OUT_MUX_13_27_port, Y(37) => 
                           OUT_MUX_13_26_port, Y(38) => OUT_MUX_13_25_port, 
                           Y(39) => OUT_MUX_13_24_port, Y(40) => 
                           OUT_MUX_13_23_port, Y(41) => OUT_MUX_13_22_port, 
                           Y(42) => OUT_MUX_13_21_port, Y(43) => 
                           OUT_MUX_13_20_port, Y(44) => OUT_MUX_13_19_port, 
                           Y(45) => OUT_MUX_13_18_port, Y(46) => 
                           OUT_MUX_13_17_port, Y(47) => OUT_MUX_13_16_port, 
                           Y(48) => OUT_MUX_13_15_port, Y(49) => 
                           OUT_MUX_13_14_port, Y(50) => OUT_MUX_13_13_port, 
                           Y(51) => OUT_MUX_13_12_port, Y(52) => 
                           OUT_MUX_13_11_port, Y(53) => OUT_MUX_13_10_port, 
                           Y(54) => OUT_MUX_13_9_port, Y(55) => 
                           OUT_MUX_13_8_port, Y(56) => OUT_MUX_13_7_port, Y(57)
                           => OUT_MUX_13_6_port, Y(58) => OUT_MUX_13_5_port, 
                           Y(59) => OUT_MUX_13_4_port, Y(60) => 
                           OUT_MUX_13_3_port, Y(61) => OUT_MUX_13_2_port, Y(62)
                           => OUT_MUX_13_1_port, Y(63) => OUT_MUX_13_0_port);
   MUXi_14 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_2 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_13_63_port, INPUT(65) => 
                           A_pos_shifted_by2_13_62_port, INPUT(66) => 
                           A_pos_shifted_by2_13_61_port, INPUT(67) => 
                           A_pos_shifted_by2_13_60_port, INPUT(68) => 
                           A_pos_shifted_by2_13_59_port, INPUT(69) => 
                           A_pos_shifted_by2_13_58_port, INPUT(70) => 
                           A_pos_shifted_by2_13_57_port, INPUT(71) => 
                           A_pos_shifted_by2_13_56_port, INPUT(72) => 
                           A_pos_shifted_by2_13_55_port, INPUT(73) => 
                           A_pos_shifted_by2_13_54_port, INPUT(74) => 
                           A_pos_shifted_by2_13_53_port, INPUT(75) => 
                           A_pos_shifted_by2_13_52_port, INPUT(76) => 
                           A_pos_shifted_by2_13_51_port, INPUT(77) => 
                           A_pos_shifted_by2_13_50_port, INPUT(78) => 
                           A_pos_shifted_by2_13_49_port, INPUT(79) => 
                           A_pos_shifted_by2_13_48_port, INPUT(80) => 
                           A_pos_shifted_by2_13_47_port, INPUT(81) => 
                           A_pos_shifted_by2_13_46_port, INPUT(82) => 
                           A_pos_shifted_by2_13_45_port, INPUT(83) => 
                           A_pos_shifted_by2_13_44_port, INPUT(84) => 
                           A_pos_shifted_by2_13_43_port, INPUT(85) => 
                           A_pos_shifted_by2_13_42_port, INPUT(86) => 
                           A_pos_shifted_by2_13_41_port, INPUT(87) => 
                           A_pos_shifted_by2_13_40_port, INPUT(88) => 
                           A_pos_shifted_by2_13_39_port, INPUT(89) => 
                           A_pos_shifted_by2_13_38_port, INPUT(90) => 
                           A_pos_shifted_by2_13_37_port, INPUT(91) => 
                           A_pos_shifted_by2_13_36_port, INPUT(92) => 
                           A_pos_shifted_by2_13_35_port, INPUT(93) => 
                           A_pos_shifted_by2_13_34_port, INPUT(94) => 
                           A_pos_shifted_by2_13_33_port, INPUT(95) => 
                           A_pos_shifted_by2_13_32_port, INPUT(96) => 
                           A_pos_shifted_by2_13_31_port, INPUT(97) => 
                           A_pos_shifted_by2_13_30_port, INPUT(98) => 
                           A_pos_shifted_by2_13_29_port, INPUT(99) => 
                           A_pos_shifted_by2_13_28_port, INPUT(100) => 
                           A_pos_shifted_by2_13_27_port, INPUT(101) => 
                           A_pos_shifted_by2_13_26_port, INPUT(102) => 
                           A_pos_shifted_by2_13_25_port, INPUT(103) => 
                           A_pos_shifted_by2_13_24_port, INPUT(104) => 
                           A_pos_shifted_by2_13_23_port, INPUT(105) => 
                           A_pos_shifted_by2_13_22_port, INPUT(106) => 
                           A_pos_shifted_by2_13_21_port, INPUT(107) => 
                           A_pos_shifted_by2_13_20_port, INPUT(108) => 
                           A_pos_shifted_by2_13_19_port, INPUT(109) => 
                           A_pos_shifted_by2_13_18_port, INPUT(110) => 
                           A_pos_shifted_by2_13_17_port, INPUT(111) => 
                           A_pos_shifted_by2_13_16_port, INPUT(112) => 
                           A_pos_shifted_by2_13_15_port, INPUT(113) => 
                           A_pos_shifted_by2_13_14_port, INPUT(114) => 
                           A_pos_shifted_by2_13_13_port, INPUT(115) => 
                           A_pos_shifted_by2_13_12_port, INPUT(116) => 
                           A_pos_shifted_by2_13_11_port, INPUT(117) => 
                           A_pos_shifted_by2_13_10_port, INPUT(118) => 
                           A_pos_shifted_by2_13_9_port, INPUT(119) => 
                           A_pos_shifted_by2_13_8_port, INPUT(120) => 
                           A_pos_shifted_by2_13_7_port, INPUT(121) => 
                           A_pos_shifted_by2_13_6_port, INPUT(122) => 
                           A_pos_shifted_by2_13_5_port, INPUT(123) => 
                           A_pos_shifted_by2_13_4_port, INPUT(124) => 
                           A_pos_shifted_by2_13_3_port, INPUT(125) => 
                           A_pos_shifted_by2_13_2_port, INPUT(126) => 
                           A_pos_shifted_by2_13_1_port, INPUT(127) => 
                           A_pos_shifted_by2_13_0_port, INPUT(128) => 
                           A_neg_shifted_by2_13_63_port, INPUT(129) => 
                           A_neg_shifted_by2_13_62_port, INPUT(130) => 
                           A_neg_shifted_by2_13_61_port, INPUT(131) => 
                           A_neg_shifted_by2_13_60_port, INPUT(132) => 
                           A_neg_shifted_by2_13_59_port, INPUT(133) => 
                           A_neg_shifted_by2_13_58_port, INPUT(134) => 
                           A_neg_shifted_by2_13_57_port, INPUT(135) => 
                           A_neg_shifted_by2_13_56_port, INPUT(136) => 
                           A_neg_shifted_by2_13_55_port, INPUT(137) => 
                           A_neg_shifted_by2_13_54_port, INPUT(138) => 
                           A_neg_shifted_by2_13_53_port, INPUT(139) => 
                           A_neg_shifted_by2_13_52_port, INPUT(140) => 
                           A_neg_shifted_by2_13_51_port, INPUT(141) => 
                           A_neg_shifted_by2_13_50_port, INPUT(142) => 
                           A_neg_shifted_by2_13_49_port, INPUT(143) => 
                           A_neg_shifted_by2_13_48_port, INPUT(144) => 
                           A_neg_shifted_by2_13_47_port, INPUT(145) => 
                           A_neg_shifted_by2_13_46_port, INPUT(146) => 
                           A_neg_shifted_by2_13_45_port, INPUT(147) => 
                           A_neg_shifted_by2_13_44_port, INPUT(148) => 
                           A_neg_shifted_by2_13_43_port, INPUT(149) => 
                           A_neg_shifted_by2_13_42_port, INPUT(150) => 
                           A_neg_shifted_by2_13_41_port, INPUT(151) => 
                           A_neg_shifted_by2_13_40_port, INPUT(152) => 
                           A_neg_shifted_by2_13_39_port, INPUT(153) => 
                           A_neg_shifted_by2_13_38_port, INPUT(154) => 
                           A_neg_shifted_by2_13_37_port, INPUT(155) => 
                           A_neg_shifted_by2_13_36_port, INPUT(156) => 
                           A_neg_shifted_by2_13_35_port, INPUT(157) => 
                           A_neg_shifted_by2_13_34_port, INPUT(158) => 
                           A_neg_shifted_by2_13_33_port, INPUT(159) => 
                           A_neg_shifted_by2_13_32_port, INPUT(160) => 
                           A_neg_shifted_by2_13_31_port, INPUT(161) => 
                           A_neg_shifted_by2_13_30_port, INPUT(162) => 
                           A_neg_shifted_by2_13_29_port, INPUT(163) => 
                           A_neg_shifted_by2_13_28_port, INPUT(164) => 
                           A_neg_shifted_by2_13_27_port, INPUT(165) => 
                           A_neg_shifted_by2_13_26_port, INPUT(166) => 
                           A_neg_shifted_by2_13_25_port, INPUT(167) => 
                           A_neg_shifted_by2_13_24_port, INPUT(168) => 
                           A_neg_shifted_by2_13_23_port, INPUT(169) => 
                           A_neg_shifted_by2_13_22_port, INPUT(170) => 
                           A_neg_shifted_by2_13_21_port, INPUT(171) => 
                           A_neg_shifted_by2_13_20_port, INPUT(172) => 
                           A_neg_shifted_by2_13_19_port, INPUT(173) => 
                           A_neg_shifted_by2_13_18_port, INPUT(174) => 
                           A_neg_shifted_by2_13_17_port, INPUT(175) => 
                           A_neg_shifted_by2_13_16_port, INPUT(176) => 
                           A_neg_shifted_by2_13_15_port, INPUT(177) => 
                           A_neg_shifted_by2_13_14_port, INPUT(178) => 
                           A_neg_shifted_by2_13_13_port, INPUT(179) => 
                           A_neg_shifted_by2_13_12_port, INPUT(180) => 
                           A_neg_shifted_by2_13_11_port, INPUT(181) => 
                           A_neg_shifted_by2_13_10_port, INPUT(182) => 
                           A_neg_shifted_by2_13_9_port, INPUT(183) => 
                           A_neg_shifted_by2_13_8_port, INPUT(184) => 
                           A_neg_shifted_by2_13_7_port, INPUT(185) => 
                           A_neg_shifted_by2_13_6_port, INPUT(186) => 
                           A_neg_shifted_by2_13_5_port, INPUT(187) => 
                           A_neg_shifted_by2_13_4_port, INPUT(188) => 
                           A_neg_shifted_by2_13_3_port, INPUT(189) => 
                           A_neg_shifted_by2_13_2_port, INPUT(190) => 
                           A_neg_shifted_by2_13_1_port, INPUT(191) => 
                           A_neg_shifted_by2_13_0_port, INPUT(192) => 
                           A_pos_shifted_by1_14_63_port, INPUT(193) => 
                           A_pos_shifted_by1_14_62_port, INPUT(194) => 
                           A_pos_shifted_by1_14_61_port, INPUT(195) => 
                           A_pos_shifted_by1_14_60_port, INPUT(196) => 
                           A_pos_shifted_by1_14_59_port, INPUT(197) => 
                           A_pos_shifted_by1_14_58_port, INPUT(198) => 
                           A_pos_shifted_by1_14_57_port, INPUT(199) => 
                           A_pos_shifted_by1_14_56_port, INPUT(200) => 
                           A_pos_shifted_by1_14_55_port, INPUT(201) => 
                           A_pos_shifted_by1_14_54_port, INPUT(202) => 
                           A_pos_shifted_by1_14_53_port, INPUT(203) => 
                           A_pos_shifted_by1_14_52_port, INPUT(204) => 
                           A_pos_shifted_by1_14_51_port, INPUT(205) => 
                           A_pos_shifted_by1_14_50_port, INPUT(206) => 
                           A_pos_shifted_by1_14_49_port, INPUT(207) => 
                           A_pos_shifted_by1_14_48_port, INPUT(208) => 
                           A_pos_shifted_by1_14_47_port, INPUT(209) => 
                           A_pos_shifted_by1_14_46_port, INPUT(210) => 
                           A_pos_shifted_by1_14_45_port, INPUT(211) => 
                           A_pos_shifted_by1_14_44_port, INPUT(212) => 
                           A_pos_shifted_by1_14_43_port, INPUT(213) => 
                           A_pos_shifted_by1_14_42_port, INPUT(214) => 
                           A_pos_shifted_by1_14_41_port, INPUT(215) => 
                           A_pos_shifted_by1_14_40_port, INPUT(216) => 
                           A_pos_shifted_by1_14_39_port, INPUT(217) => 
                           A_pos_shifted_by1_14_38_port, INPUT(218) => 
                           A_pos_shifted_by1_14_37_port, INPUT(219) => 
                           A_pos_shifted_by1_14_36_port, INPUT(220) => 
                           A_pos_shifted_by1_14_35_port, INPUT(221) => 
                           A_pos_shifted_by1_14_34_port, INPUT(222) => 
                           A_pos_shifted_by1_14_33_port, INPUT(223) => 
                           A_pos_shifted_by1_14_32_port, INPUT(224) => 
                           A_pos_shifted_by1_14_31_port, INPUT(225) => 
                           A_pos_shifted_by1_14_30_port, INPUT(226) => 
                           A_pos_shifted_by1_14_29_port, INPUT(227) => 
                           A_pos_shifted_by1_14_28_port, INPUT(228) => 
                           A_pos_shifted_by1_14_27_port, INPUT(229) => 
                           A_pos_shifted_by1_14_26_port, INPUT(230) => 
                           A_pos_shifted_by1_14_25_port, INPUT(231) => 
                           A_pos_shifted_by1_14_24_port, INPUT(232) => 
                           A_pos_shifted_by1_14_23_port, INPUT(233) => 
                           A_pos_shifted_by1_14_22_port, INPUT(234) => 
                           A_pos_shifted_by1_14_21_port, INPUT(235) => 
                           A_pos_shifted_by1_14_20_port, INPUT(236) => 
                           A_pos_shifted_by1_14_19_port, INPUT(237) => 
                           A_pos_shifted_by1_14_18_port, INPUT(238) => 
                           A_pos_shifted_by1_14_17_port, INPUT(239) => 
                           A_pos_shifted_by1_14_16_port, INPUT(240) => 
                           A_pos_shifted_by1_14_15_port, INPUT(241) => 
                           A_pos_shifted_by1_14_14_port, INPUT(242) => 
                           A_pos_shifted_by1_14_13_port, INPUT(243) => 
                           A_pos_shifted_by1_14_12_port, INPUT(244) => 
                           A_pos_shifted_by1_14_11_port, INPUT(245) => 
                           A_pos_shifted_by1_14_10_port, INPUT(246) => 
                           A_pos_shifted_by1_14_9_port, INPUT(247) => 
                           A_pos_shifted_by1_14_8_port, INPUT(248) => 
                           A_pos_shifted_by1_14_7_port, INPUT(249) => 
                           A_pos_shifted_by1_14_6_port, INPUT(250) => 
                           A_pos_shifted_by1_14_5_port, INPUT(251) => 
                           A_pos_shifted_by1_14_4_port, INPUT(252) => 
                           A_pos_shifted_by1_14_3_port, INPUT(253) => 
                           A_pos_shifted_by1_14_2_port, INPUT(254) => 
                           A_pos_shifted_by1_14_1_port, INPUT(255) => 
                           A_pos_shifted_by1_14_0_port, INPUT(256) => 
                           A_neg_shifted_by1_14_63_port, INPUT(257) => 
                           A_neg_shifted_by1_14_62_port, INPUT(258) => 
                           A_neg_shifted_by1_14_61_port, INPUT(259) => 
                           A_neg_shifted_by1_14_60_port, INPUT(260) => 
                           A_neg_shifted_by1_14_59_port, INPUT(261) => 
                           A_neg_shifted_by1_14_58_port, INPUT(262) => 
                           A_neg_shifted_by1_14_57_port, INPUT(263) => 
                           A_neg_shifted_by1_14_56_port, INPUT(264) => 
                           A_neg_shifted_by1_14_55_port, INPUT(265) => 
                           A_neg_shifted_by1_14_54_port, INPUT(266) => 
                           A_neg_shifted_by1_14_53_port, INPUT(267) => 
                           A_neg_shifted_by1_14_52_port, INPUT(268) => 
                           A_neg_shifted_by1_14_51_port, INPUT(269) => 
                           A_neg_shifted_by1_14_50_port, INPUT(270) => 
                           A_neg_shifted_by1_14_49_port, INPUT(271) => 
                           A_neg_shifted_by1_14_48_port, INPUT(272) => 
                           A_neg_shifted_by1_14_47_port, INPUT(273) => 
                           A_neg_shifted_by1_14_46_port, INPUT(274) => 
                           A_neg_shifted_by1_14_45_port, INPUT(275) => 
                           A_neg_shifted_by1_14_44_port, INPUT(276) => 
                           A_neg_shifted_by1_14_43_port, INPUT(277) => 
                           A_neg_shifted_by1_14_42_port, INPUT(278) => 
                           A_neg_shifted_by1_14_41_port, INPUT(279) => 
                           A_neg_shifted_by1_14_40_port, INPUT(280) => 
                           A_neg_shifted_by1_14_39_port, INPUT(281) => 
                           A_neg_shifted_by1_14_38_port, INPUT(282) => 
                           A_neg_shifted_by1_14_37_port, INPUT(283) => 
                           A_neg_shifted_by1_14_36_port, INPUT(284) => 
                           A_neg_shifted_by1_14_35_port, INPUT(285) => 
                           A_neg_shifted_by1_14_34_port, INPUT(286) => 
                           A_neg_shifted_by1_14_33_port, INPUT(287) => 
                           A_neg_shifted_by1_14_32_port, INPUT(288) => 
                           A_neg_shifted_by1_14_31_port, INPUT(289) => 
                           A_neg_shifted_by1_14_30_port, INPUT(290) => 
                           A_neg_shifted_by1_14_29_port, INPUT(291) => 
                           A_neg_shifted_by1_14_28_port, INPUT(292) => 
                           A_neg_shifted_by1_14_27_port, INPUT(293) => 
                           A_neg_shifted_by1_14_26_port, INPUT(294) => 
                           A_neg_shifted_by1_14_25_port, INPUT(295) => 
                           A_neg_shifted_by1_14_24_port, INPUT(296) => 
                           A_neg_shifted_by1_14_23_port, INPUT(297) => 
                           A_neg_shifted_by1_14_22_port, INPUT(298) => 
                           A_neg_shifted_by1_14_21_port, INPUT(299) => 
                           A_neg_shifted_by1_14_20_port, INPUT(300) => 
                           A_neg_shifted_by1_14_19_port, INPUT(301) => 
                           A_neg_shifted_by1_14_18_port, INPUT(302) => 
                           A_neg_shifted_by1_14_17_port, INPUT(303) => 
                           A_neg_shifted_by1_14_16_port, INPUT(304) => 
                           A_neg_shifted_by1_14_15_port, INPUT(305) => 
                           A_neg_shifted_by1_14_14_port, INPUT(306) => 
                           A_neg_shifted_by1_14_13_port, INPUT(307) => 
                           A_neg_shifted_by1_14_12_port, INPUT(308) => 
                           A_neg_shifted_by1_14_11_port, INPUT(309) => 
                           A_neg_shifted_by1_14_10_port, INPUT(310) => 
                           A_neg_shifted_by1_14_9_port, INPUT(311) => 
                           A_neg_shifted_by1_14_8_port, INPUT(312) => 
                           A_neg_shifted_by1_14_7_port, INPUT(313) => 
                           A_neg_shifted_by1_14_6_port, INPUT(314) => 
                           A_neg_shifted_by1_14_5_port, INPUT(315) => 
                           A_neg_shifted_by1_14_4_port, INPUT(316) => 
                           A_neg_shifted_by1_14_3_port, INPUT(317) => 
                           A_neg_shifted_by1_14_2_port, INPUT(318) => 
                           A_neg_shifted_by1_14_1_port, INPUT(319) => 
                           A_neg_shifted_by1_14_0_port, SEL(0) => 
                           selection_signal_14_2_port, SEL(1) => 
                           selection_signal_14_1_port, SEL(2) => 
                           selection_signal_14_0_port, Y(0) => 
                           OUT_MUX_14_63_port, Y(1) => OUT_MUX_14_62_port, Y(2)
                           => OUT_MUX_14_61_port, Y(3) => OUT_MUX_14_60_port, 
                           Y(4) => OUT_MUX_14_59_port, Y(5) => 
                           OUT_MUX_14_58_port, Y(6) => OUT_MUX_14_57_port, Y(7)
                           => OUT_MUX_14_56_port, Y(8) => OUT_MUX_14_55_port, 
                           Y(9) => OUT_MUX_14_54_port, Y(10) => 
                           OUT_MUX_14_53_port, Y(11) => OUT_MUX_14_52_port, 
                           Y(12) => OUT_MUX_14_51_port, Y(13) => 
                           OUT_MUX_14_50_port, Y(14) => OUT_MUX_14_49_port, 
                           Y(15) => OUT_MUX_14_48_port, Y(16) => 
                           OUT_MUX_14_47_port, Y(17) => OUT_MUX_14_46_port, 
                           Y(18) => OUT_MUX_14_45_port, Y(19) => 
                           OUT_MUX_14_44_port, Y(20) => OUT_MUX_14_43_port, 
                           Y(21) => OUT_MUX_14_42_port, Y(22) => 
                           OUT_MUX_14_41_port, Y(23) => OUT_MUX_14_40_port, 
                           Y(24) => OUT_MUX_14_39_port, Y(25) => 
                           OUT_MUX_14_38_port, Y(26) => OUT_MUX_14_37_port, 
                           Y(27) => OUT_MUX_14_36_port, Y(28) => 
                           OUT_MUX_14_35_port, Y(29) => OUT_MUX_14_34_port, 
                           Y(30) => OUT_MUX_14_33_port, Y(31) => 
                           OUT_MUX_14_32_port, Y(32) => OUT_MUX_14_31_port, 
                           Y(33) => OUT_MUX_14_30_port, Y(34) => 
                           OUT_MUX_14_29_port, Y(35) => OUT_MUX_14_28_port, 
                           Y(36) => OUT_MUX_14_27_port, Y(37) => 
                           OUT_MUX_14_26_port, Y(38) => OUT_MUX_14_25_port, 
                           Y(39) => OUT_MUX_14_24_port, Y(40) => 
                           OUT_MUX_14_23_port, Y(41) => OUT_MUX_14_22_port, 
                           Y(42) => OUT_MUX_14_21_port, Y(43) => 
                           OUT_MUX_14_20_port, Y(44) => OUT_MUX_14_19_port, 
                           Y(45) => OUT_MUX_14_18_port, Y(46) => 
                           OUT_MUX_14_17_port, Y(47) => OUT_MUX_14_16_port, 
                           Y(48) => OUT_MUX_14_15_port, Y(49) => 
                           OUT_MUX_14_14_port, Y(50) => OUT_MUX_14_13_port, 
                           Y(51) => OUT_MUX_14_12_port, Y(52) => 
                           OUT_MUX_14_11_port, Y(53) => OUT_MUX_14_10_port, 
                           Y(54) => OUT_MUX_14_9_port, Y(55) => 
                           OUT_MUX_14_8_port, Y(56) => OUT_MUX_14_7_port, Y(57)
                           => OUT_MUX_14_6_port, Y(58) => OUT_MUX_14_5_port, 
                           Y(59) => OUT_MUX_14_4_port, Y(60) => 
                           OUT_MUX_14_3_port, Y(61) => OUT_MUX_14_2_port, Y(62)
                           => OUT_MUX_14_1_port, Y(63) => OUT_MUX_14_0_port);
   MUXi_15 : MUX_GENERIC_NBIT64_INPUTS5_NBIT_SEL3_1 port map( INPUT(0) => 
                           X_Logic0_port, INPUT(1) => X_Logic0_port, INPUT(2) 
                           => X_Logic0_port, INPUT(3) => X_Logic0_port, 
                           INPUT(4) => X_Logic0_port, INPUT(5) => X_Logic0_port
                           , INPUT(6) => X_Logic0_port, INPUT(7) => 
                           X_Logic0_port, INPUT(8) => X_Logic0_port, INPUT(9) 
                           => X_Logic0_port, INPUT(10) => X_Logic0_port, 
                           INPUT(11) => X_Logic0_port, INPUT(12) => 
                           X_Logic0_port, INPUT(13) => X_Logic0_port, INPUT(14)
                           => X_Logic0_port, INPUT(15) => X_Logic0_port, 
                           INPUT(16) => X_Logic0_port, INPUT(17) => 
                           X_Logic0_port, INPUT(18) => X_Logic0_port, INPUT(19)
                           => X_Logic0_port, INPUT(20) => X_Logic0_port, 
                           INPUT(21) => X_Logic0_port, INPUT(22) => 
                           X_Logic0_port, INPUT(23) => X_Logic0_port, INPUT(24)
                           => X_Logic0_port, INPUT(25) => X_Logic0_port, 
                           INPUT(26) => X_Logic0_port, INPUT(27) => 
                           X_Logic0_port, INPUT(28) => X_Logic0_port, INPUT(29)
                           => X_Logic0_port, INPUT(30) => X_Logic0_port, 
                           INPUT(31) => X_Logic0_port, INPUT(32) => 
                           X_Logic0_port, INPUT(33) => X_Logic0_port, INPUT(34)
                           => X_Logic0_port, INPUT(35) => X_Logic0_port, 
                           INPUT(36) => X_Logic0_port, INPUT(37) => 
                           X_Logic0_port, INPUT(38) => X_Logic0_port, INPUT(39)
                           => X_Logic0_port, INPUT(40) => X_Logic0_port, 
                           INPUT(41) => X_Logic0_port, INPUT(42) => 
                           X_Logic0_port, INPUT(43) => X_Logic0_port, INPUT(44)
                           => X_Logic0_port, INPUT(45) => X_Logic0_port, 
                           INPUT(46) => X_Logic0_port, INPUT(47) => 
                           X_Logic0_port, INPUT(48) => X_Logic0_port, INPUT(49)
                           => X_Logic0_port, INPUT(50) => X_Logic0_port, 
                           INPUT(51) => X_Logic0_port, INPUT(52) => 
                           X_Logic0_port, INPUT(53) => X_Logic0_port, INPUT(54)
                           => X_Logic0_port, INPUT(55) => X_Logic0_port, 
                           INPUT(56) => X_Logic0_port, INPUT(57) => 
                           X_Logic0_port, INPUT(58) => X_Logic0_port, INPUT(59)
                           => X_Logic0_port, INPUT(60) => X_Logic0_port, 
                           INPUT(61) => X_Logic0_port, INPUT(62) => 
                           X_Logic0_port, INPUT(63) => X_Logic0_port, INPUT(64)
                           => A_pos_shifted_by2_14_63_port, INPUT(65) => 
                           A_pos_shifted_by2_14_62_port, INPUT(66) => 
                           A_pos_shifted_by2_14_61_port, INPUT(67) => 
                           A_pos_shifted_by2_14_60_port, INPUT(68) => 
                           A_pos_shifted_by2_14_59_port, INPUT(69) => 
                           A_pos_shifted_by2_14_58_port, INPUT(70) => 
                           A_pos_shifted_by2_14_57_port, INPUT(71) => 
                           A_pos_shifted_by2_14_56_port, INPUT(72) => 
                           A_pos_shifted_by2_14_55_port, INPUT(73) => 
                           A_pos_shifted_by2_14_54_port, INPUT(74) => 
                           A_pos_shifted_by2_14_53_port, INPUT(75) => 
                           A_pos_shifted_by2_14_52_port, INPUT(76) => 
                           A_pos_shifted_by2_14_51_port, INPUT(77) => 
                           A_pos_shifted_by2_14_50_port, INPUT(78) => 
                           A_pos_shifted_by2_14_49_port, INPUT(79) => 
                           A_pos_shifted_by2_14_48_port, INPUT(80) => 
                           A_pos_shifted_by2_14_47_port, INPUT(81) => 
                           A_pos_shifted_by2_14_46_port, INPUT(82) => 
                           A_pos_shifted_by2_14_45_port, INPUT(83) => 
                           A_pos_shifted_by2_14_44_port, INPUT(84) => 
                           A_pos_shifted_by2_14_43_port, INPUT(85) => 
                           A_pos_shifted_by2_14_42_port, INPUT(86) => 
                           A_pos_shifted_by2_14_41_port, INPUT(87) => 
                           A_pos_shifted_by2_14_40_port, INPUT(88) => 
                           A_pos_shifted_by2_14_39_port, INPUT(89) => 
                           A_pos_shifted_by2_14_38_port, INPUT(90) => 
                           A_pos_shifted_by2_14_37_port, INPUT(91) => 
                           A_pos_shifted_by2_14_36_port, INPUT(92) => 
                           A_pos_shifted_by2_14_35_port, INPUT(93) => 
                           A_pos_shifted_by2_14_34_port, INPUT(94) => 
                           A_pos_shifted_by2_14_33_port, INPUT(95) => 
                           A_pos_shifted_by2_14_32_port, INPUT(96) => 
                           A_pos_shifted_by2_14_31_port, INPUT(97) => 
                           A_pos_shifted_by2_14_30_port, INPUT(98) => 
                           A_pos_shifted_by2_14_29_port, INPUT(99) => 
                           A_pos_shifted_by2_14_28_port, INPUT(100) => 
                           A_pos_shifted_by2_14_27_port, INPUT(101) => 
                           A_pos_shifted_by2_14_26_port, INPUT(102) => 
                           A_pos_shifted_by2_14_25_port, INPUT(103) => 
                           A_pos_shifted_by2_14_24_port, INPUT(104) => 
                           A_pos_shifted_by2_14_23_port, INPUT(105) => 
                           A_pos_shifted_by2_14_22_port, INPUT(106) => 
                           A_pos_shifted_by2_14_21_port, INPUT(107) => 
                           A_pos_shifted_by2_14_20_port, INPUT(108) => 
                           A_pos_shifted_by2_14_19_port, INPUT(109) => 
                           A_pos_shifted_by2_14_18_port, INPUT(110) => 
                           A_pos_shifted_by2_14_17_port, INPUT(111) => 
                           A_pos_shifted_by2_14_16_port, INPUT(112) => 
                           A_pos_shifted_by2_14_15_port, INPUT(113) => 
                           A_pos_shifted_by2_14_14_port, INPUT(114) => 
                           A_pos_shifted_by2_14_13_port, INPUT(115) => 
                           A_pos_shifted_by2_14_12_port, INPUT(116) => 
                           A_pos_shifted_by2_14_11_port, INPUT(117) => 
                           A_pos_shifted_by2_14_10_port, INPUT(118) => 
                           A_pos_shifted_by2_14_9_port, INPUT(119) => 
                           A_pos_shifted_by2_14_8_port, INPUT(120) => 
                           A_pos_shifted_by2_14_7_port, INPUT(121) => 
                           A_pos_shifted_by2_14_6_port, INPUT(122) => 
                           A_pos_shifted_by2_14_5_port, INPUT(123) => 
                           A_pos_shifted_by2_14_4_port, INPUT(124) => 
                           A_pos_shifted_by2_14_3_port, INPUT(125) => 
                           A_pos_shifted_by2_14_2_port, INPUT(126) => 
                           A_pos_shifted_by2_14_1_port, INPUT(127) => 
                           A_pos_shifted_by2_14_0_port, INPUT(128) => 
                           A_neg_shifted_by2_14_63_port, INPUT(129) => 
                           A_neg_shifted_by2_14_62_port, INPUT(130) => 
                           A_neg_shifted_by2_14_61_port, INPUT(131) => 
                           A_neg_shifted_by2_14_60_port, INPUT(132) => 
                           A_neg_shifted_by2_14_59_port, INPUT(133) => 
                           A_neg_shifted_by2_14_58_port, INPUT(134) => 
                           A_neg_shifted_by2_14_57_port, INPUT(135) => 
                           A_neg_shifted_by2_14_56_port, INPUT(136) => 
                           A_neg_shifted_by2_14_55_port, INPUT(137) => 
                           A_neg_shifted_by2_14_54_port, INPUT(138) => 
                           A_neg_shifted_by2_14_53_port, INPUT(139) => 
                           A_neg_shifted_by2_14_52_port, INPUT(140) => 
                           A_neg_shifted_by2_14_51_port, INPUT(141) => 
                           A_neg_shifted_by2_14_50_port, INPUT(142) => 
                           A_neg_shifted_by2_14_49_port, INPUT(143) => 
                           A_neg_shifted_by2_14_48_port, INPUT(144) => 
                           A_neg_shifted_by2_14_47_port, INPUT(145) => 
                           A_neg_shifted_by2_14_46_port, INPUT(146) => 
                           A_neg_shifted_by2_14_45_port, INPUT(147) => 
                           A_neg_shifted_by2_14_44_port, INPUT(148) => 
                           A_neg_shifted_by2_14_43_port, INPUT(149) => 
                           A_neg_shifted_by2_14_42_port, INPUT(150) => 
                           A_neg_shifted_by2_14_41_port, INPUT(151) => 
                           A_neg_shifted_by2_14_40_port, INPUT(152) => 
                           A_neg_shifted_by2_14_39_port, INPUT(153) => 
                           A_neg_shifted_by2_14_38_port, INPUT(154) => 
                           A_neg_shifted_by2_14_37_port, INPUT(155) => 
                           A_neg_shifted_by2_14_36_port, INPUT(156) => 
                           A_neg_shifted_by2_14_35_port, INPUT(157) => 
                           A_neg_shifted_by2_14_34_port, INPUT(158) => 
                           A_neg_shifted_by2_14_33_port, INPUT(159) => 
                           A_neg_shifted_by2_14_32_port, INPUT(160) => 
                           A_neg_shifted_by2_14_31_port, INPUT(161) => 
                           A_neg_shifted_by2_14_30_port, INPUT(162) => 
                           A_neg_shifted_by2_14_29_port, INPUT(163) => 
                           A_neg_shifted_by2_14_28_port, INPUT(164) => 
                           A_neg_shifted_by2_14_27_port, INPUT(165) => 
                           A_neg_shifted_by2_14_26_port, INPUT(166) => 
                           A_neg_shifted_by2_14_25_port, INPUT(167) => 
                           A_neg_shifted_by2_14_24_port, INPUT(168) => 
                           A_neg_shifted_by2_14_23_port, INPUT(169) => 
                           A_neg_shifted_by2_14_22_port, INPUT(170) => 
                           A_neg_shifted_by2_14_21_port, INPUT(171) => 
                           A_neg_shifted_by2_14_20_port, INPUT(172) => 
                           A_neg_shifted_by2_14_19_port, INPUT(173) => 
                           A_neg_shifted_by2_14_18_port, INPUT(174) => 
                           A_neg_shifted_by2_14_17_port, INPUT(175) => 
                           A_neg_shifted_by2_14_16_port, INPUT(176) => 
                           A_neg_shifted_by2_14_15_port, INPUT(177) => 
                           A_neg_shifted_by2_14_14_port, INPUT(178) => 
                           A_neg_shifted_by2_14_13_port, INPUT(179) => 
                           A_neg_shifted_by2_14_12_port, INPUT(180) => 
                           A_neg_shifted_by2_14_11_port, INPUT(181) => 
                           A_neg_shifted_by2_14_10_port, INPUT(182) => 
                           A_neg_shifted_by2_14_9_port, INPUT(183) => 
                           A_neg_shifted_by2_14_8_port, INPUT(184) => 
                           A_neg_shifted_by2_14_7_port, INPUT(185) => 
                           A_neg_shifted_by2_14_6_port, INPUT(186) => 
                           A_neg_shifted_by2_14_5_port, INPUT(187) => 
                           A_neg_shifted_by2_14_4_port, INPUT(188) => 
                           A_neg_shifted_by2_14_3_port, INPUT(189) => 
                           A_neg_shifted_by2_14_2_port, INPUT(190) => 
                           A_neg_shifted_by2_14_1_port, INPUT(191) => 
                           A_neg_shifted_by2_14_0_port, INPUT(192) => 
                           A_pos_shifted_by1_15_63_port, INPUT(193) => 
                           A_pos_shifted_by1_15_62_port, INPUT(194) => 
                           A_pos_shifted_by1_15_61_port, INPUT(195) => 
                           A_pos_shifted_by1_15_60_port, INPUT(196) => 
                           A_pos_shifted_by1_15_59_port, INPUT(197) => 
                           A_pos_shifted_by1_15_58_port, INPUT(198) => 
                           A_pos_shifted_by1_15_57_port, INPUT(199) => 
                           A_pos_shifted_by1_15_56_port, INPUT(200) => 
                           A_pos_shifted_by1_15_55_port, INPUT(201) => 
                           A_pos_shifted_by1_15_54_port, INPUT(202) => 
                           A_pos_shifted_by1_15_53_port, INPUT(203) => 
                           A_pos_shifted_by1_15_52_port, INPUT(204) => 
                           A_pos_shifted_by1_15_51_port, INPUT(205) => 
                           A_pos_shifted_by1_15_50_port, INPUT(206) => 
                           A_pos_shifted_by1_15_49_port, INPUT(207) => 
                           A_pos_shifted_by1_15_48_port, INPUT(208) => 
                           A_pos_shifted_by1_15_47_port, INPUT(209) => 
                           A_pos_shifted_by1_15_46_port, INPUT(210) => 
                           A_pos_shifted_by1_15_45_port, INPUT(211) => 
                           A_pos_shifted_by1_15_44_port, INPUT(212) => 
                           A_pos_shifted_by1_15_43_port, INPUT(213) => 
                           A_pos_shifted_by1_15_42_port, INPUT(214) => 
                           A_pos_shifted_by1_15_41_port, INPUT(215) => 
                           A_pos_shifted_by1_15_40_port, INPUT(216) => 
                           A_pos_shifted_by1_15_39_port, INPUT(217) => 
                           A_pos_shifted_by1_15_38_port, INPUT(218) => 
                           A_pos_shifted_by1_15_37_port, INPUT(219) => 
                           A_pos_shifted_by1_15_36_port, INPUT(220) => 
                           A_pos_shifted_by1_15_35_port, INPUT(221) => 
                           A_pos_shifted_by1_15_34_port, INPUT(222) => 
                           A_pos_shifted_by1_15_33_port, INPUT(223) => 
                           A_pos_shifted_by1_15_32_port, INPUT(224) => 
                           A_pos_shifted_by1_15_31_port, INPUT(225) => 
                           A_pos_shifted_by1_15_30_port, INPUT(226) => 
                           A_pos_shifted_by1_15_29_port, INPUT(227) => 
                           A_pos_shifted_by1_15_28_port, INPUT(228) => 
                           A_pos_shifted_by1_15_27_port, INPUT(229) => 
                           A_pos_shifted_by1_15_26_port, INPUT(230) => 
                           A_pos_shifted_by1_15_25_port, INPUT(231) => 
                           A_pos_shifted_by1_15_24_port, INPUT(232) => 
                           A_pos_shifted_by1_15_23_port, INPUT(233) => 
                           A_pos_shifted_by1_15_22_port, INPUT(234) => 
                           A_pos_shifted_by1_15_21_port, INPUT(235) => 
                           A_pos_shifted_by1_15_20_port, INPUT(236) => 
                           A_pos_shifted_by1_15_19_port, INPUT(237) => 
                           A_pos_shifted_by1_15_18_port, INPUT(238) => 
                           A_pos_shifted_by1_15_17_port, INPUT(239) => 
                           A_pos_shifted_by1_15_16_port, INPUT(240) => 
                           A_pos_shifted_by1_15_15_port, INPUT(241) => 
                           A_pos_shifted_by1_15_14_port, INPUT(242) => 
                           A_pos_shifted_by1_15_13_port, INPUT(243) => 
                           A_pos_shifted_by1_15_12_port, INPUT(244) => 
                           A_pos_shifted_by1_15_11_port, INPUT(245) => 
                           A_pos_shifted_by1_15_10_port, INPUT(246) => 
                           A_pos_shifted_by1_15_9_port, INPUT(247) => 
                           A_pos_shifted_by1_15_8_port, INPUT(248) => 
                           A_pos_shifted_by1_15_7_port, INPUT(249) => 
                           A_pos_shifted_by1_15_6_port, INPUT(250) => 
                           A_pos_shifted_by1_15_5_port, INPUT(251) => 
                           A_pos_shifted_by1_15_4_port, INPUT(252) => 
                           A_pos_shifted_by1_15_3_port, INPUT(253) => 
                           A_pos_shifted_by1_15_2_port, INPUT(254) => 
                           A_pos_shifted_by1_15_1_port, INPUT(255) => 
                           A_pos_shifted_by1_15_0_port, INPUT(256) => 
                           A_neg_shifted_by1_15_63_port, INPUT(257) => 
                           A_neg_shifted_by1_15_62_port, INPUT(258) => 
                           A_neg_shifted_by1_15_61_port, INPUT(259) => 
                           A_neg_shifted_by1_15_60_port, INPUT(260) => 
                           A_neg_shifted_by1_15_59_port, INPUT(261) => 
                           A_neg_shifted_by1_15_58_port, INPUT(262) => 
                           A_neg_shifted_by1_15_57_port, INPUT(263) => 
                           A_neg_shifted_by1_15_56_port, INPUT(264) => 
                           A_neg_shifted_by1_15_55_port, INPUT(265) => 
                           A_neg_shifted_by1_15_54_port, INPUT(266) => 
                           A_neg_shifted_by1_15_53_port, INPUT(267) => 
                           A_neg_shifted_by1_15_52_port, INPUT(268) => 
                           A_neg_shifted_by1_15_51_port, INPUT(269) => 
                           A_neg_shifted_by1_15_50_port, INPUT(270) => 
                           A_neg_shifted_by1_15_49_port, INPUT(271) => 
                           A_neg_shifted_by1_15_48_port, INPUT(272) => 
                           A_neg_shifted_by1_15_47_port, INPUT(273) => 
                           A_neg_shifted_by1_15_46_port, INPUT(274) => 
                           A_neg_shifted_by1_15_45_port, INPUT(275) => 
                           A_neg_shifted_by1_15_44_port, INPUT(276) => 
                           A_neg_shifted_by1_15_43_port, INPUT(277) => 
                           A_neg_shifted_by1_15_42_port, INPUT(278) => 
                           A_neg_shifted_by1_15_41_port, INPUT(279) => 
                           A_neg_shifted_by1_15_40_port, INPUT(280) => 
                           A_neg_shifted_by1_15_39_port, INPUT(281) => 
                           A_neg_shifted_by1_15_38_port, INPUT(282) => 
                           A_neg_shifted_by1_15_37_port, INPUT(283) => 
                           A_neg_shifted_by1_15_36_port, INPUT(284) => 
                           A_neg_shifted_by1_15_35_port, INPUT(285) => 
                           A_neg_shifted_by1_15_34_port, INPUT(286) => 
                           A_neg_shifted_by1_15_33_port, INPUT(287) => 
                           A_neg_shifted_by1_15_32_port, INPUT(288) => 
                           A_neg_shifted_by1_15_31_port, INPUT(289) => 
                           A_neg_shifted_by1_15_30_port, INPUT(290) => 
                           A_neg_shifted_by1_15_29_port, INPUT(291) => 
                           A_neg_shifted_by1_15_28_port, INPUT(292) => 
                           A_neg_shifted_by1_15_27_port, INPUT(293) => 
                           A_neg_shifted_by1_15_26_port, INPUT(294) => 
                           A_neg_shifted_by1_15_25_port, INPUT(295) => 
                           A_neg_shifted_by1_15_24_port, INPUT(296) => 
                           A_neg_shifted_by1_15_23_port, INPUT(297) => 
                           A_neg_shifted_by1_15_22_port, INPUT(298) => 
                           A_neg_shifted_by1_15_21_port, INPUT(299) => 
                           A_neg_shifted_by1_15_20_port, INPUT(300) => 
                           A_neg_shifted_by1_15_19_port, INPUT(301) => 
                           A_neg_shifted_by1_15_18_port, INPUT(302) => 
                           A_neg_shifted_by1_15_17_port, INPUT(303) => 
                           A_neg_shifted_by1_15_16_port, INPUT(304) => 
                           A_neg_shifted_by1_15_15_port, INPUT(305) => 
                           A_neg_shifted_by1_15_14_port, INPUT(306) => 
                           A_neg_shifted_by1_15_13_port, INPUT(307) => 
                           A_neg_shifted_by1_15_12_port, INPUT(308) => 
                           A_neg_shifted_by1_15_11_port, INPUT(309) => 
                           A_neg_shifted_by1_15_10_port, INPUT(310) => 
                           A_neg_shifted_by1_15_9_port, INPUT(311) => 
                           A_neg_shifted_by1_15_8_port, INPUT(312) => 
                           A_neg_shifted_by1_15_7_port, INPUT(313) => 
                           A_neg_shifted_by1_15_6_port, INPUT(314) => 
                           A_neg_shifted_by1_15_5_port, INPUT(315) => 
                           A_neg_shifted_by1_15_4_port, INPUT(316) => 
                           A_neg_shifted_by1_15_3_port, INPUT(317) => 
                           A_neg_shifted_by1_15_2_port, INPUT(318) => 
                           A_neg_shifted_by1_15_1_port, INPUT(319) => 
                           A_neg_shifted_by1_15_0_port, SEL(0) => 
                           selection_signal_15_2_port, SEL(1) => 
                           selection_signal_15_1_port, SEL(2) => 
                           selection_signal_15_0_port, Y(0) => 
                           OUT_MUX_15_63_port, Y(1) => OUT_MUX_15_62_port, Y(2)
                           => OUT_MUX_15_61_port, Y(3) => OUT_MUX_15_60_port, 
                           Y(4) => OUT_MUX_15_59_port, Y(5) => 
                           OUT_MUX_15_58_port, Y(6) => OUT_MUX_15_57_port, Y(7)
                           => OUT_MUX_15_56_port, Y(8) => OUT_MUX_15_55_port, 
                           Y(9) => OUT_MUX_15_54_port, Y(10) => 
                           OUT_MUX_15_53_port, Y(11) => OUT_MUX_15_52_port, 
                           Y(12) => OUT_MUX_15_51_port, Y(13) => 
                           OUT_MUX_15_50_port, Y(14) => OUT_MUX_15_49_port, 
                           Y(15) => OUT_MUX_15_48_port, Y(16) => 
                           OUT_MUX_15_47_port, Y(17) => OUT_MUX_15_46_port, 
                           Y(18) => OUT_MUX_15_45_port, Y(19) => 
                           OUT_MUX_15_44_port, Y(20) => OUT_MUX_15_43_port, 
                           Y(21) => OUT_MUX_15_42_port, Y(22) => 
                           OUT_MUX_15_41_port, Y(23) => OUT_MUX_15_40_port, 
                           Y(24) => OUT_MUX_15_39_port, Y(25) => 
                           OUT_MUX_15_38_port, Y(26) => OUT_MUX_15_37_port, 
                           Y(27) => OUT_MUX_15_36_port, Y(28) => 
                           OUT_MUX_15_35_port, Y(29) => OUT_MUX_15_34_port, 
                           Y(30) => OUT_MUX_15_33_port, Y(31) => 
                           OUT_MUX_15_32_port, Y(32) => OUT_MUX_15_31_port, 
                           Y(33) => OUT_MUX_15_30_port, Y(34) => 
                           OUT_MUX_15_29_port, Y(35) => OUT_MUX_15_28_port, 
                           Y(36) => OUT_MUX_15_27_port, Y(37) => 
                           OUT_MUX_15_26_port, Y(38) => OUT_MUX_15_25_port, 
                           Y(39) => OUT_MUX_15_24_port, Y(40) => 
                           OUT_MUX_15_23_port, Y(41) => OUT_MUX_15_22_port, 
                           Y(42) => OUT_MUX_15_21_port, Y(43) => 
                           OUT_MUX_15_20_port, Y(44) => OUT_MUX_15_19_port, 
                           Y(45) => OUT_MUX_15_18_port, Y(46) => 
                           OUT_MUX_15_17_port, Y(47) => OUT_MUX_15_16_port, 
                           Y(48) => OUT_MUX_15_15_port, Y(49) => 
                           OUT_MUX_15_14_port, Y(50) => OUT_MUX_15_13_port, 
                           Y(51) => OUT_MUX_15_12_port, Y(52) => 
                           OUT_MUX_15_11_port, Y(53) => OUT_MUX_15_10_port, 
                           Y(54) => OUT_MUX_15_9_port, Y(55) => 
                           OUT_MUX_15_8_port, Y(56) => OUT_MUX_15_7_port, Y(57)
                           => OUT_MUX_15_6_port, Y(58) => OUT_MUX_15_5_port, 
                           Y(59) => OUT_MUX_15_4_port, Y(60) => 
                           OUT_MUX_15_3_port, Y(61) => OUT_MUX_15_2_port, Y(62)
                           => OUT_MUX_15_1_port, Y(63) => OUT_MUX_15_0_port);
   RCAi_0 : RCA_NBIT64_0 port map( A(63) => P_tmp_0_63_port, A(62) => 
                           P_tmp_0_62_port, A(61) => P_tmp_0_61_port, A(60) => 
                           P_tmp_0_60_port, A(59) => P_tmp_0_59_port, A(58) => 
                           P_tmp_0_58_port, A(57) => P_tmp_0_57_port, A(56) => 
                           P_tmp_0_56_port, A(55) => P_tmp_0_55_port, A(54) => 
                           P_tmp_0_54_port, A(53) => P_tmp_0_53_port, A(52) => 
                           P_tmp_0_52_port, A(51) => P_tmp_0_51_port, A(50) => 
                           P_tmp_0_50_port, A(49) => P_tmp_0_49_port, A(48) => 
                           P_tmp_0_48_port, A(47) => P_tmp_0_47_port, A(46) => 
                           P_tmp_0_46_port, A(45) => P_tmp_0_45_port, A(44) => 
                           P_tmp_0_44_port, A(43) => P_tmp_0_43_port, A(42) => 
                           P_tmp_0_42_port, A(41) => P_tmp_0_41_port, A(40) => 
                           P_tmp_0_40_port, A(39) => P_tmp_0_39_port, A(38) => 
                           P_tmp_0_38_port, A(37) => P_tmp_0_37_port, A(36) => 
                           P_tmp_0_36_port, A(35) => P_tmp_0_35_port, A(34) => 
                           P_tmp_0_34_port, A(33) => P_tmp_0_33_port, A(32) => 
                           P_tmp_0_32_port, A(31) => P_tmp_0_31_port, A(30) => 
                           P_tmp_0_30_port, A(29) => P_tmp_0_29_port, A(28) => 
                           P_tmp_0_28_port, A(27) => P_tmp_0_27_port, A(26) => 
                           P_tmp_0_26_port, A(25) => P_tmp_0_25_port, A(24) => 
                           P_tmp_0_24_port, A(23) => P_tmp_0_23_port, A(22) => 
                           P_tmp_0_22_port, A(21) => P_tmp_0_21_port, A(20) => 
                           P_tmp_0_20_port, A(19) => P_tmp_0_19_port, A(18) => 
                           P_tmp_0_18_port, A(17) => P_tmp_0_17_port, A(16) => 
                           P_tmp_0_16_port, A(15) => P_tmp_0_15_port, A(14) => 
                           P_tmp_0_14_port, A(13) => P_tmp_0_13_port, A(12) => 
                           P_tmp_0_12_port, A(11) => P_tmp_0_11_port, A(10) => 
                           P_tmp_0_10_port, A(9) => P_tmp_0_9_port, A(8) => 
                           P_tmp_0_8_port, A(7) => P_tmp_0_7_port, A(6) => 
                           P_tmp_0_6_port, A(5) => P_tmp_0_5_port, A(4) => 
                           P_tmp_0_4_port, A(3) => P_tmp_0_3_port, A(2) => 
                           P_tmp_0_2_port, A(1) => P_tmp_0_1_port, A(0) => 
                           P_tmp_0_0_port, B(63) => OUT_MUX_1_63_port, B(62) =>
                           OUT_MUX_1_62_port, B(61) => OUT_MUX_1_61_port, B(60)
                           => OUT_MUX_1_60_port, B(59) => OUT_MUX_1_59_port, 
                           B(58) => OUT_MUX_1_58_port, B(57) => 
                           OUT_MUX_1_57_port, B(56) => OUT_MUX_1_56_port, B(55)
                           => OUT_MUX_1_55_port, B(54) => OUT_MUX_1_54_port, 
                           B(53) => OUT_MUX_1_53_port, B(52) => 
                           OUT_MUX_1_52_port, B(51) => OUT_MUX_1_51_port, B(50)
                           => OUT_MUX_1_50_port, B(49) => OUT_MUX_1_49_port, 
                           B(48) => OUT_MUX_1_48_port, B(47) => 
                           OUT_MUX_1_47_port, B(46) => OUT_MUX_1_46_port, B(45)
                           => OUT_MUX_1_45_port, B(44) => OUT_MUX_1_44_port, 
                           B(43) => OUT_MUX_1_43_port, B(42) => 
                           OUT_MUX_1_42_port, B(41) => OUT_MUX_1_41_port, B(40)
                           => OUT_MUX_1_40_port, B(39) => OUT_MUX_1_39_port, 
                           B(38) => OUT_MUX_1_38_port, B(37) => 
                           OUT_MUX_1_37_port, B(36) => OUT_MUX_1_36_port, B(35)
                           => OUT_MUX_1_35_port, B(34) => OUT_MUX_1_34_port, 
                           B(33) => OUT_MUX_1_33_port, B(32) => 
                           OUT_MUX_1_32_port, B(31) => OUT_MUX_1_31_port, B(30)
                           => OUT_MUX_1_30_port, B(29) => OUT_MUX_1_29_port, 
                           B(28) => OUT_MUX_1_28_port, B(27) => 
                           OUT_MUX_1_27_port, B(26) => OUT_MUX_1_26_port, B(25)
                           => OUT_MUX_1_25_port, B(24) => OUT_MUX_1_24_port, 
                           B(23) => OUT_MUX_1_23_port, B(22) => 
                           OUT_MUX_1_22_port, B(21) => OUT_MUX_1_21_port, B(20)
                           => OUT_MUX_1_20_port, B(19) => OUT_MUX_1_19_port, 
                           B(18) => OUT_MUX_1_18_port, B(17) => 
                           OUT_MUX_1_17_port, B(16) => OUT_MUX_1_16_port, B(15)
                           => OUT_MUX_1_15_port, B(14) => OUT_MUX_1_14_port, 
                           B(13) => OUT_MUX_1_13_port, B(12) => 
                           OUT_MUX_1_12_port, B(11) => OUT_MUX_1_11_port, B(10)
                           => OUT_MUX_1_10_port, B(9) => OUT_MUX_1_9_port, B(8)
                           => OUT_MUX_1_8_port, B(7) => OUT_MUX_1_7_port, B(6) 
                           => OUT_MUX_1_6_port, B(5) => OUT_MUX_1_5_port, B(4) 
                           => OUT_MUX_1_4_port, B(3) => OUT_MUX_1_3_port, B(2) 
                           => OUT_MUX_1_2_port, B(1) => OUT_MUX_1_1_port, B(0) 
                           => OUT_MUX_1_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_1_63_port, S(62) => P_tmp_1_62_port, S(61) => 
                           P_tmp_1_61_port, S(60) => P_tmp_1_60_port, S(59) => 
                           P_tmp_1_59_port, S(58) => P_tmp_1_58_port, S(57) => 
                           P_tmp_1_57_port, S(56) => P_tmp_1_56_port, S(55) => 
                           P_tmp_1_55_port, S(54) => P_tmp_1_54_port, S(53) => 
                           P_tmp_1_53_port, S(52) => P_tmp_1_52_port, S(51) => 
                           P_tmp_1_51_port, S(50) => P_tmp_1_50_port, S(49) => 
                           P_tmp_1_49_port, S(48) => P_tmp_1_48_port, S(47) => 
                           P_tmp_1_47_port, S(46) => P_tmp_1_46_port, S(45) => 
                           P_tmp_1_45_port, S(44) => P_tmp_1_44_port, S(43) => 
                           P_tmp_1_43_port, S(42) => P_tmp_1_42_port, S(41) => 
                           P_tmp_1_41_port, S(40) => P_tmp_1_40_port, S(39) => 
                           P_tmp_1_39_port, S(38) => P_tmp_1_38_port, S(37) => 
                           P_tmp_1_37_port, S(36) => P_tmp_1_36_port, S(35) => 
                           P_tmp_1_35_port, S(34) => P_tmp_1_34_port, S(33) => 
                           P_tmp_1_33_port, S(32) => P_tmp_1_32_port, S(31) => 
                           P_tmp_1_31_port, S(30) => P_tmp_1_30_port, S(29) => 
                           P_tmp_1_29_port, S(28) => P_tmp_1_28_port, S(27) => 
                           P_tmp_1_27_port, S(26) => P_tmp_1_26_port, S(25) => 
                           P_tmp_1_25_port, S(24) => P_tmp_1_24_port, S(23) => 
                           P_tmp_1_23_port, S(22) => P_tmp_1_22_port, S(21) => 
                           P_tmp_1_21_port, S(20) => P_tmp_1_20_port, S(19) => 
                           P_tmp_1_19_port, S(18) => P_tmp_1_18_port, S(17) => 
                           P_tmp_1_17_port, S(16) => P_tmp_1_16_port, S(15) => 
                           P_tmp_1_15_port, S(14) => P_tmp_1_14_port, S(13) => 
                           P_tmp_1_13_port, S(12) => P_tmp_1_12_port, S(11) => 
                           P_tmp_1_11_port, S(10) => P_tmp_1_10_port, S(9) => 
                           P_tmp_1_9_port, S(8) => P_tmp_1_8_port, S(7) => 
                           P_tmp_1_7_port, S(6) => P_tmp_1_6_port, S(5) => 
                           P_tmp_1_5_port, S(4) => P_tmp_1_4_port, S(3) => 
                           P_tmp_1_3_port, S(2) => P_tmp_1_2_port, S(1) => 
                           P_tmp_1_1_port, S(0) => P_tmp_1_0_port, Co => n_1280
                           );
   RCAi_1 : RCA_NBIT64_14 port map( A(63) => P_tmp_1_63_port, A(62) => 
                           P_tmp_1_62_port, A(61) => P_tmp_1_61_port, A(60) => 
                           P_tmp_1_60_port, A(59) => P_tmp_1_59_port, A(58) => 
                           P_tmp_1_58_port, A(57) => P_tmp_1_57_port, A(56) => 
                           P_tmp_1_56_port, A(55) => P_tmp_1_55_port, A(54) => 
                           P_tmp_1_54_port, A(53) => P_tmp_1_53_port, A(52) => 
                           P_tmp_1_52_port, A(51) => P_tmp_1_51_port, A(50) => 
                           P_tmp_1_50_port, A(49) => P_tmp_1_49_port, A(48) => 
                           P_tmp_1_48_port, A(47) => P_tmp_1_47_port, A(46) => 
                           P_tmp_1_46_port, A(45) => P_tmp_1_45_port, A(44) => 
                           P_tmp_1_44_port, A(43) => P_tmp_1_43_port, A(42) => 
                           P_tmp_1_42_port, A(41) => P_tmp_1_41_port, A(40) => 
                           P_tmp_1_40_port, A(39) => P_tmp_1_39_port, A(38) => 
                           P_tmp_1_38_port, A(37) => P_tmp_1_37_port, A(36) => 
                           P_tmp_1_36_port, A(35) => P_tmp_1_35_port, A(34) => 
                           P_tmp_1_34_port, A(33) => P_tmp_1_33_port, A(32) => 
                           P_tmp_1_32_port, A(31) => P_tmp_1_31_port, A(30) => 
                           P_tmp_1_30_port, A(29) => P_tmp_1_29_port, A(28) => 
                           P_tmp_1_28_port, A(27) => P_tmp_1_27_port, A(26) => 
                           P_tmp_1_26_port, A(25) => P_tmp_1_25_port, A(24) => 
                           P_tmp_1_24_port, A(23) => P_tmp_1_23_port, A(22) => 
                           P_tmp_1_22_port, A(21) => P_tmp_1_21_port, A(20) => 
                           P_tmp_1_20_port, A(19) => P_tmp_1_19_port, A(18) => 
                           P_tmp_1_18_port, A(17) => P_tmp_1_17_port, A(16) => 
                           P_tmp_1_16_port, A(15) => P_tmp_1_15_port, A(14) => 
                           P_tmp_1_14_port, A(13) => P_tmp_1_13_port, A(12) => 
                           P_tmp_1_12_port, A(11) => P_tmp_1_11_port, A(10) => 
                           P_tmp_1_10_port, A(9) => P_tmp_1_9_port, A(8) => 
                           P_tmp_1_8_port, A(7) => P_tmp_1_7_port, A(6) => 
                           P_tmp_1_6_port, A(5) => P_tmp_1_5_port, A(4) => 
                           P_tmp_1_4_port, A(3) => P_tmp_1_3_port, A(2) => 
                           P_tmp_1_2_port, A(1) => P_tmp_1_1_port, A(0) => 
                           P_tmp_1_0_port, B(63) => OUT_MUX_2_63_port, B(62) =>
                           OUT_MUX_2_62_port, B(61) => OUT_MUX_2_61_port, B(60)
                           => OUT_MUX_2_60_port, B(59) => OUT_MUX_2_59_port, 
                           B(58) => OUT_MUX_2_58_port, B(57) => 
                           OUT_MUX_2_57_port, B(56) => OUT_MUX_2_56_port, B(55)
                           => OUT_MUX_2_55_port, B(54) => OUT_MUX_2_54_port, 
                           B(53) => OUT_MUX_2_53_port, B(52) => 
                           OUT_MUX_2_52_port, B(51) => OUT_MUX_2_51_port, B(50)
                           => OUT_MUX_2_50_port, B(49) => OUT_MUX_2_49_port, 
                           B(48) => OUT_MUX_2_48_port, B(47) => 
                           OUT_MUX_2_47_port, B(46) => OUT_MUX_2_46_port, B(45)
                           => OUT_MUX_2_45_port, B(44) => OUT_MUX_2_44_port, 
                           B(43) => OUT_MUX_2_43_port, B(42) => 
                           OUT_MUX_2_42_port, B(41) => OUT_MUX_2_41_port, B(40)
                           => OUT_MUX_2_40_port, B(39) => OUT_MUX_2_39_port, 
                           B(38) => OUT_MUX_2_38_port, B(37) => 
                           OUT_MUX_2_37_port, B(36) => OUT_MUX_2_36_port, B(35)
                           => OUT_MUX_2_35_port, B(34) => OUT_MUX_2_34_port, 
                           B(33) => OUT_MUX_2_33_port, B(32) => 
                           OUT_MUX_2_32_port, B(31) => OUT_MUX_2_31_port, B(30)
                           => OUT_MUX_2_30_port, B(29) => OUT_MUX_2_29_port, 
                           B(28) => OUT_MUX_2_28_port, B(27) => 
                           OUT_MUX_2_27_port, B(26) => OUT_MUX_2_26_port, B(25)
                           => OUT_MUX_2_25_port, B(24) => OUT_MUX_2_24_port, 
                           B(23) => OUT_MUX_2_23_port, B(22) => 
                           OUT_MUX_2_22_port, B(21) => OUT_MUX_2_21_port, B(20)
                           => OUT_MUX_2_20_port, B(19) => OUT_MUX_2_19_port, 
                           B(18) => OUT_MUX_2_18_port, B(17) => 
                           OUT_MUX_2_17_port, B(16) => OUT_MUX_2_16_port, B(15)
                           => OUT_MUX_2_15_port, B(14) => OUT_MUX_2_14_port, 
                           B(13) => OUT_MUX_2_13_port, B(12) => 
                           OUT_MUX_2_12_port, B(11) => OUT_MUX_2_11_port, B(10)
                           => OUT_MUX_2_10_port, B(9) => OUT_MUX_2_9_port, B(8)
                           => OUT_MUX_2_8_port, B(7) => OUT_MUX_2_7_port, B(6) 
                           => OUT_MUX_2_6_port, B(5) => OUT_MUX_2_5_port, B(4) 
                           => OUT_MUX_2_4_port, B(3) => OUT_MUX_2_3_port, B(2) 
                           => OUT_MUX_2_2_port, B(1) => OUT_MUX_2_1_port, B(0) 
                           => OUT_MUX_2_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_2_63_port, S(62) => P_tmp_2_62_port, S(61) => 
                           P_tmp_2_61_port, S(60) => P_tmp_2_60_port, S(59) => 
                           P_tmp_2_59_port, S(58) => P_tmp_2_58_port, S(57) => 
                           P_tmp_2_57_port, S(56) => P_tmp_2_56_port, S(55) => 
                           P_tmp_2_55_port, S(54) => P_tmp_2_54_port, S(53) => 
                           P_tmp_2_53_port, S(52) => P_tmp_2_52_port, S(51) => 
                           P_tmp_2_51_port, S(50) => P_tmp_2_50_port, S(49) => 
                           P_tmp_2_49_port, S(48) => P_tmp_2_48_port, S(47) => 
                           P_tmp_2_47_port, S(46) => P_tmp_2_46_port, S(45) => 
                           P_tmp_2_45_port, S(44) => P_tmp_2_44_port, S(43) => 
                           P_tmp_2_43_port, S(42) => P_tmp_2_42_port, S(41) => 
                           P_tmp_2_41_port, S(40) => P_tmp_2_40_port, S(39) => 
                           P_tmp_2_39_port, S(38) => P_tmp_2_38_port, S(37) => 
                           P_tmp_2_37_port, S(36) => P_tmp_2_36_port, S(35) => 
                           P_tmp_2_35_port, S(34) => P_tmp_2_34_port, S(33) => 
                           P_tmp_2_33_port, S(32) => P_tmp_2_32_port, S(31) => 
                           P_tmp_2_31_port, S(30) => P_tmp_2_30_port, S(29) => 
                           P_tmp_2_29_port, S(28) => P_tmp_2_28_port, S(27) => 
                           P_tmp_2_27_port, S(26) => P_tmp_2_26_port, S(25) => 
                           P_tmp_2_25_port, S(24) => P_tmp_2_24_port, S(23) => 
                           P_tmp_2_23_port, S(22) => P_tmp_2_22_port, S(21) => 
                           P_tmp_2_21_port, S(20) => P_tmp_2_20_port, S(19) => 
                           P_tmp_2_19_port, S(18) => P_tmp_2_18_port, S(17) => 
                           P_tmp_2_17_port, S(16) => P_tmp_2_16_port, S(15) => 
                           P_tmp_2_15_port, S(14) => P_tmp_2_14_port, S(13) => 
                           P_tmp_2_13_port, S(12) => P_tmp_2_12_port, S(11) => 
                           P_tmp_2_11_port, S(10) => P_tmp_2_10_port, S(9) => 
                           P_tmp_2_9_port, S(8) => P_tmp_2_8_port, S(7) => 
                           P_tmp_2_7_port, S(6) => P_tmp_2_6_port, S(5) => 
                           P_tmp_2_5_port, S(4) => P_tmp_2_4_port, S(3) => 
                           P_tmp_2_3_port, S(2) => P_tmp_2_2_port, S(1) => 
                           P_tmp_2_1_port, S(0) => P_tmp_2_0_port, Co => n_1281
                           );
   RCAi_2 : RCA_NBIT64_13 port map( A(63) => P_tmp_2_63_port, A(62) => 
                           P_tmp_2_62_port, A(61) => P_tmp_2_61_port, A(60) => 
                           P_tmp_2_60_port, A(59) => P_tmp_2_59_port, A(58) => 
                           P_tmp_2_58_port, A(57) => P_tmp_2_57_port, A(56) => 
                           P_tmp_2_56_port, A(55) => P_tmp_2_55_port, A(54) => 
                           P_tmp_2_54_port, A(53) => P_tmp_2_53_port, A(52) => 
                           P_tmp_2_52_port, A(51) => P_tmp_2_51_port, A(50) => 
                           P_tmp_2_50_port, A(49) => P_tmp_2_49_port, A(48) => 
                           P_tmp_2_48_port, A(47) => P_tmp_2_47_port, A(46) => 
                           P_tmp_2_46_port, A(45) => P_tmp_2_45_port, A(44) => 
                           P_tmp_2_44_port, A(43) => P_tmp_2_43_port, A(42) => 
                           P_tmp_2_42_port, A(41) => P_tmp_2_41_port, A(40) => 
                           P_tmp_2_40_port, A(39) => P_tmp_2_39_port, A(38) => 
                           P_tmp_2_38_port, A(37) => P_tmp_2_37_port, A(36) => 
                           P_tmp_2_36_port, A(35) => P_tmp_2_35_port, A(34) => 
                           P_tmp_2_34_port, A(33) => P_tmp_2_33_port, A(32) => 
                           P_tmp_2_32_port, A(31) => P_tmp_2_31_port, A(30) => 
                           P_tmp_2_30_port, A(29) => P_tmp_2_29_port, A(28) => 
                           P_tmp_2_28_port, A(27) => P_tmp_2_27_port, A(26) => 
                           P_tmp_2_26_port, A(25) => P_tmp_2_25_port, A(24) => 
                           P_tmp_2_24_port, A(23) => P_tmp_2_23_port, A(22) => 
                           P_tmp_2_22_port, A(21) => P_tmp_2_21_port, A(20) => 
                           P_tmp_2_20_port, A(19) => P_tmp_2_19_port, A(18) => 
                           P_tmp_2_18_port, A(17) => P_tmp_2_17_port, A(16) => 
                           P_tmp_2_16_port, A(15) => P_tmp_2_15_port, A(14) => 
                           P_tmp_2_14_port, A(13) => P_tmp_2_13_port, A(12) => 
                           P_tmp_2_12_port, A(11) => P_tmp_2_11_port, A(10) => 
                           P_tmp_2_10_port, A(9) => P_tmp_2_9_port, A(8) => 
                           P_tmp_2_8_port, A(7) => P_tmp_2_7_port, A(6) => 
                           P_tmp_2_6_port, A(5) => P_tmp_2_5_port, A(4) => 
                           P_tmp_2_4_port, A(3) => P_tmp_2_3_port, A(2) => 
                           P_tmp_2_2_port, A(1) => P_tmp_2_1_port, A(0) => 
                           P_tmp_2_0_port, B(63) => OUT_MUX_3_63_port, B(62) =>
                           OUT_MUX_3_62_port, B(61) => OUT_MUX_3_61_port, B(60)
                           => OUT_MUX_3_60_port, B(59) => OUT_MUX_3_59_port, 
                           B(58) => OUT_MUX_3_58_port, B(57) => 
                           OUT_MUX_3_57_port, B(56) => OUT_MUX_3_56_port, B(55)
                           => OUT_MUX_3_55_port, B(54) => OUT_MUX_3_54_port, 
                           B(53) => OUT_MUX_3_53_port, B(52) => 
                           OUT_MUX_3_52_port, B(51) => OUT_MUX_3_51_port, B(50)
                           => OUT_MUX_3_50_port, B(49) => OUT_MUX_3_49_port, 
                           B(48) => OUT_MUX_3_48_port, B(47) => 
                           OUT_MUX_3_47_port, B(46) => OUT_MUX_3_46_port, B(45)
                           => OUT_MUX_3_45_port, B(44) => OUT_MUX_3_44_port, 
                           B(43) => OUT_MUX_3_43_port, B(42) => 
                           OUT_MUX_3_42_port, B(41) => OUT_MUX_3_41_port, B(40)
                           => OUT_MUX_3_40_port, B(39) => OUT_MUX_3_39_port, 
                           B(38) => OUT_MUX_3_38_port, B(37) => 
                           OUT_MUX_3_37_port, B(36) => OUT_MUX_3_36_port, B(35)
                           => OUT_MUX_3_35_port, B(34) => OUT_MUX_3_34_port, 
                           B(33) => OUT_MUX_3_33_port, B(32) => 
                           OUT_MUX_3_32_port, B(31) => OUT_MUX_3_31_port, B(30)
                           => OUT_MUX_3_30_port, B(29) => OUT_MUX_3_29_port, 
                           B(28) => OUT_MUX_3_28_port, B(27) => 
                           OUT_MUX_3_27_port, B(26) => OUT_MUX_3_26_port, B(25)
                           => OUT_MUX_3_25_port, B(24) => OUT_MUX_3_24_port, 
                           B(23) => OUT_MUX_3_23_port, B(22) => 
                           OUT_MUX_3_22_port, B(21) => OUT_MUX_3_21_port, B(20)
                           => OUT_MUX_3_20_port, B(19) => OUT_MUX_3_19_port, 
                           B(18) => OUT_MUX_3_18_port, B(17) => 
                           OUT_MUX_3_17_port, B(16) => OUT_MUX_3_16_port, B(15)
                           => OUT_MUX_3_15_port, B(14) => OUT_MUX_3_14_port, 
                           B(13) => OUT_MUX_3_13_port, B(12) => 
                           OUT_MUX_3_12_port, B(11) => OUT_MUX_3_11_port, B(10)
                           => OUT_MUX_3_10_port, B(9) => OUT_MUX_3_9_port, B(8)
                           => OUT_MUX_3_8_port, B(7) => OUT_MUX_3_7_port, B(6) 
                           => OUT_MUX_3_6_port, B(5) => OUT_MUX_3_5_port, B(4) 
                           => OUT_MUX_3_4_port, B(3) => OUT_MUX_3_3_port, B(2) 
                           => OUT_MUX_3_2_port, B(1) => OUT_MUX_3_1_port, B(0) 
                           => OUT_MUX_3_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_3_63_port, S(62) => P_tmp_3_62_port, S(61) => 
                           P_tmp_3_61_port, S(60) => P_tmp_3_60_port, S(59) => 
                           P_tmp_3_59_port, S(58) => P_tmp_3_58_port, S(57) => 
                           P_tmp_3_57_port, S(56) => P_tmp_3_56_port, S(55) => 
                           P_tmp_3_55_port, S(54) => P_tmp_3_54_port, S(53) => 
                           P_tmp_3_53_port, S(52) => P_tmp_3_52_port, S(51) => 
                           P_tmp_3_51_port, S(50) => P_tmp_3_50_port, S(49) => 
                           P_tmp_3_49_port, S(48) => P_tmp_3_48_port, S(47) => 
                           P_tmp_3_47_port, S(46) => P_tmp_3_46_port, S(45) => 
                           P_tmp_3_45_port, S(44) => P_tmp_3_44_port, S(43) => 
                           P_tmp_3_43_port, S(42) => P_tmp_3_42_port, S(41) => 
                           P_tmp_3_41_port, S(40) => P_tmp_3_40_port, S(39) => 
                           P_tmp_3_39_port, S(38) => P_tmp_3_38_port, S(37) => 
                           P_tmp_3_37_port, S(36) => P_tmp_3_36_port, S(35) => 
                           P_tmp_3_35_port, S(34) => P_tmp_3_34_port, S(33) => 
                           P_tmp_3_33_port, S(32) => P_tmp_3_32_port, S(31) => 
                           P_tmp_3_31_port, S(30) => P_tmp_3_30_port, S(29) => 
                           P_tmp_3_29_port, S(28) => P_tmp_3_28_port, S(27) => 
                           P_tmp_3_27_port, S(26) => P_tmp_3_26_port, S(25) => 
                           P_tmp_3_25_port, S(24) => P_tmp_3_24_port, S(23) => 
                           P_tmp_3_23_port, S(22) => P_tmp_3_22_port, S(21) => 
                           P_tmp_3_21_port, S(20) => P_tmp_3_20_port, S(19) => 
                           P_tmp_3_19_port, S(18) => P_tmp_3_18_port, S(17) => 
                           P_tmp_3_17_port, S(16) => P_tmp_3_16_port, S(15) => 
                           P_tmp_3_15_port, S(14) => P_tmp_3_14_port, S(13) => 
                           P_tmp_3_13_port, S(12) => P_tmp_3_12_port, S(11) => 
                           P_tmp_3_11_port, S(10) => P_tmp_3_10_port, S(9) => 
                           P_tmp_3_9_port, S(8) => P_tmp_3_8_port, S(7) => 
                           P_tmp_3_7_port, S(6) => P_tmp_3_6_port, S(5) => 
                           P_tmp_3_5_port, S(4) => P_tmp_3_4_port, S(3) => 
                           P_tmp_3_3_port, S(2) => P_tmp_3_2_port, S(1) => 
                           P_tmp_3_1_port, S(0) => P_tmp_3_0_port, Co => n_1282
                           );
   RCAi_3 : RCA_NBIT64_12 port map( A(63) => P_tmp_3_63_port, A(62) => 
                           P_tmp_3_62_port, A(61) => P_tmp_3_61_port, A(60) => 
                           P_tmp_3_60_port, A(59) => P_tmp_3_59_port, A(58) => 
                           P_tmp_3_58_port, A(57) => P_tmp_3_57_port, A(56) => 
                           P_tmp_3_56_port, A(55) => P_tmp_3_55_port, A(54) => 
                           P_tmp_3_54_port, A(53) => P_tmp_3_53_port, A(52) => 
                           P_tmp_3_52_port, A(51) => P_tmp_3_51_port, A(50) => 
                           P_tmp_3_50_port, A(49) => P_tmp_3_49_port, A(48) => 
                           P_tmp_3_48_port, A(47) => P_tmp_3_47_port, A(46) => 
                           P_tmp_3_46_port, A(45) => P_tmp_3_45_port, A(44) => 
                           P_tmp_3_44_port, A(43) => P_tmp_3_43_port, A(42) => 
                           P_tmp_3_42_port, A(41) => P_tmp_3_41_port, A(40) => 
                           P_tmp_3_40_port, A(39) => P_tmp_3_39_port, A(38) => 
                           P_tmp_3_38_port, A(37) => P_tmp_3_37_port, A(36) => 
                           P_tmp_3_36_port, A(35) => P_tmp_3_35_port, A(34) => 
                           P_tmp_3_34_port, A(33) => P_tmp_3_33_port, A(32) => 
                           P_tmp_3_32_port, A(31) => P_tmp_3_31_port, A(30) => 
                           P_tmp_3_30_port, A(29) => P_tmp_3_29_port, A(28) => 
                           P_tmp_3_28_port, A(27) => P_tmp_3_27_port, A(26) => 
                           P_tmp_3_26_port, A(25) => P_tmp_3_25_port, A(24) => 
                           P_tmp_3_24_port, A(23) => P_tmp_3_23_port, A(22) => 
                           P_tmp_3_22_port, A(21) => P_tmp_3_21_port, A(20) => 
                           P_tmp_3_20_port, A(19) => P_tmp_3_19_port, A(18) => 
                           P_tmp_3_18_port, A(17) => P_tmp_3_17_port, A(16) => 
                           P_tmp_3_16_port, A(15) => P_tmp_3_15_port, A(14) => 
                           P_tmp_3_14_port, A(13) => P_tmp_3_13_port, A(12) => 
                           P_tmp_3_12_port, A(11) => P_tmp_3_11_port, A(10) => 
                           P_tmp_3_10_port, A(9) => P_tmp_3_9_port, A(8) => 
                           P_tmp_3_8_port, A(7) => P_tmp_3_7_port, A(6) => 
                           P_tmp_3_6_port, A(5) => P_tmp_3_5_port, A(4) => 
                           P_tmp_3_4_port, A(3) => P_tmp_3_3_port, A(2) => 
                           P_tmp_3_2_port, A(1) => P_tmp_3_1_port, A(0) => 
                           P_tmp_3_0_port, B(63) => OUT_MUX_4_63_port, B(62) =>
                           OUT_MUX_4_62_port, B(61) => OUT_MUX_4_61_port, B(60)
                           => OUT_MUX_4_60_port, B(59) => OUT_MUX_4_59_port, 
                           B(58) => OUT_MUX_4_58_port, B(57) => 
                           OUT_MUX_4_57_port, B(56) => OUT_MUX_4_56_port, B(55)
                           => OUT_MUX_4_55_port, B(54) => OUT_MUX_4_54_port, 
                           B(53) => OUT_MUX_4_53_port, B(52) => 
                           OUT_MUX_4_52_port, B(51) => OUT_MUX_4_51_port, B(50)
                           => OUT_MUX_4_50_port, B(49) => OUT_MUX_4_49_port, 
                           B(48) => OUT_MUX_4_48_port, B(47) => 
                           OUT_MUX_4_47_port, B(46) => OUT_MUX_4_46_port, B(45)
                           => OUT_MUX_4_45_port, B(44) => OUT_MUX_4_44_port, 
                           B(43) => OUT_MUX_4_43_port, B(42) => 
                           OUT_MUX_4_42_port, B(41) => OUT_MUX_4_41_port, B(40)
                           => OUT_MUX_4_40_port, B(39) => OUT_MUX_4_39_port, 
                           B(38) => OUT_MUX_4_38_port, B(37) => 
                           OUT_MUX_4_37_port, B(36) => OUT_MUX_4_36_port, B(35)
                           => OUT_MUX_4_35_port, B(34) => OUT_MUX_4_34_port, 
                           B(33) => OUT_MUX_4_33_port, B(32) => 
                           OUT_MUX_4_32_port, B(31) => OUT_MUX_4_31_port, B(30)
                           => OUT_MUX_4_30_port, B(29) => OUT_MUX_4_29_port, 
                           B(28) => OUT_MUX_4_28_port, B(27) => 
                           OUT_MUX_4_27_port, B(26) => OUT_MUX_4_26_port, B(25)
                           => OUT_MUX_4_25_port, B(24) => OUT_MUX_4_24_port, 
                           B(23) => OUT_MUX_4_23_port, B(22) => 
                           OUT_MUX_4_22_port, B(21) => OUT_MUX_4_21_port, B(20)
                           => OUT_MUX_4_20_port, B(19) => OUT_MUX_4_19_port, 
                           B(18) => OUT_MUX_4_18_port, B(17) => 
                           OUT_MUX_4_17_port, B(16) => OUT_MUX_4_16_port, B(15)
                           => OUT_MUX_4_15_port, B(14) => OUT_MUX_4_14_port, 
                           B(13) => OUT_MUX_4_13_port, B(12) => 
                           OUT_MUX_4_12_port, B(11) => OUT_MUX_4_11_port, B(10)
                           => OUT_MUX_4_10_port, B(9) => OUT_MUX_4_9_port, B(8)
                           => OUT_MUX_4_8_port, B(7) => OUT_MUX_4_7_port, B(6) 
                           => OUT_MUX_4_6_port, B(5) => OUT_MUX_4_5_port, B(4) 
                           => OUT_MUX_4_4_port, B(3) => OUT_MUX_4_3_port, B(2) 
                           => OUT_MUX_4_2_port, B(1) => OUT_MUX_4_1_port, B(0) 
                           => OUT_MUX_4_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_4_63_port, S(62) => P_tmp_4_62_port, S(61) => 
                           P_tmp_4_61_port, S(60) => P_tmp_4_60_port, S(59) => 
                           P_tmp_4_59_port, S(58) => P_tmp_4_58_port, S(57) => 
                           P_tmp_4_57_port, S(56) => P_tmp_4_56_port, S(55) => 
                           P_tmp_4_55_port, S(54) => P_tmp_4_54_port, S(53) => 
                           P_tmp_4_53_port, S(52) => P_tmp_4_52_port, S(51) => 
                           P_tmp_4_51_port, S(50) => P_tmp_4_50_port, S(49) => 
                           P_tmp_4_49_port, S(48) => P_tmp_4_48_port, S(47) => 
                           P_tmp_4_47_port, S(46) => P_tmp_4_46_port, S(45) => 
                           P_tmp_4_45_port, S(44) => P_tmp_4_44_port, S(43) => 
                           P_tmp_4_43_port, S(42) => P_tmp_4_42_port, S(41) => 
                           P_tmp_4_41_port, S(40) => P_tmp_4_40_port, S(39) => 
                           P_tmp_4_39_port, S(38) => P_tmp_4_38_port, S(37) => 
                           P_tmp_4_37_port, S(36) => P_tmp_4_36_port, S(35) => 
                           P_tmp_4_35_port, S(34) => P_tmp_4_34_port, S(33) => 
                           P_tmp_4_33_port, S(32) => P_tmp_4_32_port, S(31) => 
                           P_tmp_4_31_port, S(30) => P_tmp_4_30_port, S(29) => 
                           P_tmp_4_29_port, S(28) => P_tmp_4_28_port, S(27) => 
                           P_tmp_4_27_port, S(26) => P_tmp_4_26_port, S(25) => 
                           P_tmp_4_25_port, S(24) => P_tmp_4_24_port, S(23) => 
                           P_tmp_4_23_port, S(22) => P_tmp_4_22_port, S(21) => 
                           P_tmp_4_21_port, S(20) => P_tmp_4_20_port, S(19) => 
                           P_tmp_4_19_port, S(18) => P_tmp_4_18_port, S(17) => 
                           P_tmp_4_17_port, S(16) => P_tmp_4_16_port, S(15) => 
                           P_tmp_4_15_port, S(14) => P_tmp_4_14_port, S(13) => 
                           P_tmp_4_13_port, S(12) => P_tmp_4_12_port, S(11) => 
                           P_tmp_4_11_port, S(10) => P_tmp_4_10_port, S(9) => 
                           P_tmp_4_9_port, S(8) => P_tmp_4_8_port, S(7) => 
                           P_tmp_4_7_port, S(6) => P_tmp_4_6_port, S(5) => 
                           P_tmp_4_5_port, S(4) => P_tmp_4_4_port, S(3) => 
                           P_tmp_4_3_port, S(2) => P_tmp_4_2_port, S(1) => 
                           P_tmp_4_1_port, S(0) => P_tmp_4_0_port, Co => n_1283
                           );
   RCAi_4 : RCA_NBIT64_11 port map( A(63) => P_tmp_4_63_port, A(62) => 
                           P_tmp_4_62_port, A(61) => P_tmp_4_61_port, A(60) => 
                           P_tmp_4_60_port, A(59) => P_tmp_4_59_port, A(58) => 
                           P_tmp_4_58_port, A(57) => P_tmp_4_57_port, A(56) => 
                           P_tmp_4_56_port, A(55) => P_tmp_4_55_port, A(54) => 
                           P_tmp_4_54_port, A(53) => P_tmp_4_53_port, A(52) => 
                           P_tmp_4_52_port, A(51) => P_tmp_4_51_port, A(50) => 
                           P_tmp_4_50_port, A(49) => P_tmp_4_49_port, A(48) => 
                           P_tmp_4_48_port, A(47) => P_tmp_4_47_port, A(46) => 
                           P_tmp_4_46_port, A(45) => P_tmp_4_45_port, A(44) => 
                           P_tmp_4_44_port, A(43) => P_tmp_4_43_port, A(42) => 
                           P_tmp_4_42_port, A(41) => P_tmp_4_41_port, A(40) => 
                           P_tmp_4_40_port, A(39) => P_tmp_4_39_port, A(38) => 
                           P_tmp_4_38_port, A(37) => P_tmp_4_37_port, A(36) => 
                           P_tmp_4_36_port, A(35) => P_tmp_4_35_port, A(34) => 
                           P_tmp_4_34_port, A(33) => P_tmp_4_33_port, A(32) => 
                           P_tmp_4_32_port, A(31) => P_tmp_4_31_port, A(30) => 
                           P_tmp_4_30_port, A(29) => P_tmp_4_29_port, A(28) => 
                           P_tmp_4_28_port, A(27) => P_tmp_4_27_port, A(26) => 
                           P_tmp_4_26_port, A(25) => P_tmp_4_25_port, A(24) => 
                           P_tmp_4_24_port, A(23) => P_tmp_4_23_port, A(22) => 
                           P_tmp_4_22_port, A(21) => P_tmp_4_21_port, A(20) => 
                           P_tmp_4_20_port, A(19) => P_tmp_4_19_port, A(18) => 
                           P_tmp_4_18_port, A(17) => P_tmp_4_17_port, A(16) => 
                           P_tmp_4_16_port, A(15) => P_tmp_4_15_port, A(14) => 
                           P_tmp_4_14_port, A(13) => P_tmp_4_13_port, A(12) => 
                           P_tmp_4_12_port, A(11) => P_tmp_4_11_port, A(10) => 
                           P_tmp_4_10_port, A(9) => P_tmp_4_9_port, A(8) => 
                           P_tmp_4_8_port, A(7) => P_tmp_4_7_port, A(6) => 
                           P_tmp_4_6_port, A(5) => P_tmp_4_5_port, A(4) => 
                           P_tmp_4_4_port, A(3) => P_tmp_4_3_port, A(2) => 
                           P_tmp_4_2_port, A(1) => P_tmp_4_1_port, A(0) => 
                           P_tmp_4_0_port, B(63) => OUT_MUX_5_63_port, B(62) =>
                           OUT_MUX_5_62_port, B(61) => OUT_MUX_5_61_port, B(60)
                           => OUT_MUX_5_60_port, B(59) => OUT_MUX_5_59_port, 
                           B(58) => OUT_MUX_5_58_port, B(57) => 
                           OUT_MUX_5_57_port, B(56) => OUT_MUX_5_56_port, B(55)
                           => OUT_MUX_5_55_port, B(54) => OUT_MUX_5_54_port, 
                           B(53) => OUT_MUX_5_53_port, B(52) => 
                           OUT_MUX_5_52_port, B(51) => OUT_MUX_5_51_port, B(50)
                           => OUT_MUX_5_50_port, B(49) => OUT_MUX_5_49_port, 
                           B(48) => OUT_MUX_5_48_port, B(47) => 
                           OUT_MUX_5_47_port, B(46) => OUT_MUX_5_46_port, B(45)
                           => OUT_MUX_5_45_port, B(44) => OUT_MUX_5_44_port, 
                           B(43) => OUT_MUX_5_43_port, B(42) => 
                           OUT_MUX_5_42_port, B(41) => OUT_MUX_5_41_port, B(40)
                           => OUT_MUX_5_40_port, B(39) => OUT_MUX_5_39_port, 
                           B(38) => OUT_MUX_5_38_port, B(37) => 
                           OUT_MUX_5_37_port, B(36) => OUT_MUX_5_36_port, B(35)
                           => OUT_MUX_5_35_port, B(34) => OUT_MUX_5_34_port, 
                           B(33) => OUT_MUX_5_33_port, B(32) => 
                           OUT_MUX_5_32_port, B(31) => OUT_MUX_5_31_port, B(30)
                           => OUT_MUX_5_30_port, B(29) => OUT_MUX_5_29_port, 
                           B(28) => OUT_MUX_5_28_port, B(27) => 
                           OUT_MUX_5_27_port, B(26) => OUT_MUX_5_26_port, B(25)
                           => OUT_MUX_5_25_port, B(24) => OUT_MUX_5_24_port, 
                           B(23) => OUT_MUX_5_23_port, B(22) => 
                           OUT_MUX_5_22_port, B(21) => OUT_MUX_5_21_port, B(20)
                           => OUT_MUX_5_20_port, B(19) => OUT_MUX_5_19_port, 
                           B(18) => OUT_MUX_5_18_port, B(17) => 
                           OUT_MUX_5_17_port, B(16) => OUT_MUX_5_16_port, B(15)
                           => OUT_MUX_5_15_port, B(14) => OUT_MUX_5_14_port, 
                           B(13) => OUT_MUX_5_13_port, B(12) => 
                           OUT_MUX_5_12_port, B(11) => OUT_MUX_5_11_port, B(10)
                           => OUT_MUX_5_10_port, B(9) => OUT_MUX_5_9_port, B(8)
                           => OUT_MUX_5_8_port, B(7) => OUT_MUX_5_7_port, B(6) 
                           => OUT_MUX_5_6_port, B(5) => OUT_MUX_5_5_port, B(4) 
                           => OUT_MUX_5_4_port, B(3) => OUT_MUX_5_3_port, B(2) 
                           => OUT_MUX_5_2_port, B(1) => OUT_MUX_5_1_port, B(0) 
                           => OUT_MUX_5_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_5_63_port, S(62) => P_tmp_5_62_port, S(61) => 
                           P_tmp_5_61_port, S(60) => P_tmp_5_60_port, S(59) => 
                           P_tmp_5_59_port, S(58) => P_tmp_5_58_port, S(57) => 
                           P_tmp_5_57_port, S(56) => P_tmp_5_56_port, S(55) => 
                           P_tmp_5_55_port, S(54) => P_tmp_5_54_port, S(53) => 
                           P_tmp_5_53_port, S(52) => P_tmp_5_52_port, S(51) => 
                           P_tmp_5_51_port, S(50) => P_tmp_5_50_port, S(49) => 
                           P_tmp_5_49_port, S(48) => P_tmp_5_48_port, S(47) => 
                           P_tmp_5_47_port, S(46) => P_tmp_5_46_port, S(45) => 
                           P_tmp_5_45_port, S(44) => P_tmp_5_44_port, S(43) => 
                           P_tmp_5_43_port, S(42) => P_tmp_5_42_port, S(41) => 
                           P_tmp_5_41_port, S(40) => P_tmp_5_40_port, S(39) => 
                           P_tmp_5_39_port, S(38) => P_tmp_5_38_port, S(37) => 
                           P_tmp_5_37_port, S(36) => P_tmp_5_36_port, S(35) => 
                           P_tmp_5_35_port, S(34) => P_tmp_5_34_port, S(33) => 
                           P_tmp_5_33_port, S(32) => P_tmp_5_32_port, S(31) => 
                           P_tmp_5_31_port, S(30) => P_tmp_5_30_port, S(29) => 
                           P_tmp_5_29_port, S(28) => P_tmp_5_28_port, S(27) => 
                           P_tmp_5_27_port, S(26) => P_tmp_5_26_port, S(25) => 
                           P_tmp_5_25_port, S(24) => P_tmp_5_24_port, S(23) => 
                           P_tmp_5_23_port, S(22) => P_tmp_5_22_port, S(21) => 
                           P_tmp_5_21_port, S(20) => P_tmp_5_20_port, S(19) => 
                           P_tmp_5_19_port, S(18) => P_tmp_5_18_port, S(17) => 
                           P_tmp_5_17_port, S(16) => P_tmp_5_16_port, S(15) => 
                           P_tmp_5_15_port, S(14) => P_tmp_5_14_port, S(13) => 
                           P_tmp_5_13_port, S(12) => P_tmp_5_12_port, S(11) => 
                           P_tmp_5_11_port, S(10) => P_tmp_5_10_port, S(9) => 
                           P_tmp_5_9_port, S(8) => P_tmp_5_8_port, S(7) => 
                           P_tmp_5_7_port, S(6) => P_tmp_5_6_port, S(5) => 
                           P_tmp_5_5_port, S(4) => P_tmp_5_4_port, S(3) => 
                           P_tmp_5_3_port, S(2) => P_tmp_5_2_port, S(1) => 
                           P_tmp_5_1_port, S(0) => P_tmp_5_0_port, Co => n_1284
                           );
   RCAi_5 : RCA_NBIT64_10 port map( A(63) => P_tmp_5_63_port, A(62) => 
                           P_tmp_5_62_port, A(61) => P_tmp_5_61_port, A(60) => 
                           P_tmp_5_60_port, A(59) => P_tmp_5_59_port, A(58) => 
                           P_tmp_5_58_port, A(57) => P_tmp_5_57_port, A(56) => 
                           P_tmp_5_56_port, A(55) => P_tmp_5_55_port, A(54) => 
                           P_tmp_5_54_port, A(53) => P_tmp_5_53_port, A(52) => 
                           P_tmp_5_52_port, A(51) => P_tmp_5_51_port, A(50) => 
                           P_tmp_5_50_port, A(49) => P_tmp_5_49_port, A(48) => 
                           P_tmp_5_48_port, A(47) => P_tmp_5_47_port, A(46) => 
                           P_tmp_5_46_port, A(45) => P_tmp_5_45_port, A(44) => 
                           P_tmp_5_44_port, A(43) => P_tmp_5_43_port, A(42) => 
                           P_tmp_5_42_port, A(41) => P_tmp_5_41_port, A(40) => 
                           P_tmp_5_40_port, A(39) => P_tmp_5_39_port, A(38) => 
                           P_tmp_5_38_port, A(37) => P_tmp_5_37_port, A(36) => 
                           P_tmp_5_36_port, A(35) => P_tmp_5_35_port, A(34) => 
                           P_tmp_5_34_port, A(33) => P_tmp_5_33_port, A(32) => 
                           P_tmp_5_32_port, A(31) => P_tmp_5_31_port, A(30) => 
                           P_tmp_5_30_port, A(29) => P_tmp_5_29_port, A(28) => 
                           P_tmp_5_28_port, A(27) => P_tmp_5_27_port, A(26) => 
                           P_tmp_5_26_port, A(25) => P_tmp_5_25_port, A(24) => 
                           P_tmp_5_24_port, A(23) => P_tmp_5_23_port, A(22) => 
                           P_tmp_5_22_port, A(21) => P_tmp_5_21_port, A(20) => 
                           P_tmp_5_20_port, A(19) => P_tmp_5_19_port, A(18) => 
                           P_tmp_5_18_port, A(17) => P_tmp_5_17_port, A(16) => 
                           P_tmp_5_16_port, A(15) => P_tmp_5_15_port, A(14) => 
                           P_tmp_5_14_port, A(13) => P_tmp_5_13_port, A(12) => 
                           P_tmp_5_12_port, A(11) => P_tmp_5_11_port, A(10) => 
                           P_tmp_5_10_port, A(9) => P_tmp_5_9_port, A(8) => 
                           P_tmp_5_8_port, A(7) => P_tmp_5_7_port, A(6) => 
                           P_tmp_5_6_port, A(5) => P_tmp_5_5_port, A(4) => 
                           P_tmp_5_4_port, A(3) => P_tmp_5_3_port, A(2) => 
                           P_tmp_5_2_port, A(1) => P_tmp_5_1_port, A(0) => 
                           P_tmp_5_0_port, B(63) => OUT_MUX_6_63_port, B(62) =>
                           OUT_MUX_6_62_port, B(61) => OUT_MUX_6_61_port, B(60)
                           => OUT_MUX_6_60_port, B(59) => OUT_MUX_6_59_port, 
                           B(58) => OUT_MUX_6_58_port, B(57) => 
                           OUT_MUX_6_57_port, B(56) => OUT_MUX_6_56_port, B(55)
                           => OUT_MUX_6_55_port, B(54) => OUT_MUX_6_54_port, 
                           B(53) => OUT_MUX_6_53_port, B(52) => 
                           OUT_MUX_6_52_port, B(51) => OUT_MUX_6_51_port, B(50)
                           => OUT_MUX_6_50_port, B(49) => OUT_MUX_6_49_port, 
                           B(48) => OUT_MUX_6_48_port, B(47) => 
                           OUT_MUX_6_47_port, B(46) => OUT_MUX_6_46_port, B(45)
                           => OUT_MUX_6_45_port, B(44) => OUT_MUX_6_44_port, 
                           B(43) => OUT_MUX_6_43_port, B(42) => 
                           OUT_MUX_6_42_port, B(41) => OUT_MUX_6_41_port, B(40)
                           => OUT_MUX_6_40_port, B(39) => OUT_MUX_6_39_port, 
                           B(38) => OUT_MUX_6_38_port, B(37) => 
                           OUT_MUX_6_37_port, B(36) => OUT_MUX_6_36_port, B(35)
                           => OUT_MUX_6_35_port, B(34) => OUT_MUX_6_34_port, 
                           B(33) => OUT_MUX_6_33_port, B(32) => 
                           OUT_MUX_6_32_port, B(31) => OUT_MUX_6_31_port, B(30)
                           => OUT_MUX_6_30_port, B(29) => OUT_MUX_6_29_port, 
                           B(28) => OUT_MUX_6_28_port, B(27) => 
                           OUT_MUX_6_27_port, B(26) => OUT_MUX_6_26_port, B(25)
                           => OUT_MUX_6_25_port, B(24) => OUT_MUX_6_24_port, 
                           B(23) => OUT_MUX_6_23_port, B(22) => 
                           OUT_MUX_6_22_port, B(21) => OUT_MUX_6_21_port, B(20)
                           => OUT_MUX_6_20_port, B(19) => OUT_MUX_6_19_port, 
                           B(18) => OUT_MUX_6_18_port, B(17) => 
                           OUT_MUX_6_17_port, B(16) => OUT_MUX_6_16_port, B(15)
                           => OUT_MUX_6_15_port, B(14) => OUT_MUX_6_14_port, 
                           B(13) => OUT_MUX_6_13_port, B(12) => 
                           OUT_MUX_6_12_port, B(11) => OUT_MUX_6_11_port, B(10)
                           => OUT_MUX_6_10_port, B(9) => OUT_MUX_6_9_port, B(8)
                           => OUT_MUX_6_8_port, B(7) => OUT_MUX_6_7_port, B(6) 
                           => OUT_MUX_6_6_port, B(5) => OUT_MUX_6_5_port, B(4) 
                           => OUT_MUX_6_4_port, B(3) => OUT_MUX_6_3_port, B(2) 
                           => OUT_MUX_6_2_port, B(1) => OUT_MUX_6_1_port, B(0) 
                           => OUT_MUX_6_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_6_63_port, S(62) => P_tmp_6_62_port, S(61) => 
                           P_tmp_6_61_port, S(60) => P_tmp_6_60_port, S(59) => 
                           P_tmp_6_59_port, S(58) => P_tmp_6_58_port, S(57) => 
                           P_tmp_6_57_port, S(56) => P_tmp_6_56_port, S(55) => 
                           P_tmp_6_55_port, S(54) => P_tmp_6_54_port, S(53) => 
                           P_tmp_6_53_port, S(52) => P_tmp_6_52_port, S(51) => 
                           P_tmp_6_51_port, S(50) => P_tmp_6_50_port, S(49) => 
                           P_tmp_6_49_port, S(48) => P_tmp_6_48_port, S(47) => 
                           P_tmp_6_47_port, S(46) => P_tmp_6_46_port, S(45) => 
                           P_tmp_6_45_port, S(44) => P_tmp_6_44_port, S(43) => 
                           P_tmp_6_43_port, S(42) => P_tmp_6_42_port, S(41) => 
                           P_tmp_6_41_port, S(40) => P_tmp_6_40_port, S(39) => 
                           P_tmp_6_39_port, S(38) => P_tmp_6_38_port, S(37) => 
                           P_tmp_6_37_port, S(36) => P_tmp_6_36_port, S(35) => 
                           P_tmp_6_35_port, S(34) => P_tmp_6_34_port, S(33) => 
                           P_tmp_6_33_port, S(32) => P_tmp_6_32_port, S(31) => 
                           P_tmp_6_31_port, S(30) => P_tmp_6_30_port, S(29) => 
                           P_tmp_6_29_port, S(28) => P_tmp_6_28_port, S(27) => 
                           P_tmp_6_27_port, S(26) => P_tmp_6_26_port, S(25) => 
                           P_tmp_6_25_port, S(24) => P_tmp_6_24_port, S(23) => 
                           P_tmp_6_23_port, S(22) => P_tmp_6_22_port, S(21) => 
                           P_tmp_6_21_port, S(20) => P_tmp_6_20_port, S(19) => 
                           P_tmp_6_19_port, S(18) => P_tmp_6_18_port, S(17) => 
                           P_tmp_6_17_port, S(16) => P_tmp_6_16_port, S(15) => 
                           P_tmp_6_15_port, S(14) => P_tmp_6_14_port, S(13) => 
                           P_tmp_6_13_port, S(12) => P_tmp_6_12_port, S(11) => 
                           P_tmp_6_11_port, S(10) => P_tmp_6_10_port, S(9) => 
                           P_tmp_6_9_port, S(8) => P_tmp_6_8_port, S(7) => 
                           P_tmp_6_7_port, S(6) => P_tmp_6_6_port, S(5) => 
                           P_tmp_6_5_port, S(4) => P_tmp_6_4_port, S(3) => 
                           P_tmp_6_3_port, S(2) => P_tmp_6_2_port, S(1) => 
                           P_tmp_6_1_port, S(0) => P_tmp_6_0_port, Co => n_1285
                           );
   RCAi_6 : RCA_NBIT64_9 port map( A(63) => P_tmp_6_63_port, A(62) => 
                           P_tmp_6_62_port, A(61) => P_tmp_6_61_port, A(60) => 
                           P_tmp_6_60_port, A(59) => P_tmp_6_59_port, A(58) => 
                           P_tmp_6_58_port, A(57) => P_tmp_6_57_port, A(56) => 
                           P_tmp_6_56_port, A(55) => P_tmp_6_55_port, A(54) => 
                           P_tmp_6_54_port, A(53) => P_tmp_6_53_port, A(52) => 
                           P_tmp_6_52_port, A(51) => P_tmp_6_51_port, A(50) => 
                           P_tmp_6_50_port, A(49) => P_tmp_6_49_port, A(48) => 
                           P_tmp_6_48_port, A(47) => P_tmp_6_47_port, A(46) => 
                           P_tmp_6_46_port, A(45) => P_tmp_6_45_port, A(44) => 
                           P_tmp_6_44_port, A(43) => P_tmp_6_43_port, A(42) => 
                           P_tmp_6_42_port, A(41) => P_tmp_6_41_port, A(40) => 
                           P_tmp_6_40_port, A(39) => P_tmp_6_39_port, A(38) => 
                           P_tmp_6_38_port, A(37) => P_tmp_6_37_port, A(36) => 
                           P_tmp_6_36_port, A(35) => P_tmp_6_35_port, A(34) => 
                           P_tmp_6_34_port, A(33) => P_tmp_6_33_port, A(32) => 
                           P_tmp_6_32_port, A(31) => P_tmp_6_31_port, A(30) => 
                           P_tmp_6_30_port, A(29) => P_tmp_6_29_port, A(28) => 
                           P_tmp_6_28_port, A(27) => P_tmp_6_27_port, A(26) => 
                           P_tmp_6_26_port, A(25) => P_tmp_6_25_port, A(24) => 
                           P_tmp_6_24_port, A(23) => P_tmp_6_23_port, A(22) => 
                           P_tmp_6_22_port, A(21) => P_tmp_6_21_port, A(20) => 
                           P_tmp_6_20_port, A(19) => P_tmp_6_19_port, A(18) => 
                           P_tmp_6_18_port, A(17) => P_tmp_6_17_port, A(16) => 
                           P_tmp_6_16_port, A(15) => P_tmp_6_15_port, A(14) => 
                           P_tmp_6_14_port, A(13) => P_tmp_6_13_port, A(12) => 
                           P_tmp_6_12_port, A(11) => P_tmp_6_11_port, A(10) => 
                           P_tmp_6_10_port, A(9) => P_tmp_6_9_port, A(8) => 
                           P_tmp_6_8_port, A(7) => P_tmp_6_7_port, A(6) => 
                           P_tmp_6_6_port, A(5) => P_tmp_6_5_port, A(4) => 
                           P_tmp_6_4_port, A(3) => P_tmp_6_3_port, A(2) => 
                           P_tmp_6_2_port, A(1) => P_tmp_6_1_port, A(0) => 
                           P_tmp_6_0_port, B(63) => OUT_MUX_7_63_port, B(62) =>
                           OUT_MUX_7_62_port, B(61) => OUT_MUX_7_61_port, B(60)
                           => OUT_MUX_7_60_port, B(59) => OUT_MUX_7_59_port, 
                           B(58) => OUT_MUX_7_58_port, B(57) => 
                           OUT_MUX_7_57_port, B(56) => OUT_MUX_7_56_port, B(55)
                           => OUT_MUX_7_55_port, B(54) => OUT_MUX_7_54_port, 
                           B(53) => OUT_MUX_7_53_port, B(52) => 
                           OUT_MUX_7_52_port, B(51) => OUT_MUX_7_51_port, B(50)
                           => OUT_MUX_7_50_port, B(49) => OUT_MUX_7_49_port, 
                           B(48) => OUT_MUX_7_48_port, B(47) => 
                           OUT_MUX_7_47_port, B(46) => OUT_MUX_7_46_port, B(45)
                           => OUT_MUX_7_45_port, B(44) => OUT_MUX_7_44_port, 
                           B(43) => OUT_MUX_7_43_port, B(42) => 
                           OUT_MUX_7_42_port, B(41) => OUT_MUX_7_41_port, B(40)
                           => OUT_MUX_7_40_port, B(39) => OUT_MUX_7_39_port, 
                           B(38) => OUT_MUX_7_38_port, B(37) => 
                           OUT_MUX_7_37_port, B(36) => OUT_MUX_7_36_port, B(35)
                           => OUT_MUX_7_35_port, B(34) => OUT_MUX_7_34_port, 
                           B(33) => OUT_MUX_7_33_port, B(32) => 
                           OUT_MUX_7_32_port, B(31) => OUT_MUX_7_31_port, B(30)
                           => OUT_MUX_7_30_port, B(29) => OUT_MUX_7_29_port, 
                           B(28) => OUT_MUX_7_28_port, B(27) => 
                           OUT_MUX_7_27_port, B(26) => OUT_MUX_7_26_port, B(25)
                           => OUT_MUX_7_25_port, B(24) => OUT_MUX_7_24_port, 
                           B(23) => OUT_MUX_7_23_port, B(22) => 
                           OUT_MUX_7_22_port, B(21) => OUT_MUX_7_21_port, B(20)
                           => OUT_MUX_7_20_port, B(19) => OUT_MUX_7_19_port, 
                           B(18) => OUT_MUX_7_18_port, B(17) => 
                           OUT_MUX_7_17_port, B(16) => OUT_MUX_7_16_port, B(15)
                           => OUT_MUX_7_15_port, B(14) => OUT_MUX_7_14_port, 
                           B(13) => OUT_MUX_7_13_port, B(12) => 
                           OUT_MUX_7_12_port, B(11) => OUT_MUX_7_11_port, B(10)
                           => OUT_MUX_7_10_port, B(9) => OUT_MUX_7_9_port, B(8)
                           => OUT_MUX_7_8_port, B(7) => OUT_MUX_7_7_port, B(6) 
                           => OUT_MUX_7_6_port, B(5) => OUT_MUX_7_5_port, B(4) 
                           => OUT_MUX_7_4_port, B(3) => OUT_MUX_7_3_port, B(2) 
                           => OUT_MUX_7_2_port, B(1) => OUT_MUX_7_1_port, B(0) 
                           => OUT_MUX_7_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_7_63_port, S(62) => P_tmp_7_62_port, S(61) => 
                           P_tmp_7_61_port, S(60) => P_tmp_7_60_port, S(59) => 
                           P_tmp_7_59_port, S(58) => P_tmp_7_58_port, S(57) => 
                           P_tmp_7_57_port, S(56) => P_tmp_7_56_port, S(55) => 
                           P_tmp_7_55_port, S(54) => P_tmp_7_54_port, S(53) => 
                           P_tmp_7_53_port, S(52) => P_tmp_7_52_port, S(51) => 
                           P_tmp_7_51_port, S(50) => P_tmp_7_50_port, S(49) => 
                           P_tmp_7_49_port, S(48) => P_tmp_7_48_port, S(47) => 
                           P_tmp_7_47_port, S(46) => P_tmp_7_46_port, S(45) => 
                           P_tmp_7_45_port, S(44) => P_tmp_7_44_port, S(43) => 
                           P_tmp_7_43_port, S(42) => P_tmp_7_42_port, S(41) => 
                           P_tmp_7_41_port, S(40) => P_tmp_7_40_port, S(39) => 
                           P_tmp_7_39_port, S(38) => P_tmp_7_38_port, S(37) => 
                           P_tmp_7_37_port, S(36) => P_tmp_7_36_port, S(35) => 
                           P_tmp_7_35_port, S(34) => P_tmp_7_34_port, S(33) => 
                           P_tmp_7_33_port, S(32) => P_tmp_7_32_port, S(31) => 
                           P_tmp_7_31_port, S(30) => P_tmp_7_30_port, S(29) => 
                           P_tmp_7_29_port, S(28) => P_tmp_7_28_port, S(27) => 
                           P_tmp_7_27_port, S(26) => P_tmp_7_26_port, S(25) => 
                           P_tmp_7_25_port, S(24) => P_tmp_7_24_port, S(23) => 
                           P_tmp_7_23_port, S(22) => P_tmp_7_22_port, S(21) => 
                           P_tmp_7_21_port, S(20) => P_tmp_7_20_port, S(19) => 
                           P_tmp_7_19_port, S(18) => P_tmp_7_18_port, S(17) => 
                           P_tmp_7_17_port, S(16) => P_tmp_7_16_port, S(15) => 
                           P_tmp_7_15_port, S(14) => P_tmp_7_14_port, S(13) => 
                           P_tmp_7_13_port, S(12) => P_tmp_7_12_port, S(11) => 
                           P_tmp_7_11_port, S(10) => P_tmp_7_10_port, S(9) => 
                           P_tmp_7_9_port, S(8) => P_tmp_7_8_port, S(7) => 
                           P_tmp_7_7_port, S(6) => P_tmp_7_6_port, S(5) => 
                           P_tmp_7_5_port, S(4) => P_tmp_7_4_port, S(3) => 
                           P_tmp_7_3_port, S(2) => P_tmp_7_2_port, S(1) => 
                           P_tmp_7_1_port, S(0) => P_tmp_7_0_port, Co => n_1286
                           );
   RCAi_7 : RCA_NBIT64_8 port map( A(63) => P_tmp_7_63_port, A(62) => 
                           P_tmp_7_62_port, A(61) => P_tmp_7_61_port, A(60) => 
                           P_tmp_7_60_port, A(59) => P_tmp_7_59_port, A(58) => 
                           P_tmp_7_58_port, A(57) => P_tmp_7_57_port, A(56) => 
                           P_tmp_7_56_port, A(55) => P_tmp_7_55_port, A(54) => 
                           P_tmp_7_54_port, A(53) => P_tmp_7_53_port, A(52) => 
                           P_tmp_7_52_port, A(51) => P_tmp_7_51_port, A(50) => 
                           P_tmp_7_50_port, A(49) => P_tmp_7_49_port, A(48) => 
                           P_tmp_7_48_port, A(47) => P_tmp_7_47_port, A(46) => 
                           P_tmp_7_46_port, A(45) => P_tmp_7_45_port, A(44) => 
                           P_tmp_7_44_port, A(43) => P_tmp_7_43_port, A(42) => 
                           P_tmp_7_42_port, A(41) => P_tmp_7_41_port, A(40) => 
                           P_tmp_7_40_port, A(39) => P_tmp_7_39_port, A(38) => 
                           P_tmp_7_38_port, A(37) => P_tmp_7_37_port, A(36) => 
                           P_tmp_7_36_port, A(35) => P_tmp_7_35_port, A(34) => 
                           P_tmp_7_34_port, A(33) => P_tmp_7_33_port, A(32) => 
                           P_tmp_7_32_port, A(31) => P_tmp_7_31_port, A(30) => 
                           P_tmp_7_30_port, A(29) => P_tmp_7_29_port, A(28) => 
                           P_tmp_7_28_port, A(27) => P_tmp_7_27_port, A(26) => 
                           P_tmp_7_26_port, A(25) => P_tmp_7_25_port, A(24) => 
                           P_tmp_7_24_port, A(23) => P_tmp_7_23_port, A(22) => 
                           P_tmp_7_22_port, A(21) => P_tmp_7_21_port, A(20) => 
                           P_tmp_7_20_port, A(19) => P_tmp_7_19_port, A(18) => 
                           P_tmp_7_18_port, A(17) => P_tmp_7_17_port, A(16) => 
                           P_tmp_7_16_port, A(15) => P_tmp_7_15_port, A(14) => 
                           P_tmp_7_14_port, A(13) => P_tmp_7_13_port, A(12) => 
                           P_tmp_7_12_port, A(11) => P_tmp_7_11_port, A(10) => 
                           P_tmp_7_10_port, A(9) => P_tmp_7_9_port, A(8) => 
                           P_tmp_7_8_port, A(7) => P_tmp_7_7_port, A(6) => 
                           P_tmp_7_6_port, A(5) => P_tmp_7_5_port, A(4) => 
                           P_tmp_7_4_port, A(3) => P_tmp_7_3_port, A(2) => 
                           P_tmp_7_2_port, A(1) => P_tmp_7_1_port, A(0) => 
                           P_tmp_7_0_port, B(63) => OUT_MUX_8_63_port, B(62) =>
                           OUT_MUX_8_62_port, B(61) => OUT_MUX_8_61_port, B(60)
                           => OUT_MUX_8_60_port, B(59) => OUT_MUX_8_59_port, 
                           B(58) => OUT_MUX_8_58_port, B(57) => 
                           OUT_MUX_8_57_port, B(56) => OUT_MUX_8_56_port, B(55)
                           => OUT_MUX_8_55_port, B(54) => OUT_MUX_8_54_port, 
                           B(53) => OUT_MUX_8_53_port, B(52) => 
                           OUT_MUX_8_52_port, B(51) => OUT_MUX_8_51_port, B(50)
                           => OUT_MUX_8_50_port, B(49) => OUT_MUX_8_49_port, 
                           B(48) => OUT_MUX_8_48_port, B(47) => 
                           OUT_MUX_8_47_port, B(46) => OUT_MUX_8_46_port, B(45)
                           => OUT_MUX_8_45_port, B(44) => OUT_MUX_8_44_port, 
                           B(43) => OUT_MUX_8_43_port, B(42) => 
                           OUT_MUX_8_42_port, B(41) => OUT_MUX_8_41_port, B(40)
                           => OUT_MUX_8_40_port, B(39) => OUT_MUX_8_39_port, 
                           B(38) => OUT_MUX_8_38_port, B(37) => 
                           OUT_MUX_8_37_port, B(36) => OUT_MUX_8_36_port, B(35)
                           => OUT_MUX_8_35_port, B(34) => OUT_MUX_8_34_port, 
                           B(33) => OUT_MUX_8_33_port, B(32) => 
                           OUT_MUX_8_32_port, B(31) => OUT_MUX_8_31_port, B(30)
                           => OUT_MUX_8_30_port, B(29) => OUT_MUX_8_29_port, 
                           B(28) => OUT_MUX_8_28_port, B(27) => 
                           OUT_MUX_8_27_port, B(26) => OUT_MUX_8_26_port, B(25)
                           => OUT_MUX_8_25_port, B(24) => OUT_MUX_8_24_port, 
                           B(23) => OUT_MUX_8_23_port, B(22) => 
                           OUT_MUX_8_22_port, B(21) => OUT_MUX_8_21_port, B(20)
                           => OUT_MUX_8_20_port, B(19) => OUT_MUX_8_19_port, 
                           B(18) => OUT_MUX_8_18_port, B(17) => 
                           OUT_MUX_8_17_port, B(16) => OUT_MUX_8_16_port, B(15)
                           => OUT_MUX_8_15_port, B(14) => OUT_MUX_8_14_port, 
                           B(13) => OUT_MUX_8_13_port, B(12) => 
                           OUT_MUX_8_12_port, B(11) => OUT_MUX_8_11_port, B(10)
                           => OUT_MUX_8_10_port, B(9) => OUT_MUX_8_9_port, B(8)
                           => OUT_MUX_8_8_port, B(7) => OUT_MUX_8_7_port, B(6) 
                           => OUT_MUX_8_6_port, B(5) => OUT_MUX_8_5_port, B(4) 
                           => OUT_MUX_8_4_port, B(3) => OUT_MUX_8_3_port, B(2) 
                           => OUT_MUX_8_2_port, B(1) => OUT_MUX_8_1_port, B(0) 
                           => OUT_MUX_8_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_8_63_port, S(62) => P_tmp_8_62_port, S(61) => 
                           P_tmp_8_61_port, S(60) => P_tmp_8_60_port, S(59) => 
                           P_tmp_8_59_port, S(58) => P_tmp_8_58_port, S(57) => 
                           P_tmp_8_57_port, S(56) => P_tmp_8_56_port, S(55) => 
                           P_tmp_8_55_port, S(54) => P_tmp_8_54_port, S(53) => 
                           P_tmp_8_53_port, S(52) => P_tmp_8_52_port, S(51) => 
                           P_tmp_8_51_port, S(50) => P_tmp_8_50_port, S(49) => 
                           P_tmp_8_49_port, S(48) => P_tmp_8_48_port, S(47) => 
                           P_tmp_8_47_port, S(46) => P_tmp_8_46_port, S(45) => 
                           P_tmp_8_45_port, S(44) => P_tmp_8_44_port, S(43) => 
                           P_tmp_8_43_port, S(42) => P_tmp_8_42_port, S(41) => 
                           P_tmp_8_41_port, S(40) => P_tmp_8_40_port, S(39) => 
                           P_tmp_8_39_port, S(38) => P_tmp_8_38_port, S(37) => 
                           P_tmp_8_37_port, S(36) => P_tmp_8_36_port, S(35) => 
                           P_tmp_8_35_port, S(34) => P_tmp_8_34_port, S(33) => 
                           P_tmp_8_33_port, S(32) => P_tmp_8_32_port, S(31) => 
                           P_tmp_8_31_port, S(30) => P_tmp_8_30_port, S(29) => 
                           P_tmp_8_29_port, S(28) => P_tmp_8_28_port, S(27) => 
                           P_tmp_8_27_port, S(26) => P_tmp_8_26_port, S(25) => 
                           P_tmp_8_25_port, S(24) => P_tmp_8_24_port, S(23) => 
                           P_tmp_8_23_port, S(22) => P_tmp_8_22_port, S(21) => 
                           P_tmp_8_21_port, S(20) => P_tmp_8_20_port, S(19) => 
                           P_tmp_8_19_port, S(18) => P_tmp_8_18_port, S(17) => 
                           P_tmp_8_17_port, S(16) => P_tmp_8_16_port, S(15) => 
                           P_tmp_8_15_port, S(14) => P_tmp_8_14_port, S(13) => 
                           P_tmp_8_13_port, S(12) => P_tmp_8_12_port, S(11) => 
                           P_tmp_8_11_port, S(10) => P_tmp_8_10_port, S(9) => 
                           P_tmp_8_9_port, S(8) => P_tmp_8_8_port, S(7) => 
                           P_tmp_8_7_port, S(6) => P_tmp_8_6_port, S(5) => 
                           P_tmp_8_5_port, S(4) => P_tmp_8_4_port, S(3) => 
                           P_tmp_8_3_port, S(2) => P_tmp_8_2_port, S(1) => 
                           P_tmp_8_1_port, S(0) => P_tmp_8_0_port, Co => n_1287
                           );
   RCAi_8 : RCA_NBIT64_7 port map( A(63) => P_tmp_8_63_port, A(62) => 
                           P_tmp_8_62_port, A(61) => P_tmp_8_61_port, A(60) => 
                           P_tmp_8_60_port, A(59) => P_tmp_8_59_port, A(58) => 
                           P_tmp_8_58_port, A(57) => P_tmp_8_57_port, A(56) => 
                           P_tmp_8_56_port, A(55) => P_tmp_8_55_port, A(54) => 
                           P_tmp_8_54_port, A(53) => P_tmp_8_53_port, A(52) => 
                           P_tmp_8_52_port, A(51) => P_tmp_8_51_port, A(50) => 
                           P_tmp_8_50_port, A(49) => P_tmp_8_49_port, A(48) => 
                           P_tmp_8_48_port, A(47) => P_tmp_8_47_port, A(46) => 
                           P_tmp_8_46_port, A(45) => P_tmp_8_45_port, A(44) => 
                           P_tmp_8_44_port, A(43) => P_tmp_8_43_port, A(42) => 
                           P_tmp_8_42_port, A(41) => P_tmp_8_41_port, A(40) => 
                           P_tmp_8_40_port, A(39) => P_tmp_8_39_port, A(38) => 
                           P_tmp_8_38_port, A(37) => P_tmp_8_37_port, A(36) => 
                           P_tmp_8_36_port, A(35) => P_tmp_8_35_port, A(34) => 
                           P_tmp_8_34_port, A(33) => P_tmp_8_33_port, A(32) => 
                           P_tmp_8_32_port, A(31) => P_tmp_8_31_port, A(30) => 
                           P_tmp_8_30_port, A(29) => P_tmp_8_29_port, A(28) => 
                           P_tmp_8_28_port, A(27) => P_tmp_8_27_port, A(26) => 
                           P_tmp_8_26_port, A(25) => P_tmp_8_25_port, A(24) => 
                           P_tmp_8_24_port, A(23) => P_tmp_8_23_port, A(22) => 
                           P_tmp_8_22_port, A(21) => P_tmp_8_21_port, A(20) => 
                           P_tmp_8_20_port, A(19) => P_tmp_8_19_port, A(18) => 
                           P_tmp_8_18_port, A(17) => P_tmp_8_17_port, A(16) => 
                           P_tmp_8_16_port, A(15) => P_tmp_8_15_port, A(14) => 
                           P_tmp_8_14_port, A(13) => P_tmp_8_13_port, A(12) => 
                           P_tmp_8_12_port, A(11) => P_tmp_8_11_port, A(10) => 
                           P_tmp_8_10_port, A(9) => P_tmp_8_9_port, A(8) => 
                           P_tmp_8_8_port, A(7) => P_tmp_8_7_port, A(6) => 
                           P_tmp_8_6_port, A(5) => P_tmp_8_5_port, A(4) => 
                           P_tmp_8_4_port, A(3) => P_tmp_8_3_port, A(2) => 
                           P_tmp_8_2_port, A(1) => P_tmp_8_1_port, A(0) => 
                           P_tmp_8_0_port, B(63) => OUT_MUX_9_63_port, B(62) =>
                           OUT_MUX_9_62_port, B(61) => OUT_MUX_9_61_port, B(60)
                           => OUT_MUX_9_60_port, B(59) => OUT_MUX_9_59_port, 
                           B(58) => OUT_MUX_9_58_port, B(57) => 
                           OUT_MUX_9_57_port, B(56) => OUT_MUX_9_56_port, B(55)
                           => OUT_MUX_9_55_port, B(54) => OUT_MUX_9_54_port, 
                           B(53) => OUT_MUX_9_53_port, B(52) => 
                           OUT_MUX_9_52_port, B(51) => OUT_MUX_9_51_port, B(50)
                           => OUT_MUX_9_50_port, B(49) => OUT_MUX_9_49_port, 
                           B(48) => OUT_MUX_9_48_port, B(47) => 
                           OUT_MUX_9_47_port, B(46) => OUT_MUX_9_46_port, B(45)
                           => OUT_MUX_9_45_port, B(44) => OUT_MUX_9_44_port, 
                           B(43) => OUT_MUX_9_43_port, B(42) => 
                           OUT_MUX_9_42_port, B(41) => OUT_MUX_9_41_port, B(40)
                           => OUT_MUX_9_40_port, B(39) => OUT_MUX_9_39_port, 
                           B(38) => OUT_MUX_9_38_port, B(37) => 
                           OUT_MUX_9_37_port, B(36) => OUT_MUX_9_36_port, B(35)
                           => OUT_MUX_9_35_port, B(34) => OUT_MUX_9_34_port, 
                           B(33) => OUT_MUX_9_33_port, B(32) => 
                           OUT_MUX_9_32_port, B(31) => OUT_MUX_9_31_port, B(30)
                           => OUT_MUX_9_30_port, B(29) => OUT_MUX_9_29_port, 
                           B(28) => OUT_MUX_9_28_port, B(27) => 
                           OUT_MUX_9_27_port, B(26) => OUT_MUX_9_26_port, B(25)
                           => OUT_MUX_9_25_port, B(24) => OUT_MUX_9_24_port, 
                           B(23) => OUT_MUX_9_23_port, B(22) => 
                           OUT_MUX_9_22_port, B(21) => OUT_MUX_9_21_port, B(20)
                           => OUT_MUX_9_20_port, B(19) => OUT_MUX_9_19_port, 
                           B(18) => OUT_MUX_9_18_port, B(17) => 
                           OUT_MUX_9_17_port, B(16) => OUT_MUX_9_16_port, B(15)
                           => OUT_MUX_9_15_port, B(14) => OUT_MUX_9_14_port, 
                           B(13) => OUT_MUX_9_13_port, B(12) => 
                           OUT_MUX_9_12_port, B(11) => OUT_MUX_9_11_port, B(10)
                           => OUT_MUX_9_10_port, B(9) => OUT_MUX_9_9_port, B(8)
                           => OUT_MUX_9_8_port, B(7) => OUT_MUX_9_7_port, B(6) 
                           => OUT_MUX_9_6_port, B(5) => OUT_MUX_9_5_port, B(4) 
                           => OUT_MUX_9_4_port, B(3) => OUT_MUX_9_3_port, B(2) 
                           => OUT_MUX_9_2_port, B(1) => OUT_MUX_9_1_port, B(0) 
                           => OUT_MUX_9_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_9_63_port, S(62) => P_tmp_9_62_port, S(61) => 
                           P_tmp_9_61_port, S(60) => P_tmp_9_60_port, S(59) => 
                           P_tmp_9_59_port, S(58) => P_tmp_9_58_port, S(57) => 
                           P_tmp_9_57_port, S(56) => P_tmp_9_56_port, S(55) => 
                           P_tmp_9_55_port, S(54) => P_tmp_9_54_port, S(53) => 
                           P_tmp_9_53_port, S(52) => P_tmp_9_52_port, S(51) => 
                           P_tmp_9_51_port, S(50) => P_tmp_9_50_port, S(49) => 
                           P_tmp_9_49_port, S(48) => P_tmp_9_48_port, S(47) => 
                           P_tmp_9_47_port, S(46) => P_tmp_9_46_port, S(45) => 
                           P_tmp_9_45_port, S(44) => P_tmp_9_44_port, S(43) => 
                           P_tmp_9_43_port, S(42) => P_tmp_9_42_port, S(41) => 
                           P_tmp_9_41_port, S(40) => P_tmp_9_40_port, S(39) => 
                           P_tmp_9_39_port, S(38) => P_tmp_9_38_port, S(37) => 
                           P_tmp_9_37_port, S(36) => P_tmp_9_36_port, S(35) => 
                           P_tmp_9_35_port, S(34) => P_tmp_9_34_port, S(33) => 
                           P_tmp_9_33_port, S(32) => P_tmp_9_32_port, S(31) => 
                           P_tmp_9_31_port, S(30) => P_tmp_9_30_port, S(29) => 
                           P_tmp_9_29_port, S(28) => P_tmp_9_28_port, S(27) => 
                           P_tmp_9_27_port, S(26) => P_tmp_9_26_port, S(25) => 
                           P_tmp_9_25_port, S(24) => P_tmp_9_24_port, S(23) => 
                           P_tmp_9_23_port, S(22) => P_tmp_9_22_port, S(21) => 
                           P_tmp_9_21_port, S(20) => P_tmp_9_20_port, S(19) => 
                           P_tmp_9_19_port, S(18) => P_tmp_9_18_port, S(17) => 
                           P_tmp_9_17_port, S(16) => P_tmp_9_16_port, S(15) => 
                           P_tmp_9_15_port, S(14) => P_tmp_9_14_port, S(13) => 
                           P_tmp_9_13_port, S(12) => P_tmp_9_12_port, S(11) => 
                           P_tmp_9_11_port, S(10) => P_tmp_9_10_port, S(9) => 
                           P_tmp_9_9_port, S(8) => P_tmp_9_8_port, S(7) => 
                           P_tmp_9_7_port, S(6) => P_tmp_9_6_port, S(5) => 
                           P_tmp_9_5_port, S(4) => P_tmp_9_4_port, S(3) => 
                           P_tmp_9_3_port, S(2) => P_tmp_9_2_port, S(1) => 
                           P_tmp_9_1_port, S(0) => P_tmp_9_0_port, Co => n_1288
                           );
   RCAi_9 : RCA_NBIT64_6 port map( A(63) => P_tmp_9_63_port, A(62) => 
                           P_tmp_9_62_port, A(61) => P_tmp_9_61_port, A(60) => 
                           P_tmp_9_60_port, A(59) => P_tmp_9_59_port, A(58) => 
                           P_tmp_9_58_port, A(57) => P_tmp_9_57_port, A(56) => 
                           P_tmp_9_56_port, A(55) => P_tmp_9_55_port, A(54) => 
                           P_tmp_9_54_port, A(53) => P_tmp_9_53_port, A(52) => 
                           P_tmp_9_52_port, A(51) => P_tmp_9_51_port, A(50) => 
                           P_tmp_9_50_port, A(49) => P_tmp_9_49_port, A(48) => 
                           P_tmp_9_48_port, A(47) => P_tmp_9_47_port, A(46) => 
                           P_tmp_9_46_port, A(45) => P_tmp_9_45_port, A(44) => 
                           P_tmp_9_44_port, A(43) => P_tmp_9_43_port, A(42) => 
                           P_tmp_9_42_port, A(41) => P_tmp_9_41_port, A(40) => 
                           P_tmp_9_40_port, A(39) => P_tmp_9_39_port, A(38) => 
                           P_tmp_9_38_port, A(37) => P_tmp_9_37_port, A(36) => 
                           P_tmp_9_36_port, A(35) => P_tmp_9_35_port, A(34) => 
                           P_tmp_9_34_port, A(33) => P_tmp_9_33_port, A(32) => 
                           P_tmp_9_32_port, A(31) => P_tmp_9_31_port, A(30) => 
                           P_tmp_9_30_port, A(29) => P_tmp_9_29_port, A(28) => 
                           P_tmp_9_28_port, A(27) => P_tmp_9_27_port, A(26) => 
                           P_tmp_9_26_port, A(25) => P_tmp_9_25_port, A(24) => 
                           P_tmp_9_24_port, A(23) => P_tmp_9_23_port, A(22) => 
                           P_tmp_9_22_port, A(21) => P_tmp_9_21_port, A(20) => 
                           P_tmp_9_20_port, A(19) => P_tmp_9_19_port, A(18) => 
                           P_tmp_9_18_port, A(17) => P_tmp_9_17_port, A(16) => 
                           P_tmp_9_16_port, A(15) => P_tmp_9_15_port, A(14) => 
                           P_tmp_9_14_port, A(13) => P_tmp_9_13_port, A(12) => 
                           P_tmp_9_12_port, A(11) => P_tmp_9_11_port, A(10) => 
                           P_tmp_9_10_port, A(9) => P_tmp_9_9_port, A(8) => 
                           P_tmp_9_8_port, A(7) => P_tmp_9_7_port, A(6) => 
                           P_tmp_9_6_port, A(5) => P_tmp_9_5_port, A(4) => 
                           P_tmp_9_4_port, A(3) => P_tmp_9_3_port, A(2) => 
                           P_tmp_9_2_port, A(1) => P_tmp_9_1_port, A(0) => 
                           P_tmp_9_0_port, B(63) => OUT_MUX_10_63_port, B(62) 
                           => OUT_MUX_10_62_port, B(61) => OUT_MUX_10_61_port, 
                           B(60) => OUT_MUX_10_60_port, B(59) => 
                           OUT_MUX_10_59_port, B(58) => OUT_MUX_10_58_port, 
                           B(57) => OUT_MUX_10_57_port, B(56) => 
                           OUT_MUX_10_56_port, B(55) => OUT_MUX_10_55_port, 
                           B(54) => OUT_MUX_10_54_port, B(53) => 
                           OUT_MUX_10_53_port, B(52) => OUT_MUX_10_52_port, 
                           B(51) => OUT_MUX_10_51_port, B(50) => 
                           OUT_MUX_10_50_port, B(49) => OUT_MUX_10_49_port, 
                           B(48) => OUT_MUX_10_48_port, B(47) => 
                           OUT_MUX_10_47_port, B(46) => OUT_MUX_10_46_port, 
                           B(45) => OUT_MUX_10_45_port, B(44) => 
                           OUT_MUX_10_44_port, B(43) => OUT_MUX_10_43_port, 
                           B(42) => OUT_MUX_10_42_port, B(41) => 
                           OUT_MUX_10_41_port, B(40) => OUT_MUX_10_40_port, 
                           B(39) => OUT_MUX_10_39_port, B(38) => 
                           OUT_MUX_10_38_port, B(37) => OUT_MUX_10_37_port, 
                           B(36) => OUT_MUX_10_36_port, B(35) => 
                           OUT_MUX_10_35_port, B(34) => OUT_MUX_10_34_port, 
                           B(33) => OUT_MUX_10_33_port, B(32) => 
                           OUT_MUX_10_32_port, B(31) => OUT_MUX_10_31_port, 
                           B(30) => OUT_MUX_10_30_port, B(29) => 
                           OUT_MUX_10_29_port, B(28) => OUT_MUX_10_28_port, 
                           B(27) => OUT_MUX_10_27_port, B(26) => 
                           OUT_MUX_10_26_port, B(25) => OUT_MUX_10_25_port, 
                           B(24) => OUT_MUX_10_24_port, B(23) => 
                           OUT_MUX_10_23_port, B(22) => OUT_MUX_10_22_port, 
                           B(21) => OUT_MUX_10_21_port, B(20) => 
                           OUT_MUX_10_20_port, B(19) => OUT_MUX_10_19_port, 
                           B(18) => OUT_MUX_10_18_port, B(17) => 
                           OUT_MUX_10_17_port, B(16) => OUT_MUX_10_16_port, 
                           B(15) => OUT_MUX_10_15_port, B(14) => 
                           OUT_MUX_10_14_port, B(13) => OUT_MUX_10_13_port, 
                           B(12) => OUT_MUX_10_12_port, B(11) => 
                           OUT_MUX_10_11_port, B(10) => OUT_MUX_10_10_port, 
                           B(9) => OUT_MUX_10_9_port, B(8) => OUT_MUX_10_8_port
                           , B(7) => OUT_MUX_10_7_port, B(6) => 
                           OUT_MUX_10_6_port, B(5) => OUT_MUX_10_5_port, B(4) 
                           => OUT_MUX_10_4_port, B(3) => OUT_MUX_10_3_port, 
                           B(2) => OUT_MUX_10_2_port, B(1) => OUT_MUX_10_1_port
                           , B(0) => OUT_MUX_10_0_port, Ci => X_Logic0_port, 
                           S(63) => P_tmp_10_63_port, S(62) => P_tmp_10_62_port
                           , S(61) => P_tmp_10_61_port, S(60) => 
                           P_tmp_10_60_port, S(59) => P_tmp_10_59_port, S(58) 
                           => P_tmp_10_58_port, S(57) => P_tmp_10_57_port, 
                           S(56) => P_tmp_10_56_port, S(55) => P_tmp_10_55_port
                           , S(54) => P_tmp_10_54_port, S(53) => 
                           P_tmp_10_53_port, S(52) => P_tmp_10_52_port, S(51) 
                           => P_tmp_10_51_port, S(50) => P_tmp_10_50_port, 
                           S(49) => P_tmp_10_49_port, S(48) => P_tmp_10_48_port
                           , S(47) => P_tmp_10_47_port, S(46) => 
                           P_tmp_10_46_port, S(45) => P_tmp_10_45_port, S(44) 
                           => P_tmp_10_44_port, S(43) => P_tmp_10_43_port, 
                           S(42) => P_tmp_10_42_port, S(41) => P_tmp_10_41_port
                           , S(40) => P_tmp_10_40_port, S(39) => 
                           P_tmp_10_39_port, S(38) => P_tmp_10_38_port, S(37) 
                           => P_tmp_10_37_port, S(36) => P_tmp_10_36_port, 
                           S(35) => P_tmp_10_35_port, S(34) => P_tmp_10_34_port
                           , S(33) => P_tmp_10_33_port, S(32) => 
                           P_tmp_10_32_port, S(31) => P_tmp_10_31_port, S(30) 
                           => P_tmp_10_30_port, S(29) => P_tmp_10_29_port, 
                           S(28) => P_tmp_10_28_port, S(27) => P_tmp_10_27_port
                           , S(26) => P_tmp_10_26_port, S(25) => 
                           P_tmp_10_25_port, S(24) => P_tmp_10_24_port, S(23) 
                           => P_tmp_10_23_port, S(22) => P_tmp_10_22_port, 
                           S(21) => P_tmp_10_21_port, S(20) => P_tmp_10_20_port
                           , S(19) => P_tmp_10_19_port, S(18) => 
                           P_tmp_10_18_port, S(17) => P_tmp_10_17_port, S(16) 
                           => P_tmp_10_16_port, S(15) => P_tmp_10_15_port, 
                           S(14) => P_tmp_10_14_port, S(13) => P_tmp_10_13_port
                           , S(12) => P_tmp_10_12_port, S(11) => 
                           P_tmp_10_11_port, S(10) => P_tmp_10_10_port, S(9) =>
                           P_tmp_10_9_port, S(8) => P_tmp_10_8_port, S(7) => 
                           P_tmp_10_7_port, S(6) => P_tmp_10_6_port, S(5) => 
                           P_tmp_10_5_port, S(4) => P_tmp_10_4_port, S(3) => 
                           P_tmp_10_3_port, S(2) => P_tmp_10_2_port, S(1) => 
                           P_tmp_10_1_port, S(0) => P_tmp_10_0_port, Co => 
                           n_1289);
   RCAi_10 : RCA_NBIT64_5 port map( A(63) => P_tmp_10_63_port, A(62) => 
                           P_tmp_10_62_port, A(61) => P_tmp_10_61_port, A(60) 
                           => P_tmp_10_60_port, A(59) => P_tmp_10_59_port, 
                           A(58) => P_tmp_10_58_port, A(57) => P_tmp_10_57_port
                           , A(56) => P_tmp_10_56_port, A(55) => 
                           P_tmp_10_55_port, A(54) => P_tmp_10_54_port, A(53) 
                           => P_tmp_10_53_port, A(52) => P_tmp_10_52_port, 
                           A(51) => P_tmp_10_51_port, A(50) => P_tmp_10_50_port
                           , A(49) => P_tmp_10_49_port, A(48) => 
                           P_tmp_10_48_port, A(47) => P_tmp_10_47_port, A(46) 
                           => P_tmp_10_46_port, A(45) => P_tmp_10_45_port, 
                           A(44) => P_tmp_10_44_port, A(43) => P_tmp_10_43_port
                           , A(42) => P_tmp_10_42_port, A(41) => 
                           P_tmp_10_41_port, A(40) => P_tmp_10_40_port, A(39) 
                           => P_tmp_10_39_port, A(38) => P_tmp_10_38_port, 
                           A(37) => P_tmp_10_37_port, A(36) => P_tmp_10_36_port
                           , A(35) => P_tmp_10_35_port, A(34) => 
                           P_tmp_10_34_port, A(33) => P_tmp_10_33_port, A(32) 
                           => P_tmp_10_32_port, A(31) => P_tmp_10_31_port, 
                           A(30) => P_tmp_10_30_port, A(29) => P_tmp_10_29_port
                           , A(28) => P_tmp_10_28_port, A(27) => 
                           P_tmp_10_27_port, A(26) => P_tmp_10_26_port, A(25) 
                           => P_tmp_10_25_port, A(24) => P_tmp_10_24_port, 
                           A(23) => P_tmp_10_23_port, A(22) => P_tmp_10_22_port
                           , A(21) => P_tmp_10_21_port, A(20) => 
                           P_tmp_10_20_port, A(19) => P_tmp_10_19_port, A(18) 
                           => P_tmp_10_18_port, A(17) => P_tmp_10_17_port, 
                           A(16) => P_tmp_10_16_port, A(15) => P_tmp_10_15_port
                           , A(14) => P_tmp_10_14_port, A(13) => 
                           P_tmp_10_13_port, A(12) => P_tmp_10_12_port, A(11) 
                           => P_tmp_10_11_port, A(10) => P_tmp_10_10_port, A(9)
                           => P_tmp_10_9_port, A(8) => P_tmp_10_8_port, A(7) =>
                           P_tmp_10_7_port, A(6) => P_tmp_10_6_port, A(5) => 
                           P_tmp_10_5_port, A(4) => P_tmp_10_4_port, A(3) => 
                           P_tmp_10_3_port, A(2) => P_tmp_10_2_port, A(1) => 
                           P_tmp_10_1_port, A(0) => P_tmp_10_0_port, B(63) => 
                           OUT_MUX_11_63_port, B(62) => OUT_MUX_11_62_port, 
                           B(61) => OUT_MUX_11_61_port, B(60) => 
                           OUT_MUX_11_60_port, B(59) => OUT_MUX_11_59_port, 
                           B(58) => OUT_MUX_11_58_port, B(57) => 
                           OUT_MUX_11_57_port, B(56) => OUT_MUX_11_56_port, 
                           B(55) => OUT_MUX_11_55_port, B(54) => 
                           OUT_MUX_11_54_port, B(53) => OUT_MUX_11_53_port, 
                           B(52) => OUT_MUX_11_52_port, B(51) => 
                           OUT_MUX_11_51_port, B(50) => OUT_MUX_11_50_port, 
                           B(49) => OUT_MUX_11_49_port, B(48) => 
                           OUT_MUX_11_48_port, B(47) => OUT_MUX_11_47_port, 
                           B(46) => OUT_MUX_11_46_port, B(45) => 
                           OUT_MUX_11_45_port, B(44) => OUT_MUX_11_44_port, 
                           B(43) => OUT_MUX_11_43_port, B(42) => 
                           OUT_MUX_11_42_port, B(41) => OUT_MUX_11_41_port, 
                           B(40) => OUT_MUX_11_40_port, B(39) => 
                           OUT_MUX_11_39_port, B(38) => OUT_MUX_11_38_port, 
                           B(37) => OUT_MUX_11_37_port, B(36) => 
                           OUT_MUX_11_36_port, B(35) => OUT_MUX_11_35_port, 
                           B(34) => OUT_MUX_11_34_port, B(33) => 
                           OUT_MUX_11_33_port, B(32) => OUT_MUX_11_32_port, 
                           B(31) => OUT_MUX_11_31_port, B(30) => 
                           OUT_MUX_11_30_port, B(29) => OUT_MUX_11_29_port, 
                           B(28) => OUT_MUX_11_28_port, B(27) => 
                           OUT_MUX_11_27_port, B(26) => OUT_MUX_11_26_port, 
                           B(25) => OUT_MUX_11_25_port, B(24) => 
                           OUT_MUX_11_24_port, B(23) => OUT_MUX_11_23_port, 
                           B(22) => OUT_MUX_11_22_port, B(21) => 
                           OUT_MUX_11_21_port, B(20) => OUT_MUX_11_20_port, 
                           B(19) => OUT_MUX_11_19_port, B(18) => 
                           OUT_MUX_11_18_port, B(17) => OUT_MUX_11_17_port, 
                           B(16) => OUT_MUX_11_16_port, B(15) => 
                           OUT_MUX_11_15_port, B(14) => OUT_MUX_11_14_port, 
                           B(13) => OUT_MUX_11_13_port, B(12) => 
                           OUT_MUX_11_12_port, B(11) => OUT_MUX_11_11_port, 
                           B(10) => OUT_MUX_11_10_port, B(9) => 
                           OUT_MUX_11_9_port, B(8) => OUT_MUX_11_8_port, B(7) 
                           => OUT_MUX_11_7_port, B(6) => OUT_MUX_11_6_port, 
                           B(5) => OUT_MUX_11_5_port, B(4) => OUT_MUX_11_4_port
                           , B(3) => OUT_MUX_11_3_port, B(2) => 
                           OUT_MUX_11_2_port, B(1) => OUT_MUX_11_1_port, B(0) 
                           => OUT_MUX_11_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_11_63_port, S(62) => P_tmp_11_62_port, S(61) 
                           => P_tmp_11_61_port, S(60) => P_tmp_11_60_port, 
                           S(59) => P_tmp_11_59_port, S(58) => P_tmp_11_58_port
                           , S(57) => P_tmp_11_57_port, S(56) => 
                           P_tmp_11_56_port, S(55) => P_tmp_11_55_port, S(54) 
                           => P_tmp_11_54_port, S(53) => P_tmp_11_53_port, 
                           S(52) => P_tmp_11_52_port, S(51) => P_tmp_11_51_port
                           , S(50) => P_tmp_11_50_port, S(49) => 
                           P_tmp_11_49_port, S(48) => P_tmp_11_48_port, S(47) 
                           => P_tmp_11_47_port, S(46) => P_tmp_11_46_port, 
                           S(45) => P_tmp_11_45_port, S(44) => P_tmp_11_44_port
                           , S(43) => P_tmp_11_43_port, S(42) => 
                           P_tmp_11_42_port, S(41) => P_tmp_11_41_port, S(40) 
                           => P_tmp_11_40_port, S(39) => P_tmp_11_39_port, 
                           S(38) => P_tmp_11_38_port, S(37) => P_tmp_11_37_port
                           , S(36) => P_tmp_11_36_port, S(35) => 
                           P_tmp_11_35_port, S(34) => P_tmp_11_34_port, S(33) 
                           => P_tmp_11_33_port, S(32) => P_tmp_11_32_port, 
                           S(31) => P_tmp_11_31_port, S(30) => P_tmp_11_30_port
                           , S(29) => P_tmp_11_29_port, S(28) => 
                           P_tmp_11_28_port, S(27) => P_tmp_11_27_port, S(26) 
                           => P_tmp_11_26_port, S(25) => P_tmp_11_25_port, 
                           S(24) => P_tmp_11_24_port, S(23) => P_tmp_11_23_port
                           , S(22) => P_tmp_11_22_port, S(21) => 
                           P_tmp_11_21_port, S(20) => P_tmp_11_20_port, S(19) 
                           => P_tmp_11_19_port, S(18) => P_tmp_11_18_port, 
                           S(17) => P_tmp_11_17_port, S(16) => P_tmp_11_16_port
                           , S(15) => P_tmp_11_15_port, S(14) => 
                           P_tmp_11_14_port, S(13) => P_tmp_11_13_port, S(12) 
                           => P_tmp_11_12_port, S(11) => P_tmp_11_11_port, 
                           S(10) => P_tmp_11_10_port, S(9) => P_tmp_11_9_port, 
                           S(8) => P_tmp_11_8_port, S(7) => P_tmp_11_7_port, 
                           S(6) => P_tmp_11_6_port, S(5) => P_tmp_11_5_port, 
                           S(4) => P_tmp_11_4_port, S(3) => P_tmp_11_3_port, 
                           S(2) => P_tmp_11_2_port, S(1) => P_tmp_11_1_port, 
                           S(0) => P_tmp_11_0_port, Co => n_1290);
   RCAi_11 : RCA_NBIT64_4 port map( A(63) => P_tmp_11_63_port, A(62) => 
                           P_tmp_11_62_port, A(61) => P_tmp_11_61_port, A(60) 
                           => P_tmp_11_60_port, A(59) => P_tmp_11_59_port, 
                           A(58) => P_tmp_11_58_port, A(57) => P_tmp_11_57_port
                           , A(56) => P_tmp_11_56_port, A(55) => 
                           P_tmp_11_55_port, A(54) => P_tmp_11_54_port, A(53) 
                           => P_tmp_11_53_port, A(52) => P_tmp_11_52_port, 
                           A(51) => P_tmp_11_51_port, A(50) => P_tmp_11_50_port
                           , A(49) => P_tmp_11_49_port, A(48) => 
                           P_tmp_11_48_port, A(47) => P_tmp_11_47_port, A(46) 
                           => P_tmp_11_46_port, A(45) => P_tmp_11_45_port, 
                           A(44) => P_tmp_11_44_port, A(43) => P_tmp_11_43_port
                           , A(42) => P_tmp_11_42_port, A(41) => 
                           P_tmp_11_41_port, A(40) => P_tmp_11_40_port, A(39) 
                           => P_tmp_11_39_port, A(38) => P_tmp_11_38_port, 
                           A(37) => P_tmp_11_37_port, A(36) => P_tmp_11_36_port
                           , A(35) => P_tmp_11_35_port, A(34) => 
                           P_tmp_11_34_port, A(33) => P_tmp_11_33_port, A(32) 
                           => P_tmp_11_32_port, A(31) => P_tmp_11_31_port, 
                           A(30) => P_tmp_11_30_port, A(29) => P_tmp_11_29_port
                           , A(28) => P_tmp_11_28_port, A(27) => 
                           P_tmp_11_27_port, A(26) => P_tmp_11_26_port, A(25) 
                           => P_tmp_11_25_port, A(24) => P_tmp_11_24_port, 
                           A(23) => P_tmp_11_23_port, A(22) => P_tmp_11_22_port
                           , A(21) => P_tmp_11_21_port, A(20) => 
                           P_tmp_11_20_port, A(19) => P_tmp_11_19_port, A(18) 
                           => P_tmp_11_18_port, A(17) => P_tmp_11_17_port, 
                           A(16) => P_tmp_11_16_port, A(15) => P_tmp_11_15_port
                           , A(14) => P_tmp_11_14_port, A(13) => 
                           P_tmp_11_13_port, A(12) => P_tmp_11_12_port, A(11) 
                           => P_tmp_11_11_port, A(10) => P_tmp_11_10_port, A(9)
                           => P_tmp_11_9_port, A(8) => P_tmp_11_8_port, A(7) =>
                           P_tmp_11_7_port, A(6) => P_tmp_11_6_port, A(5) => 
                           P_tmp_11_5_port, A(4) => P_tmp_11_4_port, A(3) => 
                           P_tmp_11_3_port, A(2) => P_tmp_11_2_port, A(1) => 
                           P_tmp_11_1_port, A(0) => P_tmp_11_0_port, B(63) => 
                           OUT_MUX_12_63_port, B(62) => OUT_MUX_12_62_port, 
                           B(61) => OUT_MUX_12_61_port, B(60) => 
                           OUT_MUX_12_60_port, B(59) => OUT_MUX_12_59_port, 
                           B(58) => OUT_MUX_12_58_port, B(57) => 
                           OUT_MUX_12_57_port, B(56) => OUT_MUX_12_56_port, 
                           B(55) => OUT_MUX_12_55_port, B(54) => 
                           OUT_MUX_12_54_port, B(53) => OUT_MUX_12_53_port, 
                           B(52) => OUT_MUX_12_52_port, B(51) => 
                           OUT_MUX_12_51_port, B(50) => OUT_MUX_12_50_port, 
                           B(49) => OUT_MUX_12_49_port, B(48) => 
                           OUT_MUX_12_48_port, B(47) => OUT_MUX_12_47_port, 
                           B(46) => OUT_MUX_12_46_port, B(45) => 
                           OUT_MUX_12_45_port, B(44) => OUT_MUX_12_44_port, 
                           B(43) => OUT_MUX_12_43_port, B(42) => 
                           OUT_MUX_12_42_port, B(41) => OUT_MUX_12_41_port, 
                           B(40) => OUT_MUX_12_40_port, B(39) => 
                           OUT_MUX_12_39_port, B(38) => OUT_MUX_12_38_port, 
                           B(37) => OUT_MUX_12_37_port, B(36) => 
                           OUT_MUX_12_36_port, B(35) => OUT_MUX_12_35_port, 
                           B(34) => OUT_MUX_12_34_port, B(33) => 
                           OUT_MUX_12_33_port, B(32) => OUT_MUX_12_32_port, 
                           B(31) => OUT_MUX_12_31_port, B(30) => 
                           OUT_MUX_12_30_port, B(29) => OUT_MUX_12_29_port, 
                           B(28) => OUT_MUX_12_28_port, B(27) => 
                           OUT_MUX_12_27_port, B(26) => OUT_MUX_12_26_port, 
                           B(25) => OUT_MUX_12_25_port, B(24) => 
                           OUT_MUX_12_24_port, B(23) => OUT_MUX_12_23_port, 
                           B(22) => OUT_MUX_12_22_port, B(21) => 
                           OUT_MUX_12_21_port, B(20) => OUT_MUX_12_20_port, 
                           B(19) => OUT_MUX_12_19_port, B(18) => 
                           OUT_MUX_12_18_port, B(17) => OUT_MUX_12_17_port, 
                           B(16) => OUT_MUX_12_16_port, B(15) => 
                           OUT_MUX_12_15_port, B(14) => OUT_MUX_12_14_port, 
                           B(13) => OUT_MUX_12_13_port, B(12) => 
                           OUT_MUX_12_12_port, B(11) => OUT_MUX_12_11_port, 
                           B(10) => OUT_MUX_12_10_port, B(9) => 
                           OUT_MUX_12_9_port, B(8) => OUT_MUX_12_8_port, B(7) 
                           => OUT_MUX_12_7_port, B(6) => OUT_MUX_12_6_port, 
                           B(5) => OUT_MUX_12_5_port, B(4) => OUT_MUX_12_4_port
                           , B(3) => OUT_MUX_12_3_port, B(2) => 
                           OUT_MUX_12_2_port, B(1) => OUT_MUX_12_1_port, B(0) 
                           => OUT_MUX_12_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_12_63_port, S(62) => P_tmp_12_62_port, S(61) 
                           => P_tmp_12_61_port, S(60) => P_tmp_12_60_port, 
                           S(59) => P_tmp_12_59_port, S(58) => P_tmp_12_58_port
                           , S(57) => P_tmp_12_57_port, S(56) => 
                           P_tmp_12_56_port, S(55) => P_tmp_12_55_port, S(54) 
                           => P_tmp_12_54_port, S(53) => P_tmp_12_53_port, 
                           S(52) => P_tmp_12_52_port, S(51) => P_tmp_12_51_port
                           , S(50) => P_tmp_12_50_port, S(49) => 
                           P_tmp_12_49_port, S(48) => P_tmp_12_48_port, S(47) 
                           => P_tmp_12_47_port, S(46) => P_tmp_12_46_port, 
                           S(45) => P_tmp_12_45_port, S(44) => P_tmp_12_44_port
                           , S(43) => P_tmp_12_43_port, S(42) => 
                           P_tmp_12_42_port, S(41) => P_tmp_12_41_port, S(40) 
                           => P_tmp_12_40_port, S(39) => P_tmp_12_39_port, 
                           S(38) => P_tmp_12_38_port, S(37) => P_tmp_12_37_port
                           , S(36) => P_tmp_12_36_port, S(35) => 
                           P_tmp_12_35_port, S(34) => P_tmp_12_34_port, S(33) 
                           => P_tmp_12_33_port, S(32) => P_tmp_12_32_port, 
                           S(31) => P_tmp_12_31_port, S(30) => P_tmp_12_30_port
                           , S(29) => P_tmp_12_29_port, S(28) => 
                           P_tmp_12_28_port, S(27) => P_tmp_12_27_port, S(26) 
                           => P_tmp_12_26_port, S(25) => P_tmp_12_25_port, 
                           S(24) => P_tmp_12_24_port, S(23) => P_tmp_12_23_port
                           , S(22) => P_tmp_12_22_port, S(21) => 
                           P_tmp_12_21_port, S(20) => P_tmp_12_20_port, S(19) 
                           => P_tmp_12_19_port, S(18) => P_tmp_12_18_port, 
                           S(17) => P_tmp_12_17_port, S(16) => P_tmp_12_16_port
                           , S(15) => P_tmp_12_15_port, S(14) => 
                           P_tmp_12_14_port, S(13) => P_tmp_12_13_port, S(12) 
                           => P_tmp_12_12_port, S(11) => P_tmp_12_11_port, 
                           S(10) => P_tmp_12_10_port, S(9) => P_tmp_12_9_port, 
                           S(8) => P_tmp_12_8_port, S(7) => P_tmp_12_7_port, 
                           S(6) => P_tmp_12_6_port, S(5) => P_tmp_12_5_port, 
                           S(4) => P_tmp_12_4_port, S(3) => P_tmp_12_3_port, 
                           S(2) => P_tmp_12_2_port, S(1) => P_tmp_12_1_port, 
                           S(0) => P_tmp_12_0_port, Co => n_1291);
   RCAi_12 : RCA_NBIT64_3 port map( A(63) => P_tmp_12_63_port, A(62) => 
                           P_tmp_12_62_port, A(61) => P_tmp_12_61_port, A(60) 
                           => P_tmp_12_60_port, A(59) => P_tmp_12_59_port, 
                           A(58) => P_tmp_12_58_port, A(57) => P_tmp_12_57_port
                           , A(56) => P_tmp_12_56_port, A(55) => 
                           P_tmp_12_55_port, A(54) => P_tmp_12_54_port, A(53) 
                           => P_tmp_12_53_port, A(52) => P_tmp_12_52_port, 
                           A(51) => P_tmp_12_51_port, A(50) => P_tmp_12_50_port
                           , A(49) => P_tmp_12_49_port, A(48) => 
                           P_tmp_12_48_port, A(47) => P_tmp_12_47_port, A(46) 
                           => P_tmp_12_46_port, A(45) => P_tmp_12_45_port, 
                           A(44) => P_tmp_12_44_port, A(43) => P_tmp_12_43_port
                           , A(42) => P_tmp_12_42_port, A(41) => 
                           P_tmp_12_41_port, A(40) => P_tmp_12_40_port, A(39) 
                           => P_tmp_12_39_port, A(38) => P_tmp_12_38_port, 
                           A(37) => P_tmp_12_37_port, A(36) => P_tmp_12_36_port
                           , A(35) => P_tmp_12_35_port, A(34) => 
                           P_tmp_12_34_port, A(33) => P_tmp_12_33_port, A(32) 
                           => P_tmp_12_32_port, A(31) => P_tmp_12_31_port, 
                           A(30) => P_tmp_12_30_port, A(29) => P_tmp_12_29_port
                           , A(28) => P_tmp_12_28_port, A(27) => 
                           P_tmp_12_27_port, A(26) => P_tmp_12_26_port, A(25) 
                           => P_tmp_12_25_port, A(24) => P_tmp_12_24_port, 
                           A(23) => P_tmp_12_23_port, A(22) => P_tmp_12_22_port
                           , A(21) => P_tmp_12_21_port, A(20) => 
                           P_tmp_12_20_port, A(19) => P_tmp_12_19_port, A(18) 
                           => P_tmp_12_18_port, A(17) => P_tmp_12_17_port, 
                           A(16) => P_tmp_12_16_port, A(15) => P_tmp_12_15_port
                           , A(14) => P_tmp_12_14_port, A(13) => 
                           P_tmp_12_13_port, A(12) => P_tmp_12_12_port, A(11) 
                           => P_tmp_12_11_port, A(10) => P_tmp_12_10_port, A(9)
                           => P_tmp_12_9_port, A(8) => P_tmp_12_8_port, A(7) =>
                           P_tmp_12_7_port, A(6) => P_tmp_12_6_port, A(5) => 
                           P_tmp_12_5_port, A(4) => P_tmp_12_4_port, A(3) => 
                           P_tmp_12_3_port, A(2) => P_tmp_12_2_port, A(1) => 
                           P_tmp_12_1_port, A(0) => P_tmp_12_0_port, B(63) => 
                           OUT_MUX_13_63_port, B(62) => OUT_MUX_13_62_port, 
                           B(61) => OUT_MUX_13_61_port, B(60) => 
                           OUT_MUX_13_60_port, B(59) => OUT_MUX_13_59_port, 
                           B(58) => OUT_MUX_13_58_port, B(57) => 
                           OUT_MUX_13_57_port, B(56) => OUT_MUX_13_56_port, 
                           B(55) => OUT_MUX_13_55_port, B(54) => 
                           OUT_MUX_13_54_port, B(53) => OUT_MUX_13_53_port, 
                           B(52) => OUT_MUX_13_52_port, B(51) => 
                           OUT_MUX_13_51_port, B(50) => OUT_MUX_13_50_port, 
                           B(49) => OUT_MUX_13_49_port, B(48) => 
                           OUT_MUX_13_48_port, B(47) => OUT_MUX_13_47_port, 
                           B(46) => OUT_MUX_13_46_port, B(45) => 
                           OUT_MUX_13_45_port, B(44) => OUT_MUX_13_44_port, 
                           B(43) => OUT_MUX_13_43_port, B(42) => 
                           OUT_MUX_13_42_port, B(41) => OUT_MUX_13_41_port, 
                           B(40) => OUT_MUX_13_40_port, B(39) => 
                           OUT_MUX_13_39_port, B(38) => OUT_MUX_13_38_port, 
                           B(37) => OUT_MUX_13_37_port, B(36) => 
                           OUT_MUX_13_36_port, B(35) => OUT_MUX_13_35_port, 
                           B(34) => OUT_MUX_13_34_port, B(33) => 
                           OUT_MUX_13_33_port, B(32) => OUT_MUX_13_32_port, 
                           B(31) => OUT_MUX_13_31_port, B(30) => 
                           OUT_MUX_13_30_port, B(29) => OUT_MUX_13_29_port, 
                           B(28) => OUT_MUX_13_28_port, B(27) => 
                           OUT_MUX_13_27_port, B(26) => OUT_MUX_13_26_port, 
                           B(25) => OUT_MUX_13_25_port, B(24) => 
                           OUT_MUX_13_24_port, B(23) => OUT_MUX_13_23_port, 
                           B(22) => OUT_MUX_13_22_port, B(21) => 
                           OUT_MUX_13_21_port, B(20) => OUT_MUX_13_20_port, 
                           B(19) => OUT_MUX_13_19_port, B(18) => 
                           OUT_MUX_13_18_port, B(17) => OUT_MUX_13_17_port, 
                           B(16) => OUT_MUX_13_16_port, B(15) => 
                           OUT_MUX_13_15_port, B(14) => OUT_MUX_13_14_port, 
                           B(13) => OUT_MUX_13_13_port, B(12) => 
                           OUT_MUX_13_12_port, B(11) => OUT_MUX_13_11_port, 
                           B(10) => OUT_MUX_13_10_port, B(9) => 
                           OUT_MUX_13_9_port, B(8) => OUT_MUX_13_8_port, B(7) 
                           => OUT_MUX_13_7_port, B(6) => OUT_MUX_13_6_port, 
                           B(5) => OUT_MUX_13_5_port, B(4) => OUT_MUX_13_4_port
                           , B(3) => OUT_MUX_13_3_port, B(2) => 
                           OUT_MUX_13_2_port, B(1) => OUT_MUX_13_1_port, B(0) 
                           => OUT_MUX_13_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_13_63_port, S(62) => P_tmp_13_62_port, S(61) 
                           => P_tmp_13_61_port, S(60) => P_tmp_13_60_port, 
                           S(59) => P_tmp_13_59_port, S(58) => P_tmp_13_58_port
                           , S(57) => P_tmp_13_57_port, S(56) => 
                           P_tmp_13_56_port, S(55) => P_tmp_13_55_port, S(54) 
                           => P_tmp_13_54_port, S(53) => P_tmp_13_53_port, 
                           S(52) => P_tmp_13_52_port, S(51) => P_tmp_13_51_port
                           , S(50) => P_tmp_13_50_port, S(49) => 
                           P_tmp_13_49_port, S(48) => P_tmp_13_48_port, S(47) 
                           => P_tmp_13_47_port, S(46) => P_tmp_13_46_port, 
                           S(45) => P_tmp_13_45_port, S(44) => P_tmp_13_44_port
                           , S(43) => P_tmp_13_43_port, S(42) => 
                           P_tmp_13_42_port, S(41) => P_tmp_13_41_port, S(40) 
                           => P_tmp_13_40_port, S(39) => P_tmp_13_39_port, 
                           S(38) => P_tmp_13_38_port, S(37) => P_tmp_13_37_port
                           , S(36) => P_tmp_13_36_port, S(35) => 
                           P_tmp_13_35_port, S(34) => P_tmp_13_34_port, S(33) 
                           => P_tmp_13_33_port, S(32) => P_tmp_13_32_port, 
                           S(31) => P_tmp_13_31_port, S(30) => P_tmp_13_30_port
                           , S(29) => P_tmp_13_29_port, S(28) => 
                           P_tmp_13_28_port, S(27) => P_tmp_13_27_port, S(26) 
                           => P_tmp_13_26_port, S(25) => P_tmp_13_25_port, 
                           S(24) => P_tmp_13_24_port, S(23) => P_tmp_13_23_port
                           , S(22) => P_tmp_13_22_port, S(21) => 
                           P_tmp_13_21_port, S(20) => P_tmp_13_20_port, S(19) 
                           => P_tmp_13_19_port, S(18) => P_tmp_13_18_port, 
                           S(17) => P_tmp_13_17_port, S(16) => P_tmp_13_16_port
                           , S(15) => P_tmp_13_15_port, S(14) => 
                           P_tmp_13_14_port, S(13) => P_tmp_13_13_port, S(12) 
                           => P_tmp_13_12_port, S(11) => P_tmp_13_11_port, 
                           S(10) => P_tmp_13_10_port, S(9) => P_tmp_13_9_port, 
                           S(8) => P_tmp_13_8_port, S(7) => P_tmp_13_7_port, 
                           S(6) => P_tmp_13_6_port, S(5) => P_tmp_13_5_port, 
                           S(4) => P_tmp_13_4_port, S(3) => P_tmp_13_3_port, 
                           S(2) => P_tmp_13_2_port, S(1) => P_tmp_13_1_port, 
                           S(0) => P_tmp_13_0_port, Co => n_1292);
   RCAi_13 : RCA_NBIT64_2 port map( A(63) => P_tmp_13_63_port, A(62) => 
                           P_tmp_13_62_port, A(61) => P_tmp_13_61_port, A(60) 
                           => P_tmp_13_60_port, A(59) => P_tmp_13_59_port, 
                           A(58) => P_tmp_13_58_port, A(57) => P_tmp_13_57_port
                           , A(56) => P_tmp_13_56_port, A(55) => 
                           P_tmp_13_55_port, A(54) => P_tmp_13_54_port, A(53) 
                           => P_tmp_13_53_port, A(52) => P_tmp_13_52_port, 
                           A(51) => P_tmp_13_51_port, A(50) => P_tmp_13_50_port
                           , A(49) => P_tmp_13_49_port, A(48) => 
                           P_tmp_13_48_port, A(47) => P_tmp_13_47_port, A(46) 
                           => P_tmp_13_46_port, A(45) => P_tmp_13_45_port, 
                           A(44) => P_tmp_13_44_port, A(43) => P_tmp_13_43_port
                           , A(42) => P_tmp_13_42_port, A(41) => 
                           P_tmp_13_41_port, A(40) => P_tmp_13_40_port, A(39) 
                           => P_tmp_13_39_port, A(38) => P_tmp_13_38_port, 
                           A(37) => P_tmp_13_37_port, A(36) => P_tmp_13_36_port
                           , A(35) => P_tmp_13_35_port, A(34) => 
                           P_tmp_13_34_port, A(33) => P_tmp_13_33_port, A(32) 
                           => P_tmp_13_32_port, A(31) => P_tmp_13_31_port, 
                           A(30) => P_tmp_13_30_port, A(29) => P_tmp_13_29_port
                           , A(28) => P_tmp_13_28_port, A(27) => 
                           P_tmp_13_27_port, A(26) => P_tmp_13_26_port, A(25) 
                           => P_tmp_13_25_port, A(24) => P_tmp_13_24_port, 
                           A(23) => P_tmp_13_23_port, A(22) => P_tmp_13_22_port
                           , A(21) => P_tmp_13_21_port, A(20) => 
                           P_tmp_13_20_port, A(19) => P_tmp_13_19_port, A(18) 
                           => P_tmp_13_18_port, A(17) => P_tmp_13_17_port, 
                           A(16) => P_tmp_13_16_port, A(15) => P_tmp_13_15_port
                           , A(14) => P_tmp_13_14_port, A(13) => 
                           P_tmp_13_13_port, A(12) => P_tmp_13_12_port, A(11) 
                           => P_tmp_13_11_port, A(10) => P_tmp_13_10_port, A(9)
                           => P_tmp_13_9_port, A(8) => P_tmp_13_8_port, A(7) =>
                           P_tmp_13_7_port, A(6) => P_tmp_13_6_port, A(5) => 
                           P_tmp_13_5_port, A(4) => P_tmp_13_4_port, A(3) => 
                           P_tmp_13_3_port, A(2) => P_tmp_13_2_port, A(1) => 
                           P_tmp_13_1_port, A(0) => P_tmp_13_0_port, B(63) => 
                           OUT_MUX_14_63_port, B(62) => OUT_MUX_14_62_port, 
                           B(61) => OUT_MUX_14_61_port, B(60) => 
                           OUT_MUX_14_60_port, B(59) => OUT_MUX_14_59_port, 
                           B(58) => OUT_MUX_14_58_port, B(57) => 
                           OUT_MUX_14_57_port, B(56) => OUT_MUX_14_56_port, 
                           B(55) => OUT_MUX_14_55_port, B(54) => 
                           OUT_MUX_14_54_port, B(53) => OUT_MUX_14_53_port, 
                           B(52) => OUT_MUX_14_52_port, B(51) => 
                           OUT_MUX_14_51_port, B(50) => OUT_MUX_14_50_port, 
                           B(49) => OUT_MUX_14_49_port, B(48) => 
                           OUT_MUX_14_48_port, B(47) => OUT_MUX_14_47_port, 
                           B(46) => OUT_MUX_14_46_port, B(45) => 
                           OUT_MUX_14_45_port, B(44) => OUT_MUX_14_44_port, 
                           B(43) => OUT_MUX_14_43_port, B(42) => 
                           OUT_MUX_14_42_port, B(41) => OUT_MUX_14_41_port, 
                           B(40) => OUT_MUX_14_40_port, B(39) => 
                           OUT_MUX_14_39_port, B(38) => OUT_MUX_14_38_port, 
                           B(37) => OUT_MUX_14_37_port, B(36) => 
                           OUT_MUX_14_36_port, B(35) => OUT_MUX_14_35_port, 
                           B(34) => OUT_MUX_14_34_port, B(33) => 
                           OUT_MUX_14_33_port, B(32) => OUT_MUX_14_32_port, 
                           B(31) => OUT_MUX_14_31_port, B(30) => 
                           OUT_MUX_14_30_port, B(29) => OUT_MUX_14_29_port, 
                           B(28) => OUT_MUX_14_28_port, B(27) => 
                           OUT_MUX_14_27_port, B(26) => OUT_MUX_14_26_port, 
                           B(25) => OUT_MUX_14_25_port, B(24) => 
                           OUT_MUX_14_24_port, B(23) => OUT_MUX_14_23_port, 
                           B(22) => OUT_MUX_14_22_port, B(21) => 
                           OUT_MUX_14_21_port, B(20) => OUT_MUX_14_20_port, 
                           B(19) => OUT_MUX_14_19_port, B(18) => 
                           OUT_MUX_14_18_port, B(17) => OUT_MUX_14_17_port, 
                           B(16) => OUT_MUX_14_16_port, B(15) => 
                           OUT_MUX_14_15_port, B(14) => OUT_MUX_14_14_port, 
                           B(13) => OUT_MUX_14_13_port, B(12) => 
                           OUT_MUX_14_12_port, B(11) => OUT_MUX_14_11_port, 
                           B(10) => OUT_MUX_14_10_port, B(9) => 
                           OUT_MUX_14_9_port, B(8) => OUT_MUX_14_8_port, B(7) 
                           => OUT_MUX_14_7_port, B(6) => OUT_MUX_14_6_port, 
                           B(5) => OUT_MUX_14_5_port, B(4) => OUT_MUX_14_4_port
                           , B(3) => OUT_MUX_14_3_port, B(2) => 
                           OUT_MUX_14_2_port, B(1) => OUT_MUX_14_1_port, B(0) 
                           => OUT_MUX_14_0_port, Ci => X_Logic0_port, S(63) => 
                           P_tmp_14_63_port, S(62) => P_tmp_14_62_port, S(61) 
                           => P_tmp_14_61_port, S(60) => P_tmp_14_60_port, 
                           S(59) => P_tmp_14_59_port, S(58) => P_tmp_14_58_port
                           , S(57) => P_tmp_14_57_port, S(56) => 
                           P_tmp_14_56_port, S(55) => P_tmp_14_55_port, S(54) 
                           => P_tmp_14_54_port, S(53) => P_tmp_14_53_port, 
                           S(52) => P_tmp_14_52_port, S(51) => P_tmp_14_51_port
                           , S(50) => P_tmp_14_50_port, S(49) => 
                           P_tmp_14_49_port, S(48) => P_tmp_14_48_port, S(47) 
                           => P_tmp_14_47_port, S(46) => P_tmp_14_46_port, 
                           S(45) => P_tmp_14_45_port, S(44) => P_tmp_14_44_port
                           , S(43) => P_tmp_14_43_port, S(42) => 
                           P_tmp_14_42_port, S(41) => P_tmp_14_41_port, S(40) 
                           => P_tmp_14_40_port, S(39) => P_tmp_14_39_port, 
                           S(38) => P_tmp_14_38_port, S(37) => P_tmp_14_37_port
                           , S(36) => P_tmp_14_36_port, S(35) => 
                           P_tmp_14_35_port, S(34) => P_tmp_14_34_port, S(33) 
                           => P_tmp_14_33_port, S(32) => P_tmp_14_32_port, 
                           S(31) => P_tmp_14_31_port, S(30) => P_tmp_14_30_port
                           , S(29) => P_tmp_14_29_port, S(28) => 
                           P_tmp_14_28_port, S(27) => P_tmp_14_27_port, S(26) 
                           => P_tmp_14_26_port, S(25) => P_tmp_14_25_port, 
                           S(24) => P_tmp_14_24_port, S(23) => P_tmp_14_23_port
                           , S(22) => P_tmp_14_22_port, S(21) => 
                           P_tmp_14_21_port, S(20) => P_tmp_14_20_port, S(19) 
                           => P_tmp_14_19_port, S(18) => P_tmp_14_18_port, 
                           S(17) => P_tmp_14_17_port, S(16) => P_tmp_14_16_port
                           , S(15) => P_tmp_14_15_port, S(14) => 
                           P_tmp_14_14_port, S(13) => P_tmp_14_13_port, S(12) 
                           => P_tmp_14_12_port, S(11) => P_tmp_14_11_port, 
                           S(10) => P_tmp_14_10_port, S(9) => P_tmp_14_9_port, 
                           S(8) => P_tmp_14_8_port, S(7) => P_tmp_14_7_port, 
                           S(6) => P_tmp_14_6_port, S(5) => P_tmp_14_5_port, 
                           S(4) => P_tmp_14_4_port, S(3) => P_tmp_14_3_port, 
                           S(2) => P_tmp_14_2_port, S(1) => P_tmp_14_1_port, 
                           S(0) => P_tmp_14_0_port, Co => n_1293);
   RCAi_14 : RCA_NBIT64_1 port map( A(63) => P_tmp_14_63_port, A(62) => 
                           P_tmp_14_62_port, A(61) => P_tmp_14_61_port, A(60) 
                           => P_tmp_14_60_port, A(59) => P_tmp_14_59_port, 
                           A(58) => P_tmp_14_58_port, A(57) => P_tmp_14_57_port
                           , A(56) => P_tmp_14_56_port, A(55) => 
                           P_tmp_14_55_port, A(54) => P_tmp_14_54_port, A(53) 
                           => P_tmp_14_53_port, A(52) => P_tmp_14_52_port, 
                           A(51) => P_tmp_14_51_port, A(50) => P_tmp_14_50_port
                           , A(49) => P_tmp_14_49_port, A(48) => 
                           P_tmp_14_48_port, A(47) => P_tmp_14_47_port, A(46) 
                           => P_tmp_14_46_port, A(45) => P_tmp_14_45_port, 
                           A(44) => P_tmp_14_44_port, A(43) => P_tmp_14_43_port
                           , A(42) => P_tmp_14_42_port, A(41) => 
                           P_tmp_14_41_port, A(40) => P_tmp_14_40_port, A(39) 
                           => P_tmp_14_39_port, A(38) => P_tmp_14_38_port, 
                           A(37) => P_tmp_14_37_port, A(36) => P_tmp_14_36_port
                           , A(35) => P_tmp_14_35_port, A(34) => 
                           P_tmp_14_34_port, A(33) => P_tmp_14_33_port, A(32) 
                           => P_tmp_14_32_port, A(31) => P_tmp_14_31_port, 
                           A(30) => P_tmp_14_30_port, A(29) => P_tmp_14_29_port
                           , A(28) => P_tmp_14_28_port, A(27) => 
                           P_tmp_14_27_port, A(26) => P_tmp_14_26_port, A(25) 
                           => P_tmp_14_25_port, A(24) => P_tmp_14_24_port, 
                           A(23) => P_tmp_14_23_port, A(22) => P_tmp_14_22_port
                           , A(21) => P_tmp_14_21_port, A(20) => 
                           P_tmp_14_20_port, A(19) => P_tmp_14_19_port, A(18) 
                           => P_tmp_14_18_port, A(17) => P_tmp_14_17_port, 
                           A(16) => P_tmp_14_16_port, A(15) => P_tmp_14_15_port
                           , A(14) => P_tmp_14_14_port, A(13) => 
                           P_tmp_14_13_port, A(12) => P_tmp_14_12_port, A(11) 
                           => P_tmp_14_11_port, A(10) => P_tmp_14_10_port, A(9)
                           => P_tmp_14_9_port, A(8) => P_tmp_14_8_port, A(7) =>
                           P_tmp_14_7_port, A(6) => P_tmp_14_6_port, A(5) => 
                           P_tmp_14_5_port, A(4) => P_tmp_14_4_port, A(3) => 
                           P_tmp_14_3_port, A(2) => P_tmp_14_2_port, A(1) => 
                           P_tmp_14_1_port, A(0) => P_tmp_14_0_port, B(63) => 
                           OUT_MUX_15_63_port, B(62) => OUT_MUX_15_62_port, 
                           B(61) => OUT_MUX_15_61_port, B(60) => 
                           OUT_MUX_15_60_port, B(59) => OUT_MUX_15_59_port, 
                           B(58) => OUT_MUX_15_58_port, B(57) => 
                           OUT_MUX_15_57_port, B(56) => OUT_MUX_15_56_port, 
                           B(55) => OUT_MUX_15_55_port, B(54) => 
                           OUT_MUX_15_54_port, B(53) => OUT_MUX_15_53_port, 
                           B(52) => OUT_MUX_15_52_port, B(51) => 
                           OUT_MUX_15_51_port, B(50) => OUT_MUX_15_50_port, 
                           B(49) => OUT_MUX_15_49_port, B(48) => 
                           OUT_MUX_15_48_port, B(47) => OUT_MUX_15_47_port, 
                           B(46) => OUT_MUX_15_46_port, B(45) => 
                           OUT_MUX_15_45_port, B(44) => OUT_MUX_15_44_port, 
                           B(43) => OUT_MUX_15_43_port, B(42) => 
                           OUT_MUX_15_42_port, B(41) => OUT_MUX_15_41_port, 
                           B(40) => OUT_MUX_15_40_port, B(39) => 
                           OUT_MUX_15_39_port, B(38) => OUT_MUX_15_38_port, 
                           B(37) => OUT_MUX_15_37_port, B(36) => 
                           OUT_MUX_15_36_port, B(35) => OUT_MUX_15_35_port, 
                           B(34) => OUT_MUX_15_34_port, B(33) => 
                           OUT_MUX_15_33_port, B(32) => OUT_MUX_15_32_port, 
                           B(31) => OUT_MUX_15_31_port, B(30) => 
                           OUT_MUX_15_30_port, B(29) => OUT_MUX_15_29_port, 
                           B(28) => OUT_MUX_15_28_port, B(27) => 
                           OUT_MUX_15_27_port, B(26) => OUT_MUX_15_26_port, 
                           B(25) => OUT_MUX_15_25_port, B(24) => 
                           OUT_MUX_15_24_port, B(23) => OUT_MUX_15_23_port, 
                           B(22) => OUT_MUX_15_22_port, B(21) => 
                           OUT_MUX_15_21_port, B(20) => OUT_MUX_15_20_port, 
                           B(19) => OUT_MUX_15_19_port, B(18) => 
                           OUT_MUX_15_18_port, B(17) => OUT_MUX_15_17_port, 
                           B(16) => OUT_MUX_15_16_port, B(15) => 
                           OUT_MUX_15_15_port, B(14) => OUT_MUX_15_14_port, 
                           B(13) => OUT_MUX_15_13_port, B(12) => 
                           OUT_MUX_15_12_port, B(11) => OUT_MUX_15_11_port, 
                           B(10) => OUT_MUX_15_10_port, B(9) => 
                           OUT_MUX_15_9_port, B(8) => OUT_MUX_15_8_port, B(7) 
                           => OUT_MUX_15_7_port, B(6) => OUT_MUX_15_6_port, 
                           B(5) => OUT_MUX_15_5_port, B(4) => OUT_MUX_15_4_port
                           , B(3) => OUT_MUX_15_3_port, B(2) => 
                           OUT_MUX_15_2_port, B(1) => OUT_MUX_15_1_port, B(0) 
                           => OUT_MUX_15_0_port, Ci => X_Logic0_port, S(63) => 
                           P(63), S(62) => P(62), S(61) => P(61), S(60) => 
                           P(60), S(59) => P(59), S(58) => P(58), S(57) => 
                           P(57), S(56) => P(56), S(55) => P(55), S(54) => 
                           P(54), S(53) => P(53), S(52) => P(52), S(51) => 
                           P(51), S(50) => P(50), S(49) => P(49), S(48) => 
                           P(48), S(47) => P(47), S(46) => P(46), S(45) => 
                           P(45), S(44) => P(44), S(43) => P(43), S(42) => 
                           P(42), S(41) => P(41), S(40) => P(40), S(39) => 
                           P(39), S(38) => P(38), S(37) => P(37), S(36) => 
                           P(36), S(35) => P(35), S(34) => P(34), S(33) => 
                           P(33), S(32) => P(32), S(31) => P(31), S(30) => 
                           P(30), S(29) => P(29), S(28) => P(28), S(27) => 
                           P(27), S(26) => P(26), S(25) => P(25), S(24) => 
                           P(24), S(23) => P(23), S(22) => P(22), S(21) => 
                           P(21), S(20) => P(20), S(19) => P(19), S(18) => 
                           P(18), S(17) => P(17), S(16) => P(16), S(15) => 
                           P(15), S(14) => P(14), S(13) => P(13), S(12) => 
                           P(12), S(11) => P(11), S(10) => P(10), S(9) => P(9),
                           S(8) => P(8), S(7) => P(7), S(6) => P(6), S(5) => 
                           P(5), S(4) => P(4), S(3) => P(3), S(2) => P(2), S(1)
                           => P(1), S(0) => P(0), Co => n_1294);
   add_88 : BOOTHMUL_DW01_inc_0 port map( A(31) => n235, A(30) => n229, A(29) 
                           => n166, A(28) => n156, A(27) => n223, A(26) => n221
                           , A(25) => n179, A(24) => n154, A(23) => n145, A(22)
                           => n144, A(21) => n140, A(20) => net15411, A(19) => 
                           net15417, A(18) => n147, A(17) => n141, A(16) => 
                           net15435, A(15) => net15441, A(14) => net15447, 
                           A(13) => net15453, A(12) => net17026, A(11) => n158,
                           A(10) => net18009, A(9) => net15477, A(8) => 
                           net15483, A(7) => n165, A(6) => net15495, A(5) => 
                           n181, A(4) => n189, A(3) => n180, A(2) => n184, A(1)
                           => net15525, A(0) => net15535, SUM(31) => N97, 
                           SUM(30) => N96, SUM(29) => N95, SUM(28) => N94, 
                           SUM(27) => N93, SUM(26) => N92, SUM(25) => N91, 
                           SUM(24) => N90, SUM(23) => N89, SUM(22) => N88, 
                           SUM(21) => N87, SUM(20) => N86, SUM(19) => N85, 
                           SUM(18) => N84, SUM(17) => N83, SUM(16) => N82, 
                           SUM(15) => N81, SUM(14) => N80, SUM(13) => N79, 
                           SUM(12) => N78, SUM(11) => N77, SUM(10) => N76, 
                           SUM(9) => N75, SUM(8) => N74, SUM(7) => N73, SUM(6) 
                           => N72, SUM(5) => N71, SUM(4) => N70, SUM(3) => N69,
                           SUM(2) => N68, SUM(1) => N67, SUM(0) => N66);
   U155 : BUF_X4 port map( A => net15837, Z => net25715);
   U156 : BUF_X1 port map( A => net17729, Z => net15837);
   U157 : INV_X1 port map( A => A(27), ZN => n138);
   U158 : AND4_X2 port map( A1 => n235, A2 => n211, A3 => n213, A4 => n215, ZN 
                           => n139);
   U159 : AND4_X1 port map( A1 => n235, A2 => n211, A3 => n213, A4 => n215, ZN 
                           => net17036);
   U160 : INV_X1 port map( A => net15403, ZN => n140);
   U161 : INV_X1 port map( A => net15427, ZN => n141);
   U162 : CLKBUF_X1 port map( A => A_neg_tmp_1_port, Z => n142);
   U255 : BUF_X1 port map( A => net17729, Z => n143);
   U256 : INV_X2 port map( A => A(3), ZN => n180);
   U257 : INV_X2 port map( A => A(2), ZN => n184);
   U258 : AND4_X1 port map( A1 => n217, A2 => n219, A3 => n191, A4 => n192, ZN 
                           => net17038);
   U259 : AND2_X2 port map( A1 => N71, A2 => net25715, ZN => n186);
   U260 : AND2_X2 port map( A1 => net17729, A2 => N68, ZN => n178);
   U261 : AND2_X2 port map( A1 => N76, A2 => net25715, ZN => A_neg_tmp_10_port)
                           ;
   U262 : BUF_X4 port map( A => A_neg_tmp_63_port, Z => n199);
   U263 : AND2_X4 port map( A1 => N74, A2 => net25715, ZN => A_neg_tmp_8_port);
   U264 : INV_X1 port map( A => A(28), ZN => n156);
   U265 : AND2_X2 port map( A1 => N77, A2 => net25715, ZN => A_neg_tmp_11_port)
                           ;
   U266 : INV_X2 port map( A => n234, ZN => n233);
   U267 : INV_X1 port map( A => A(28), ZN => n225);
   U268 : AND4_X2 port map( A1 => net17613, A2 => net17614, A3 => net17616, A4 
                           => n174, ZN => n128);
   U269 : AND4_X2 port map( A1 => n169, A2 => n170, A3 => n171, A4 => n172, ZN 
                           => n174);
   U270 : INV_X1 port map( A => net15397, ZN => n144);
   U271 : INV_X1 port map( A => net15391, ZN => n145);
   U272 : INV_X1 port map( A => A(0), ZN => n146);
   U273 : AND2_X2 port map( A1 => N70, A2 => n143, ZN => n194);
   U274 : INV_X1 port map( A => net15421, ZN => n147);
   U275 : AND4_X1 port map( A1 => n225, A2 => n227, A3 => n209, A4 => n190, ZN 
                           => n148);
   U276 : AND4_X1 port map( A1 => n225, A2 => n227, A3 => n209, A4 => n190, ZN 
                           => net18025);
   U277 : AND2_X1 port map( A1 => n152, A2 => n149, ZN => n157);
   U278 : NOR2_X1 port map( A1 => A(19), A2 => A(1), ZN => n149);
   U279 : INV_X1 port map( A => A(29), ZN => n150);
   U280 : INV_X1 port map( A => A(29), ZN => n166);
   U281 : NOR4_X1 port map( A1 => A(20), A2 => A(21), A3 => A(22), A4 => A(23),
                           ZN => n153);
   U282 : INV_X1 port map( A => A(20), ZN => net15411);
   U283 : INV_X1 port map( A => A(21), ZN => net15405);
   U284 : INV_X1 port map( A => A(22), ZN => net15399);
   U285 : INV_X1 port map( A => A(23), ZN => net15393);
   U286 : AND2_X1 port map( A1 => N72, A2 => n143, ZN => A_neg_tmp_6_port);
   U287 : INV_X1 port map( A => A(10), ZN => n151);
   U288 : INV_X1 port map( A => A(29), ZN => n227);
   U289 : NOR2_X1 port map( A1 => A(17), A2 => A(18), ZN => n152);
   U290 : AND4_X1 port map( A1 => net15411, A2 => net15405, A3 => net15399, A4 
                           => net15393, ZN => net17613);
   U291 : INV_X1 port map( A => A(17), ZN => net15429);
   U292 : INV_X1 port map( A => A(24), ZN => n154);
   U293 : INV_X1 port map( A => A(24), ZN => n217);
   U294 : AND4_X1 port map( A1 => n217, A2 => n219, A3 => n191, A4 => n138, ZN 
                           => net98228);
   U295 : INV_X1 port map( A => A(3), ZN => n155);
   U296 : AND4_X1 port map( A1 => net15429, A2 => net15525, A3 => n175, A4 => 
                           net15423, ZN => net17614);
   U297 : INV_X1 port map( A => A(18), ZN => net15423);
   U298 : INV_X1 port map( A => A(11), ZN => n158);
   U299 : AND4_X2 port map( A1 => n161, A2 => n139, A3 => n148, A4 => net17038,
                           ZN => net18732);
   U300 : AND4_X2 port map( A1 => net17036, A2 => net18025, A3 => net98228, A4 
                           => n161, ZN => n129);
   U301 : INV_X1 port map( A => A(4), ZN => n159);
   U302 : INV_X1 port map( A => A(5), ZN => n160);
   U303 : AND2_X1 port map( A1 => n162, A2 => n163, ZN => n161);
   U304 : NOR2_X1 port map( A1 => A(8), A2 => A(9), ZN => n163);
   U305 : NOR2_X1 port map( A1 => A(6), A2 => A(7), ZN => n162);
   U306 : INV_X1 port map( A => A(8), ZN => net15483);
   U307 : INV_X1 port map( A => A(9), ZN => net15477);
   U308 : INV_X1 port map( A => net15495, ZN => net15493);
   U309 : INV_X1 port map( A => A(7), ZN => net15489);
   U310 : INV_X1 port map( A => A(7), ZN => n165);
   U311 : INV_X1 port map( A => A(6), ZN => net15495);
   U312 : NAND2_X1 port map( A1 => n167, A2 => net18732, ZN => n164);
   U313 : INV_X1 port map( A => net15483, ZN => net15481);
   U314 : AND4_X2 port map( A1 => n153, A2 => n157, A3 => net17616, A4 => n174,
                           ZN => n167);
   U315 : AND4_X2 port map( A1 => n176, A2 => net15471, A3 => net15465, A4 => 
                           n173, ZN => net17616);
   U316 : AND2_X2 port map( A1 => n127, A2 => N66, ZN => A_neg_tmp_0_port);
   U317 : AOI21_X2 port map( B1 => n128, B2 => n129, A => n168, ZN => 
                           A_neg_tmp_1_port);
   U318 : INV_X1 port map( A => N67, ZN => n168);
   U319 : INV_X1 port map( A => A(13), ZN => n169);
   U320 : INV_X1 port map( A => A(14), ZN => n170);
   U321 : INV_X1 port map( A => A(15), ZN => n171);
   U322 : INV_X1 port map( A => A(16), ZN => n172);
   U323 : NAND2_X1 port map( A1 => n167, A2 => net18732, ZN => net17729);
   U324 : NAND2_X1 port map( A1 => n167, A2 => net18016, ZN => n127);
   U325 : INV_X1 port map( A => A(12), ZN => n173);
   U326 : INV_X1 port map( A => A(11), ZN => net15465);
   U327 : INV_X1 port map( A => A(10), ZN => net15471);
   U328 : INV_X1 port map( A => A(0), ZN => n176);
   U329 : INV_X1 port map( A => n146, ZN => net15533);
   U330 : INV_X1 port map( A => A(1), ZN => net15525);
   U331 : INV_X1 port map( A => A(19), ZN => n175);
   U332 : INV_X1 port map( A => net15423, ZN => net15421);
   U333 : INV_X1 port map( A => net15429, ZN => net15427);
   U334 : INV_X1 port map( A => net15393, ZN => net15391);
   U335 : INV_X1 port map( A => net15399, ZN => net15397);
   U336 : INV_X1 port map( A => net15405, ZN => net15403);
   U337 : INV_X1 port map( A => net15411, ZN => net15409);
   U338 : INV_X1 port map( A => A(13), ZN => net15453);
   U339 : INV_X1 port map( A => A(14), ZN => net15447);
   U340 : INV_X1 port map( A => A(15), ZN => net15441);
   U341 : INV_X1 port map( A => A(16), ZN => net15435);
   U342 : CLKBUF_X3 port map( A => A_neg_tmp_7_port, Z => n177);
   U343 : AND2_X1 port map( A1 => N73, A2 => net25715, ZN => A_neg_tmp_7_port);
   U344 : INV_X2 port map( A => net15489, ZN => net15487);
   U345 : INV_X1 port map( A => A(25), ZN => n179);
   U346 : INV_X1 port map( A => A(25), ZN => n219);
   U347 : INV_X1 port map( A => A(3), ZN => n211);
   U348 : INV_X1 port map( A => A(5), ZN => n181);
   U349 : INV_X1 port map( A => A(5), ZN => n215);
   U350 : CLKBUF_X3 port map( A => A_neg_tmp_9_port, Z => n182);
   U351 : AND2_X2 port map( A1 => N69, A2 => n143, ZN => n188);
   U352 : AND2_X1 port map( A1 => N71, A2 => n143, ZN => A_neg_tmp_5_port);
   U353 : INV_X1 port map( A => A(2), ZN => n183);
   U354 : INV_X1 port map( A => A(2), ZN => n209);
   U355 : AND2_X2 port map( A1 => N72, A2 => net25715, ZN => n185);
   U356 : BUF_X2 port map( A => A_neg_shifted_by2_0_2_port, Z => n187);
   U357 : AND2_X1 port map( A1 => n164, A2 => N68, ZN => A_neg_tmp_2_port);
   U358 : AND2_X1 port map( A1 => net17729, A2 => N69, ZN => A_neg_tmp_3_port);
   U359 : AND4_X1 port map( A1 => n156, A2 => n150, A3 => n183, A4 => n229, ZN 
                           => n195);
   U360 : INV_X1 port map( A => A(4), ZN => n189);
   U361 : INV_X1 port map( A => A(4), ZN => n213);
   U362 : INV_X1 port map( A => A(19), ZN => net15417);
   U363 : AND4_X1 port map( A1 => n139, A2 => n161, A3 => n195, A4 => net17038,
                           ZN => net18016);
   U364 : INV_X1 port map( A => A(30), ZN => n190);
   U365 : INV_X1 port map( A => A(10), ZN => net18009);
   U366 : INV_X1 port map( A => A(1), ZN => net18006);
   U367 : INV_X1 port map( A => A(26), ZN => n191);
   U368 : INV_X1 port map( A => n183, ZN => n208);
   U369 : INV_X1 port map( A => A(27), ZN => n192);
   U370 : BUF_X2 port map( A => B(1), Z => n193);
   U371 : AND2_X1 port map( A1 => N70, A2 => net15837, ZN => A_neg_tmp_4_port);
   U372 : BUF_X1 port map( A => A_neg_shifted_by2_5_47_port, Z => n203);
   U373 : BUF_X1 port map( A => A_neg_shifted_by2_3_47_port, Z => n205);
   U374 : BUF_X1 port map( A => A_neg_shifted_by2_4_47_port, Z => n204);
   U375 : BUF_X1 port map( A => A_neg_shifted_by2_6_47_port, Z => n202);
   U376 : BUF_X1 port map( A => A_neg_shifted_by2_0_47_port, Z => n207);
   U377 : BUF_X1 port map( A => A_neg_shifted_by2_1_47_port, Z => n206);
   U378 : AND2_X1 port map( A1 => N75, A2 => net25715, ZN => A_neg_tmp_9_port);
   U379 : AND2_X1 port map( A1 => N78, A2 => net25715, ZN => A_neg_tmp_12_port)
                           ;
   U380 : AND2_X1 port map( A1 => N79, A2 => net25715, ZN => A_neg_tmp_13_port)
                           ;
   U381 : AND2_X1 port map( A1 => N80, A2 => net25715, ZN => A_neg_tmp_14_port)
                           ;
   U382 : AND2_X1 port map( A1 => N81, A2 => net25715, ZN => A_neg_tmp_15_port)
                           ;
   U383 : AND2_X1 port map( A1 => N82, A2 => net25715, ZN => A_neg_tmp_16_port)
                           ;
   U384 : AND2_X1 port map( A1 => N83, A2 => net25715, ZN => A_neg_tmp_17_port)
                           ;
   U385 : AND2_X1 port map( A1 => N96, A2 => net25715, ZN => A_neg_tmp_30_port)
                           ;
   U386 : AND2_X1 port map( A1 => N95, A2 => net25715, ZN => A_neg_tmp_29_port)
                           ;
   U387 : AND2_X1 port map( A1 => N94, A2 => net25715, ZN => A_neg_tmp_28_port)
                           ;
   U388 : AND2_X1 port map( A1 => N93, A2 => net25715, ZN => A_neg_tmp_27_port)
                           ;
   U389 : AND2_X1 port map( A1 => N92, A2 => net25715, ZN => A_neg_tmp_26_port)
                           ;
   U390 : AND2_X1 port map( A1 => N91, A2 => net25715, ZN => A_neg_tmp_25_port)
                           ;
   U391 : AND2_X1 port map( A1 => N90, A2 => net25715, ZN => A_neg_tmp_24_port)
                           ;
   U392 : AND2_X1 port map( A1 => N89, A2 => net25715, ZN => A_neg_tmp_23_port)
                           ;
   U393 : AND2_X1 port map( A1 => N88, A2 => net25715, ZN => A_neg_tmp_22_port)
                           ;
   U394 : AND2_X1 port map( A1 => N84, A2 => net25715, ZN => A_neg_tmp_18_port)
                           ;
   U395 : AND2_X1 port map( A1 => N87, A2 => net25715, ZN => A_neg_tmp_21_port)
                           ;
   U396 : AND2_X1 port map( A1 => N85, A2 => net25715, ZN => A_neg_tmp_19_port)
                           ;
   U397 : AND2_X1 port map( A1 => N86, A2 => net25715, ZN => A_neg_tmp_20_port)
                           ;
   U398 : BUF_X2 port map( A => A_neg_tmp_63_port, Z => n197);
   U399 : BUF_X2 port map( A => A_neg_tmp_63_port, Z => n198);
   U400 : BUF_X2 port map( A => A_neg_tmp_63_port, Z => n196);
   U401 : BUF_X2 port map( A => A_neg_tmp_63_port, Z => n200);
   U402 : BUF_X1 port map( A => A_neg_tmp_63_port, Z => n201);
   U403 : BUF_X1 port map( A => A_pos_shifted_by2_0_47_port, Z => n242);
   U404 : BUF_X1 port map( A => A_pos_shifted_by2_1_47_port, Z => n241);
   U405 : BUF_X1 port map( A => A_pos_shifted_by2_2_47_port, Z => n240);
   U406 : BUF_X1 port map( A => A_pos_shifted_by2_4_47_port, Z => n238);
   U407 : BUF_X1 port map( A => A_pos_shifted_by2_6_47_port, Z => n236);
   U408 : BUF_X1 port map( A => A_pos_shifted_by2_5_47_port, Z => n237);
   U409 : BUF_X1 port map( A => A_pos_shifted_by2_3_47_port, Z => n239);
   U410 : INV_X1 port map( A => net15477, ZN => net15475);
   U411 : INV_X1 port map( A => net15453, ZN => net15451);
   U412 : INV_X1 port map( A => net15447, ZN => net15445);
   U413 : INV_X1 port map( A => net15417, ZN => net15415);
   U414 : INV_X1 port map( A => n154, ZN => n216);
   U415 : INV_X1 port map( A => n179, ZN => n218);
   U416 : INV_X1 port map( A => n160, ZN => n214);
   U417 : AND2_X1 port map( A1 => N97, A2 => net25715, ZN => A_neg_tmp_31_port)
                           ;
   U418 : INV_X1 port map( A => n156, ZN => n224);
   U419 : INV_X1 port map( A => n150, ZN => n226);
   U420 : INV_X1 port map( A => A(0), ZN => net15535);
   U421 : INV_X1 port map( A => A(31), ZN => n235);
   U422 : INV_X1 port map( A => A(31), ZN => n234);
   U423 : INV_X1 port map( A => net15441, ZN => net15439);
   U424 : INV_X1 port map( A => net15435, ZN => net15433);
   U425 : INV_X1 port map( A => n151, ZN => net15469);
   U426 : INV_X1 port map( A => n229, ZN => n228);
   U427 : INV_X1 port map( A => n221, ZN => n220);
   U428 : INV_X1 port map( A => A(26), ZN => n221);
   U429 : INV_X1 port map( A => A(12), ZN => net17026);
   U430 : AND2_X1 port map( A1 => n234, A2 => net25715, ZN => A_neg_tmp_63_port
                           );
   U431 : INV_X1 port map( A => n223, ZN => n222);
   U432 : INV_X1 port map( A => A(30), ZN => n229);
   U433 : INV_X1 port map( A => A(27), ZN => n223);
   U434 : INV_X2 port map( A => net18006, ZN => net15523);
   U435 : INV_X2 port map( A => n155, ZN => n210);
   U436 : INV_X2 port map( A => n159, ZN => n212);
   U437 : INV_X2 port map( A => n158, ZN => net15463);
   U438 : INV_X2 port map( A => net17026, ZN => net15457);
   U439 : INV_X4 port map( A => n234, ZN => n230);
   U440 : INV_X4 port map( A => n234, ZN => n231);
   U441 : INV_X4 port map( A => n234, ZN => n232);

end SYN_STRUCTURAL;
