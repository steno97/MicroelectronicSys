
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file;

architecture SYN_A of register_file is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n4254, 
      n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
      n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, 
      n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, 
      n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, 
      n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
      n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, 
      n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, 
      n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, 
      n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
      n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, 
      n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
      n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
      n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, 
      n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, 
      n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
      n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
      n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, 
      n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, 
      n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
      n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
      n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, 
      n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, 
      n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
      n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
      n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, 
      n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, 
      n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, 
      n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
      n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, 
      n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, 
      n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, 
      n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, 
      n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, 
      n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, 
      n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, 
      n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, 
      n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, 
      n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, 
      n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, 
      n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, 
      n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, 
      n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, 
      n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, 
      n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, 
      n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, 
      n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, 
      n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, 
      n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, 
      n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, 
      n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, 
      n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, 
      n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, 
      n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, 
      n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, 
      n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, 
      n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, 
      n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, 
      n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, 
      n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, 
      n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, 
      n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, 
      n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, 
      n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
      n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, 
      n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
      n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, 
      n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, 
      n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, 
      n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, 
      n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, 
      n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, 
      n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, 
      n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, 
      n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, 
      n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, 
      n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, 
      n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, 
      n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, 
      n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, 
      n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, 
      n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, 
      n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, 
      n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, 
      n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, 
      n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, 
      n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, 
      n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, 
      n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, 
      n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, 
      n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, 
      n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, 
      n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, 
      n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, 
      n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, 
      n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, 
      n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
      n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, 
      n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, 
      n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, 
      n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
      n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, 
      n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, 
      n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
      n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
      n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, 
      n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, 
      n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, 
      n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, 
      n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, 
      n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, 
      n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
      n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, 
      n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, 
      n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, 
      n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, 
      n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, 
      n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, 
      n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, 
      n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, 
      n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
      n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, 
      n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, 
      n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
      n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, 
      n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, 
      n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, 
      n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, 
      n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, 
      n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, 
      n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, 
      n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
      n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, 
      n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, 
      n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, 
      n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, 
      n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, 
      n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, 
      n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
      n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, 
      n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, 
      n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, 
      n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, 
      n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, 
      n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, 
      n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, 
      n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, 
      n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, 
      n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, 
      n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, 
      n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, 
      n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, 
      n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, 
      n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, 
      n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, 
      n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, 
      n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, 
      n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, 
      n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, 
      n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
      n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, 
      n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, 
      n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, 
      n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, 
      n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, 
      n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, 
      n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, 
      n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, 
      n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, 
      n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, 
      n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, 
      n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, 
      n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, 
      n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, 
      n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, 
      n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
      n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, 
      n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, 
      n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, 
      n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, 
      n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, 
      n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, 
      n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, 
      n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, 
      n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, 
      n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, 
      n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, 
      n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, 
      n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, 
      n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, 
      n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, 
      n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, 
      n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, 
      n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, 
      n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, 
      n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, 
      n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, 
      n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, 
      n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, 
      n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, 
      n6415, n6416, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, 
      n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6465, n6466, 
      n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, 
      n6477, n6478, n6479, n6480, n6497, n6498, n6499, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, 
      n6539, n6540, n6541, n6542, n6543, n6544, n6593, n6594, n6595, n6596, 
      n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, 
      n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, 
      n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, 
      n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, 
      n6637, n6638, n6639, n6640, n6689, n6690, n6691, n6692, n6693, n6694, 
      n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, 
      n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, 
      n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, 
      n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, 
      n6735, n6736, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, 
      n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, 
      n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, 
      n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, 
      n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, 
      n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, 
      n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, 
      n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, 
      n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, 
      n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, 
      n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, 
      n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, 
      n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, 
      n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, 
      n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, 
      n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, 
      n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, 
      n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, 
      n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, 
      n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, 
      n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, 
      n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, 
      n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, 
      n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, 
      n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, 
      n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, 
      n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, 
      n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, 
      n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, 
      n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, 
      n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, 
      n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, 
      n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, 
      n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, 
      n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, 
      n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, 
      n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, 
      n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, 
      n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, 
      n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, 
      n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, 
      n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, 
      n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, 
      n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, 
      n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, 
      n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, 
      n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, 
      n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, 
      n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, 
      n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, 
      n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, 
      n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, 
      n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, 
      n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, 
      n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, 
      n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, 
      n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, 
      n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, 
      n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, 
      n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, 
      n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, 
      n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, 
      n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, 
      n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, 
      n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, 
      n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, 
      n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, 
      n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, 
      n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, 
      n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, 
      n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, 
      n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, 
      n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, 
      n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, 
      n7581, n7582, n7583, n7584, n7585, n7586, n7587, n_1000, n_1001, n_1002, 
      n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, 
      n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, 
      n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, 
      n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, 
      n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, 
      n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, 
      n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, 
      n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, 
      n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, 
      n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, 
      n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, 
      n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, 
      n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, 
      n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, 
      n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, 
      n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, 
      n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, 
      n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, 
      n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, 
      n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, 
      n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, 
      n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, 
      n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, 
      n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, 
      n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, 
      n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, 
      n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, 
      n_1507, n_1508, n_1509, n_1510, n_1511 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3615, CK => CLK, Q => 
                           n_1000, QN => n1);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => 
                           n_1001, QN => n2);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n_1002, QN => n3);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n_1003, QN => n4);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n_1004, QN => n5);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n_1005, QN => n6);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n_1006, QN => n7);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n_1007, QN => n8);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n_1008, QN => n9);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n_1009, QN => n10);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n_1010, QN => n11);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n_1011, QN => n12);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n_1012, QN => n13);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n_1013, QN => n14);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n_1014, QN => n15);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           n_1015, QN => n16);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           n_1016, QN => n17);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           n_1017, QN => n18);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           n_1018, QN => n19);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           n_1019, QN => n20);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           n_1020, QN => n21);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           n_1021, QN => n22);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => n_1022
                           , QN => n23);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n_1023
                           , QN => n24);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n_1024
                           , QN => n25);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n_1025
                           , QN => n26);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n_1026
                           , QN => n27);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n_1027
                           , QN => n28);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n_1028
                           , QN => n29);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n_1029
                           , QN => n30);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n_1030
                           , QN => n31);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n_1031
                           , QN => n32);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => 
                           n_1032, QN => n33);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => 
                           n_1033, QN => n34);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n_1034, QN => n35);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n_1035, QN => n36);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n_1036, QN => n37);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n_1037, QN => n38);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n_1038, QN => n39);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n_1039, QN => n40);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n_1040, QN => n41);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n_1041, QN => n42);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n_1042, QN => n43);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n_1043, QN => n44);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n_1044, QN => n45);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n_1045, QN => n46);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n_1046, QN => n47);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           n_1047, QN => n48);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           n_1048, QN => n49);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           n_1049, QN => n50);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           n_1050, QN => n51);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           n_1051, QN => n52);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           n_1052, QN => n53);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           n_1053, QN => n54);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => n_1054
                           , QN => n55);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n_1055
                           , QN => n56);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n_1056
                           , QN => n57);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n_1057
                           , QN => n58);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n_1058
                           , QN => n59);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n_1059
                           , QN => n60);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n_1060
                           , QN => n61);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n_1061
                           , QN => n62);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n_1062
                           , QN => n63);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n_1063
                           , QN => n64);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => 
                           n_1064, QN => n257);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => 
                           n_1065, QN => n258);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => 
                           n_1066, QN => n259);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => 
                           n_1067, QN => n260);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => 
                           n_1068, QN => n261);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => 
                           n_1069, QN => n262);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => 
                           n_1070, QN => n263);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => 
                           n_1071, QN => n264);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => 
                           n_1072, QN => n265);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => 
                           n_1073, QN => n266);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => 
                           n_1074, QN => n267);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => 
                           n_1075, QN => n268);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => 
                           n_1076, QN => n269);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => 
                           n_1077, QN => n270);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => 
                           n_1078, QN => n271);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => 
                           n_1079, QN => n272);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => 
                           n_1080, QN => n273);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => 
                           n_1081, QN => n274);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => 
                           n_1082, QN => n275);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => 
                           n_1083, QN => n276);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => 
                           n_1084, QN => n277);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => 
                           n_1085, QN => n278);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n_1086
                           , QN => n279);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n_1087
                           , QN => n280);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n_1088
                           , QN => n281);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n_1089
                           , QN => n282);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n_1090
                           , QN => n283);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n_1091
                           , QN => n284);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n_1092
                           , QN => n285);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n_1093
                           , QN => n286);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n_1094
                           , QN => n287);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n_1095
                           , QN => n288);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => 
                           n_1096, QN => n289);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => 
                           n_1097, QN => n290);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => 
                           n_1098, QN => n291);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => 
                           n_1099, QN => n292);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => 
                           n_1100, QN => n293);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => 
                           n_1101, QN => n294);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => 
                           n_1102, QN => n295);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => 
                           n_1103, QN => n296);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => 
                           n_1104, QN => n297);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => 
                           n_1105, QN => n298);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => 
                           n_1106, QN => n299);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => 
                           n_1107, QN => n300);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => 
                           n_1108, QN => n301);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => 
                           n_1109, QN => n302);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => 
                           n_1110, QN => n303);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => 
                           n_1111, QN => n304);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => 
                           n_1112, QN => n305);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => 
                           n_1113, QN => n306);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => 
                           n_1114, QN => n307);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => 
                           n_1115, QN => n308);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => 
                           n_1116, QN => n309);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => 
                           n_1117, QN => n310);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n_1118
                           , QN => n311);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n_1119
                           , QN => n312);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n_1120
                           , QN => n313);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n_1121
                           , QN => n314);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n_1122
                           , QN => n315);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n_1123
                           , QN => n316);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n_1124
                           , QN => n317);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n_1125
                           , QN => n318);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n_1126
                           , QN => n319);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n_1127
                           , QN => n320);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => 
                           n_1128, QN => n513);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           n_1129, QN => n514);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           n_1130, QN => n515);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n_1131, QN => n516);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           n_1132, QN => n517);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n_1133, QN => n518);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           n_1134, QN => n519);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n_1135, QN => n520);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           n_1136, QN => n521);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n_1137, QN => n522);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           n_1138, QN => n523);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n_1139, QN => n524);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           n_1140, QN => n525);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n_1141, QN => n526);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           n_1142, QN => n527);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n_1143, QN => n528);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           n_1144, QN => n529);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n_1145, QN => n530);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           n_1146, QN => n531);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n_1147, QN => n532);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           n_1148, QN => n533);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n_1149, QN => n534);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           n_1150, QN => n535);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n_1151, QN => n536);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => 
                           n_1152, QN => n537);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => 
                           n_1153, QN => n538);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => 
                           n_1154, QN => n539);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => 
                           n_1155, QN => n540);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => 
                           n_1156, QN => n541);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => 
                           n_1157, QN => n542);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => 
                           n_1158, QN => n543);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => 
                           n_1159, QN => n544);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => 
                           n_1160, QN => n545);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => 
                           n_1161, QN => n546);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           n_1162, QN => n547);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n_1163, QN => n548);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           n_1164, QN => n549);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           n_1165, QN => n550);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           n_1166, QN => n551);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => 
                           n_1167, QN => n552);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           n_1168, QN => n553);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           n_1169, QN => n554);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           n_1170, QN => n555);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           n_1171, QN => n556);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           n_1172, QN => n557);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           n_1173, QN => n558);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           n_1174, QN => n559);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           n_1175, QN => n560);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           n_1176, QN => n561);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           n_1177, QN => n562);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           n_1178, QN => n563);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           n_1179, QN => n564);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           n_1180, QN => n565);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           n_1181, QN => n566);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           n_1182, QN => n567);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           n_1183, QN => n568);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => 
                           n_1184, QN => n569);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => 
                           n_1185, QN => n570);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => 
                           n_1186, QN => n571);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => 
                           n_1187, QN => n572);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => 
                           n_1188, QN => n573);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => 
                           n_1189, QN => n574);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => 
                           n_1190, QN => n575);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => 
                           n_1191, QN => n576);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n_1192, QN => n770);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n_1193, QN => n771);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n_1194, QN => n772);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n_1195, QN => n773);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n_1196, QN => n774);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n_1197, QN => n775);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n_1198, QN => n776);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n_1199, QN => n777);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n_1200, QN => n778);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n_1201, QN => n779);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n_1202, QN => n780);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n_1203, QN => n781);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n_1204, QN => n782);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n_1205, QN => n783);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n_1206, QN => n784);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n_1207, QN => n785);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n_1208, QN => n786);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n_1209, QN => n787);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n_1210, QN => n788);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n_1211, QN => n789);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n_1212, QN => n790);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n_1213, QN => n791);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => 
                           n_1214, QN => n792);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => 
                           n_1215, QN => n793);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => 
                           n_1216, QN => n794);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => 
                           n_1217, QN => n795);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => 
                           n_1218, QN => n796);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => 
                           n_1219, QN => n797);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => 
                           n_1220, QN => n798);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => 
                           n_1221, QN => n799);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => 
                           n_1222, QN => n800);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => 
                           n_1223, QN => n801);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           n_1224, QN => n802);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n_1225, QN => n803);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n_1226, QN => n804);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n_1227, QN => n805);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n_1228, QN => n806);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n_1229, QN => n807);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n_1230, QN => n808);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n_1231, QN => n809);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n_1232, QN => n810);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n_1233, QN => n811);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n_1234, QN => n812);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n_1235, QN => n813);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n_1236, QN => n814);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n_1237, QN => n815);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n_1238, QN => n816);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n_1239, QN => n817);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n_1240, QN => n818);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n_1241, QN => n819);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n_1242, QN => n820);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n_1243, QN => n821);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n_1244, QN => n822);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n_1245, QN => n823);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => 
                           n_1246, QN => n824);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => 
                           n_1247, QN => n825);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => 
                           n_1248, QN => n826);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => 
                           n_1249, QN => n827);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => 
                           n_1250, QN => n828);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => 
                           n_1251, QN => n829);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => 
                           n_1252, QN => n830);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => 
                           n_1253, QN => n831);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => 
                           n_1254, QN => n832);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => OUT2(31), QN
                           => n6992);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => OUT2(30), QN
                           => n6968);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => OUT2(29), QN
                           => n6967);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => OUT2(28), QN
                           => n6966);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => OUT2(27), QN
                           => n6965);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => OUT2(26), QN
                           => n6964);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => OUT2(25), QN
                           => n6963);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => OUT2(24), QN
                           => n6962);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => OUT2(23), QN
                           => n6961);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => OUT2(22), QN
                           => n6960);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => OUT2(21), QN
                           => n6959);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => OUT2(20), QN
                           => n6958);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => OUT2(19), QN
                           => n6957);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => OUT2(18), QN
                           => n6956);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => OUT2(17), QN
                           => n6955);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => OUT2(16), QN
                           => n6954);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => OUT2(15), QN
                           => n6953);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT2(14), QN
                           => n6952);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT2(13), QN
                           => n6951);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT2(12), QN
                           => n6950);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT2(11), QN
                           => n6949);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT2(10), QN
                           => n6948);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT2(9), QN 
                           => n6947);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT2(8), QN 
                           => n6946);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT2(7), QN 
                           => n6945);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT2(6), QN 
                           => n6944);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT2(5), QN 
                           => n6943);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2(4), QN 
                           => n6942);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2(3), QN 
                           => n6941);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2(2), QN 
                           => n6940);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2(1), QN 
                           => n6939);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(0), QN 
                           => n6938);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT1(31), QN
                           => n6929);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT1(30), QN
                           => n6991);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT1(29), QN
                           => n6990);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT1(28), QN
                           => n6989);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT1(27), QN
                           => n6988);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT1(26), QN
                           => n6987);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT1(25), QN
                           => n6986);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT1(24), QN
                           => n6985);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT1(23), QN
                           => n6984);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT1(22), QN
                           => n6983);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT1(21), QN
                           => n6982);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT1(20), QN
                           => n6981);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT1(19), QN
                           => n6980);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT1(18), QN
                           => n6979);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT1(17), QN
                           => n6978);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT1(16), QN
                           => n6977);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT1(15), QN
                           => n6976);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT1(14), QN
                           => n6975);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT1(13), QN
                           => n6974);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT1(12), QN
                           => n6973);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT1(11), QN
                           => n6972);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT1(10), QN
                           => n6971);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1(9), QN 
                           => n6970);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1(8), QN 
                           => n6969);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1(7), QN 
                           => n6937);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1(6), QN 
                           => n6936);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1(5), QN 
                           => n6935);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1(4), QN 
                           => n6934);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1(3), QN 
                           => n6933);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1(2), QN 
                           => n6932);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1(1), QN 
                           => n6931);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1(0), QN 
                           => n6930);
   U5865 : NAND3_X1 port map( A1 => n4256, A2 => n4255, A3 => n5083, ZN => 
                           n5067);
   U5866 : NAND3_X1 port map( A1 => n5083, A2 => n4255, A3 => ADD_WR(3), ZN => 
                           n5085);
   U5867 : NAND3_X1 port map( A1 => n5083, A2 => n4256, A3 => ADD_WR(4), ZN => 
                           n5094);
   U5868 : NAND3_X1 port map( A1 => n4258, A2 => n4257, A3 => n4259, ZN => 
                           n5068);
   U5869 : NAND3_X1 port map( A1 => n4258, A2 => n4257, A3 => ADD_WR(0), ZN => 
                           n5070);
   U5870 : NAND3_X1 port map( A1 => n4259, A2 => n4257, A3 => ADD_WR(1), ZN => 
                           n5072);
   U5871 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n4257, A3 => ADD_WR(1), ZN
                           => n5074);
   U5872 : NAND3_X1 port map( A1 => n4259, A2 => n4258, A3 => ADD_WR(2), ZN => 
                           n5076);
   U5873 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n4258, A3 => ADD_WR(2), ZN
                           => n5078);
   U5874 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n4259, A3 => ADD_WR(2), ZN
                           => n5080);
   U5875 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n5083, A3 => ADD_WR(4), ZN
                           => n5103);
   U5876 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n5082);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => 
                           n5002, QN => n993);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n5003, QN => n994);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n5004, QN => n995);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n5005, QN => n996);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n5006, QN => n997);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n5007, QN => n998);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           n5008, QN => n999);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           n5009, QN => n1000);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => 
                           n5010, QN => n1001);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           n5011, QN => n1002);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           n5012, QN => n1003);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n5013, QN => n1004);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => 
                           n5014, QN => n1005);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => 
                           n5015, QN => n1006);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => 
                           n5016, QN => n1007);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => 
                           n5017, QN => n1008);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => 
                           n5018, QN => n1009);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => 
                           n5019, QN => n1010);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => 
                           n5020, QN => n1011);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => 
                           n5021, QN => n1012);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => 
                           n5022, QN => n1013);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => 
                           n5023, QN => n1014);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => n5024
                           , QN => n1015);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => n5025
                           , QN => n1016);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => n5026
                           , QN => n1017);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => n5027
                           , QN => n1018);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => n5028
                           , QN => n1019);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => n5029
                           , QN => n1020);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => n5030
                           , QN => n1021);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => n5031
                           , QN => n1022);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => n5032
                           , QN => n1023);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => n5033
                           , QN => n1024);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => 
                           n4970, QN => n961);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => 
                           n4971, QN => n962);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           n4972, QN => n963);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           n4973, QN => n964);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           n4974, QN => n965);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           n4975, QN => n966);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           n4976, QN => n967);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           n4977, QN => n968);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => 
                           n4810, QN => n737);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           n4811, QN => n738);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n4812, QN => n739);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n4813, QN => n740);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n4814, QN => n741);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n4815, QN => n742);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n4816, QN => n743);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n4817, QN => n744);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => 
                           n4778, QN => n705);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => 
                           n4779, QN => n706);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n4780, QN => n707);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n4781, QN => n708);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n4782, QN => n709);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n4783, QN => n710);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n4784, QN => n711);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n4785, QN => n712);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => 
                           n4618, QN => n481);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n4619, QN => n482);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n4620, QN => n483);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n4621, QN => n484);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n4622, QN => n485);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n4623, QN => n486);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n4624, QN => n487);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n4625, QN => n488);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => 
                           n4586, QN => n449);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           n4587, QN => n450);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n4588, QN => n451);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n4589, QN => n452);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n4590, QN => n453);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n4591, QN => n454);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n4592, QN => n455);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n4593, QN => n456);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n4426
                           , QN => n225);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n4427
                           , QN => n226);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => n4428
                           , QN => n227);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => n4429
                           , QN => n228);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => n4430
                           , QN => n229);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => n4431
                           , QN => n230);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => n4432
                           , QN => n231);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => n4433
                           , QN => n232);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n4394
                           , QN => n193);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n4395
                           , QN => n194);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => n4396
                           , QN => n195);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => n4397
                           , QN => n196);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => n4398
                           , QN => n197);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => n4399
                           , QN => n198);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => n4400
                           , QN => n199);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => n4401
                           , QN => n200);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           n4978, QN => n969);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           n4979, QN => n970);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           n4980, QN => n971);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           n4981, QN => n972);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           n4982, QN => n973);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           n4983, QN => n974);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           n4984, QN => n975);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           n4985, QN => n976);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           n4986, QN => n977);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           n4987, QN => n978);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           n4988, QN => n979);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           n4989, QN => n980);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           n4990, QN => n981);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n4991, QN => n982);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => n4992
                           , QN => n983);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => n4993
                           , QN => n984);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => n4994
                           , QN => n985);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => n4995
                           , QN => n986);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => n4996
                           , QN => n987);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => n4997
                           , QN => n988);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => n4998
                           , QN => n989);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => n4999
                           , QN => n990);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => n5000
                           , QN => n991);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => n5001
                           , QN => n992);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n4818, QN => n745);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n4819, QN => n746);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n4820, QN => n747);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n4821, QN => n748);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n4822, QN => n749);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n4823, QN => n750);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n4824, QN => n751);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n4825, QN => n752);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n4826, QN => n753);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n4827, QN => n754);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n4828, QN => n755);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n4829, QN => n756);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n4830, QN => n757);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n4831, QN => n758);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => n4832
                           , QN => n759);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => n4833
                           , QN => n760);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => n4834
                           , QN => n761);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => n4835
                           , QN => n762);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => n4836
                           , QN => n763);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => n4837
                           , QN => n764);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => n4838
                           , QN => n765);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => n4839
                           , QN => n766);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => n4840
                           , QN => n767);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => n4841
                           , QN => n768);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n4786, QN => n713);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n4787, QN => n714);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n4788, QN => n715);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n4789, QN => n716);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n4790, QN => n717);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n4791, QN => n718);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n4792, QN => n719);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n4793, QN => n720);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n4794, QN => n721);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n4795, QN => n722);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n4796, QN => n723);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n4797, QN => n724);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n4798, QN => n725);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n4799, QN => n726);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => n4800
                           , QN => n727);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => n4801
                           , QN => n728);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n4802
                           , QN => n729);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => n4803
                           , QN => n730);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => n4804
                           , QN => n731);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => n4805
                           , QN => n732);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => n4806
                           , QN => n733);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => n4807
                           , QN => n734);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => n4808
                           , QN => n735);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => n4809
                           , QN => n736);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n4626, QN => n489);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n4627, QN => n490);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n4628, QN => n491);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n4629, QN => n492);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n4630, QN => n493);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n4631, QN => n494);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n4632, QN => n495);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n4633, QN => n496);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n4634, QN => n497);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n4635, QN => n498);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n4636, QN => n499);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n4637, QN => n500);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n4638, QN => n501);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n4639, QN => n502);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => n4640
                           , QN => n503);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => n4641
                           , QN => n504);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n4642
                           , QN => n505);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => n4643
                           , QN => n506);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n4644
                           , QN => n507);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => n4645
                           , QN => n508);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n4646
                           , QN => n509);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => n4647
                           , QN => n510);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n4648
                           , QN => n511);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => n4649
                           , QN => n512);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n4594, QN => n457);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n4595, QN => n458);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n4596, QN => n459);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n4597, QN => n460);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n4598, QN => n461);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n4599, QN => n462);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n4600, QN => n463);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n4601, QN => n464);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n4602, QN => n465);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n4603, QN => n466);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n4604, QN => n467);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n4605, QN => n468);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n4606, QN => n469);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n4607, QN => n470);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => n4608
                           , QN => n471);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => n4609
                           , QN => n472);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n4610
                           , QN => n473);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => n4611
                           , QN => n474);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => n4612
                           , QN => n475);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => n4613
                           , QN => n476);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => n4614
                           , QN => n477);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => n4615
                           , QN => n478);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => n4616
                           , QN => n479);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => n4617
                           , QN => n480);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => n4434
                           , QN => n233);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => n4435
                           , QN => n234);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => n4436
                           , QN => n235);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => n4437
                           , QN => n236);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => n4438
                           , QN => n237);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => n4439
                           , QN => n238);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => n4440
                           , QN => n239);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n4441
                           , QN => n240);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n4442
                           , QN => n241);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n4443
                           , QN => n242);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n4444
                           , QN => n243);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n4445
                           , QN => n244);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n4446
                           , QN => n245);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n4447
                           , QN => n246);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n4448,
                           QN => n247);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n4449,
                           QN => n248);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n4450,
                           QN => n249);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n4451,
                           QN => n250);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n4452,
                           QN => n251);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n4453,
                           QN => n252);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n4454,
                           QN => n253);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n4455,
                           QN => n254);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n4456,
                           QN => n255);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n4457,
                           QN => n256);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => n4402
                           , QN => n201);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => n4403
                           , QN => n202);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => n4404
                           , QN => n203);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => n4405
                           , QN => n204);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => n4406
                           , QN => n205);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => n4407
                           , QN => n206);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => n4408
                           , QN => n207);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n4409
                           , QN => n208);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n4410
                           , QN => n209);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n4411
                           , QN => n210);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n4412
                           , QN => n211);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n4413
                           , QN => n212);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n4414
                           , QN => n213);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n4415
                           , QN => n214);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n4416,
                           QN => n215);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n4417,
                           QN => n216);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n4418,
                           QN => n217);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n4419,
                           QN => n218);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n4420,
                           QN => n219);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n4421,
                           QN => n220);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n4422,
                           QN => n221);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n4423,
                           QN => n222);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n4424,
                           QN => n223);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n4425,
                           QN => n224);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => 
                           n_1255, QN => n769);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => 
                           n_1256, QN => n4938);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           n_1257, QN => n4939);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n_1258, QN => n4940);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n_1259, QN => n4941);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n_1260, QN => n4942);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n_1261, QN => n4943);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n_1262, QN => n4944);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n_1263, QN => n4945);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => 
                           n_1264, QN => n4746);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => 
                           n_1265, QN => n4747);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           n_1266, QN => n4748);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => 
                           n_1267, QN => n4749);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           n_1268, QN => n4750);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           n_1269, QN => n4751);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           n_1270, QN => n4752);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           n_1271, QN => n4753);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => 
                           n_1272, QN => n4554);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => 
                           n_1273, QN => n4555);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n_1274, QN => n4556);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n_1275, QN => n4557);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n_1276, QN => n4558);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n_1277, QN => n4559);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n_1278, QN => n4560);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n_1279, QN => n4561);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => 
                           n_1280, QN => n4362);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => 
                           n_1281, QN => n4363);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           n_1282, QN => n4364);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           n_1283, QN => n4365);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           n_1284, QN => n4366);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           n_1285, QN => n4367);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           n_1286, QN => n4368);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           n_1287, QN => n4369);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => 
                           n_1288, QN => n4906);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => 
                           n_1289, QN => n4907);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n_1290, QN => n4908);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n_1291, QN => n4909);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n_1292, QN => n4910);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n_1293, QN => n4911);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n_1294, QN => n4912);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n_1295, QN => n4913);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => 
                           n_1296, QN => n4714);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => 
                           n_1297, QN => n4715);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           n_1298, QN => n4716);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           n_1299, QN => n4717);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           n_1300, QN => n4718);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           n_1301, QN => n4719);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           n_1302, QN => n4720);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           n_1303, QN => n4721);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => 
                           n_1304, QN => n4522);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => 
                           n_1305, QN => n4523);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n_1306, QN => n4524);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n_1307, QN => n4525);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n_1308, QN => n4526);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n_1309, QN => n4527);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n_1310, QN => n4528);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n_1311, QN => n4529);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => 
                           n_1312, QN => n4330);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => 
                           n_1313, QN => n4331);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           n_1314, QN => n4332);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           n_1315, QN => n4333);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           n_1316, QN => n4334);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           n_1317, QN => n4335);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           n_1318, QN => n4336);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           n_1319, QN => n4337);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n_1320, QN => n4946);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n_1321, QN => n4947);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n_1322, QN => n4948);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n_1323, QN => n4949);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n_1324, QN => n4950);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n_1325, QN => n4951);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n_1326, QN => n4952);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n_1327, QN => n4953);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n_1328, QN => n4954);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n_1329, QN => n4955);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n_1330, QN => n4956);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n_1331, QN => n4957);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n_1332, QN => n4958);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n_1333, QN => n4959);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n_1334, QN => n4960);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => 
                           n_1335, QN => n4961);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => 
                           n_1336, QN => n4962);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => 
                           n_1337, QN => n4963);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => 
                           n_1338, QN => n4964);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => 
                           n_1339, QN => n4965);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => 
                           n_1340, QN => n4966);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => 
                           n_1341, QN => n4967);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => 
                           n_1342, QN => n4968);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => 
                           n_1343, QN => n4969);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           n_1344, QN => n4754);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           n_1345, QN => n4755);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           n_1346, QN => n4756);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           n_1347, QN => n4757);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           n_1348, QN => n4758);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           n_1349, QN => n4759);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           n_1350, QN => n4760);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           n_1351, QN => n4761);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           n_1352, QN => n4762);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           n_1353, QN => n4763);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           n_1354, QN => n4764);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           n_1355, QN => n4765);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           n_1356, QN => n4766);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           n_1357, QN => n4767);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           n_1358, QN => n4768);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           n_1359, QN => n4769);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => 
                           n_1360, QN => n4770);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => 
                           n_1361, QN => n4771);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => 
                           n_1362, QN => n4772);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => 
                           n_1363, QN => n4773);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => 
                           n_1364, QN => n4774);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => 
                           n_1365, QN => n4775);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => 
                           n_1366, QN => n4776);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => 
                           n_1367, QN => n4777);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n_1368, QN => n4562);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n_1369, QN => n4563);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n_1370, QN => n4564);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n_1371, QN => n4565);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n_1372, QN => n4566);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n_1373, QN => n4567);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n_1374, QN => n4568);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           n_1375, QN => n4569);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           n_1376, QN => n4570);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           n_1377, QN => n4571);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           n_1378, QN => n4572);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           n_1379, QN => n4573);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           n_1380, QN => n4574);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           n_1381, QN => n4575);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => 
                           n_1382, QN => n4576);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           n_1383, QN => n4577);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => 
                           n_1384, QN => n4578);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => 
                           n_1385, QN => n4579);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => 
                           n_1386, QN => n4580);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => 
                           n_1387, QN => n4581);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => 
                           n_1388, QN => n4582);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => 
                           n_1389, QN => n4583);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => 
                           n_1390, QN => n4584);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => 
                           n_1391, QN => n4585);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           n_1392, QN => n4370);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           n_1393, QN => n4371);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           n_1394, QN => n4372);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           n_1395, QN => n4373);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           n_1396, QN => n4374);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           n_1397, QN => n4375);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           n_1398, QN => n4376);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => 
                           n_1399, QN => n4377);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => 
                           n_1400, QN => n4378);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => 
                           n_1401, QN => n4379);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => 
                           n_1402, QN => n4380);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => 
                           n_1403, QN => n4381);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => 
                           n_1404, QN => n4382);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => 
                           n_1405, QN => n4383);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n_1406
                           , QN => n4384);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n_1407
                           , QN => n4385);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n_1408
                           , QN => n4386);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n_1409
                           , QN => n4387);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n_1410
                           , QN => n4388);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n_1411
                           , QN => n4389);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n_1412
                           , QN => n4390);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n_1413
                           , QN => n4391);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n_1414
                           , QN => n4392);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n_1415
                           , QN => n4393);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n_1416, QN => n4914);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n_1417, QN => n4915);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n_1418, QN => n4916);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n_1419, QN => n4917);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n_1420, QN => n4918);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n_1421, QN => n4919);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n_1422, QN => n4920);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n_1423, QN => n4921);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n_1424, QN => n4922);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n_1425, QN => n4923);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n_1426, QN => n4924);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n_1427, QN => n4925);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n_1428, QN => n4926);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n_1429, QN => n4927);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n_1430, QN => n4928);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => 
                           n_1431, QN => n4929);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => 
                           n_1432, QN => n4930);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => 
                           n_1433, QN => n4931);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => 
                           n_1434, QN => n4932);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => 
                           n_1435, QN => n4933);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => 
                           n_1436, QN => n4934);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => 
                           n_1437, QN => n4935);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => 
                           n_1438, QN => n4936);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => 
                           n_1439, QN => n4937);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           n_1440, QN => n4722);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           n_1441, QN => n4723);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           n_1442, QN => n4724);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           n_1443, QN => n4725);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           n_1444, QN => n4726);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           n_1445, QN => n4727);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           n_1446, QN => n4728);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           n_1447, QN => n4729);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           n_1448, QN => n4730);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           n_1449, QN => n4731);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           n_1450, QN => n4732);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           n_1451, QN => n4733);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           n_1452, QN => n4734);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           n_1453, QN => n4735);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           n_1454, QN => n4736);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           n_1455, QN => n4737);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => 
                           n_1456, QN => n4738);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => 
                           n_1457, QN => n4739);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => 
                           n_1458, QN => n4740);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => 
                           n_1459, QN => n4741);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => 
                           n_1460, QN => n4742);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => 
                           n_1461, QN => n4743);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => 
                           n_1462, QN => n4744);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => 
                           n_1463, QN => n4745);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n_1464, QN => n4530);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n_1465, QN => n4531);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n_1466, QN => n4532);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n_1467, QN => n4533);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n_1468, QN => n4534);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n_1469, QN => n4535);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n_1470, QN => n4536);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           n_1471, QN => n4537);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           n_1472, QN => n4538);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           n_1473, QN => n4539);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           n_1474, QN => n4540);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           n_1475, QN => n4541);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           n_1476, QN => n4542);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           n_1477, QN => n4543);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           n_1478, QN => n4544);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => 
                           n_1479, QN => n4545);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => 
                           n_1480, QN => n4546);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => 
                           n_1481, QN => n4547);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => 
                           n_1482, QN => n4548);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => 
                           n_1483, QN => n4549);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => 
                           n_1484, QN => n4550);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => 
                           n_1485, QN => n4551);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => 
                           n_1486, QN => n4552);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => 
                           n_1487, QN => n4553);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           n_1488, QN => n4338);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           n_1489, QN => n4339);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           n_1490, QN => n4340);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           n_1491, QN => n4341);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           n_1492, QN => n4342);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           n_1493, QN => n4343);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           n_1494, QN => n4344);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => 
                           n_1495, QN => n4345);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => 
                           n_1496, QN => n4346);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => 
                           n_1497, QN => n4347);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => 
                           n_1498, QN => n4348);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => 
                           n_1499, QN => n4349);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => 
                           n_1500, QN => n4350);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => 
                           n_1501, QN => n4351);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n_1502
                           , QN => n4352);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n_1503
                           , QN => n4353);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n_1504
                           , QN => n4354);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n_1505
                           , QN => n4355);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n_1506
                           , QN => n4356);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n_1507
                           , QN => n4357);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n_1508
                           , QN => n4358);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n_1509
                           , QN => n4359);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n_1510
                           , QN => n4360);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n_1511
                           , QN => n4361);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => 
                           n6616, QN => n4874);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => 
                           n6615, QN => n4875);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n6614, QN => n4876);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n6613, QN => n4877);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n6612, QN => n4878);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n6611, QN => n4879);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n6610, QN => n4880);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n6609, QN => n4881);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => 
                           n6712, QN => n4682);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           n6711, QN => n4683);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n6710, QN => n4684);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n6709, QN => n4685);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n6708, QN => n4686);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n6707, QN => n4687);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n6706, QN => n4688);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n6705, QN => n4689);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => 
                           n6808, QN => n4490);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           n6807, QN => n4491);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n6806, QN => n4492);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n6805, QN => n4493);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n6804, QN => n4494);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n6803, QN => n4495);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n6802, QN => n4496);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n6801, QN => n4497);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n6904
                           , QN => n4298);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n6903
                           , QN => n4299);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n6902
                           , QN => n4300);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n6901
                           , QN => n4301);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n6900
                           , QN => n4302);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n6899
                           , QN => n4303);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n6898
                           , QN => n4304);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n6897
                           , QN => n4305);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n6608, QN => n4882);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n6607, QN => n4883);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n6606, QN => n4884);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n6605, QN => n4885);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n6604, QN => n4886);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n6603, QN => n4887);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n6602, QN => n4888);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n6601, QN => n4889);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n6600, QN => n4890);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n6599, QN => n4891);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n6598, QN => n4892);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n6597, QN => n4893);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n6596, QN => n4894);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n6595, QN => n4895);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => n6594
                           , QN => n4896);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => n6593
                           , QN => n4897);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => n6440
                           , QN => n4898);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => n6439
                           , QN => n4899);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => n6438
                           , QN => n4900);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => n6437
                           , QN => n4901);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => n6436
                           , QN => n4902);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => n6435
                           , QN => n4903);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => n6434
                           , QN => n4904);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => n6433
                           , QN => n4905);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n6704, QN => n4690);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n6703, QN => n4691);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n6702, QN => n4692);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n6701, QN => n4693);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n6700, QN => n4694);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n6699, QN => n4695);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n6698, QN => n4696);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n6697, QN => n4697);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n6696, QN => n4698);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n6695, QN => n4699);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n6694, QN => n4700);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n6693, QN => n4701);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n6692, QN => n4702);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n6691, QN => n4703);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => n6690
                           , QN => n4704);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => n6689
                           , QN => n4705);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => n6472
                           , QN => n4706);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => n6471
                           , QN => n4707);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => n6470
                           , QN => n4708);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => n6469
                           , QN => n4709);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => n6468
                           , QN => n4710);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => n6467
                           , QN => n4711);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => n6466
                           , QN => n4712);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => n6465
                           , QN => n4713);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n6800, QN => n4498);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n6799, QN => n4499);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n6798, QN => n4500);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n6797, QN => n4501);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n6796, QN => n4502);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n6795, QN => n4503);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n6794, QN => n4504);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n6793, QN => n4505);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n6792, QN => n4506);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n6791, QN => n4507);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n6790, QN => n4508);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n6789, QN => n4509);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n6788, QN => n4510);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n6787, QN => n4511);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => n6786
                           , QN => n4512);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => n6785
                           , QN => n4513);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n6504
                           , QN => n4514);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n6503
                           , QN => n4515);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n6502
                           , QN => n4516);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n6501
                           , QN => n4517);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n6500
                           , QN => n4518);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n6499
                           , QN => n4519);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n6498
                           , QN => n4520);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n6497
                           , QN => n4521);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n6896
                           , QN => n4306);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n6895
                           , QN => n4307);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n6894
                           , QN => n4308);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n6893
                           , QN => n4309);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n6892
                           , QN => n4310);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n6891
                           , QN => n4311);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n6890
                           , QN => n4312);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n6889
                           , QN => n4313);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n6888
                           , QN => n4314);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n6887
                           , QN => n4315);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n6886
                           , QN => n4316);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n6885
                           , QN => n4317);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n6884
                           , QN => n4318);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n6883
                           , QN => n4319);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n6882,
                           QN => n4320);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n6881,
                           QN => n4321);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n6536,
                           QN => n4322);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n6535,
                           QN => n4323);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n6534,
                           QN => n4324);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n6533,
                           QN => n4325);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n6532,
                           QN => n4326);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n6531,
                           QN => n4327);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n6530,
                           QN => n4328);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n6529,
                           QN => n4329);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => 
                           n6640, QN => n4842);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => 
                           n6639, QN => n4843);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           n6638, QN => n4844);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           n6637, QN => n4845);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           n6636, QN => n4846);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           n6635, QN => n4847);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           n6634, QN => n4848);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           n6633, QN => n4849);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => 
                           n6736, QN => n4650);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => 
                           n6735, QN => n4651);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n6734, QN => n4652);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n6733, QN => n4653);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n6732, QN => n4654);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n6731, QN => n4655);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n6730, QN => n4656);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n6729, QN => n4657);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => 
                           n6832, QN => n4458);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => 
                           n6831, QN => n4459);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n6830, QN => n4460);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n6829, QN => n4461);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n6828, QN => n4462);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n6827, QN => n4463);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n6826, QN => n4464);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n6825, QN => n4465);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n6928
                           , QN => n4266);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n6927
                           , QN => n4267);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n6926
                           , QN => n4268);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n6925
                           , QN => n4269);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n6924
                           , QN => n4270);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n6923
                           , QN => n4271);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n6922
                           , QN => n4272);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n6921
                           , QN => n4273);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           n6632, QN => n4850);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           n6631, QN => n4851);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           n6630, QN => n4852);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           n6629, QN => n4853);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           n6628, QN => n4854);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           n6627, QN => n4855);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           n6626, QN => n4856);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => 
                           n6625, QN => n4857);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n6624, QN => n4858);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n6623, QN => n4859);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n6622, QN => n4860);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n6621, QN => n4861);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n6620, QN => n4862);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n6619, QN => n4863);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => n6618
                           , QN => n4864);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => n6617
                           , QN => n4865);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => n6448
                           , QN => n4866);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => n6447
                           , QN => n4867);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => n6446
                           , QN => n4868);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => n6445
                           , QN => n4869);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => n6444
                           , QN => n4870);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => n6443
                           , QN => n4871);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => n6442
                           , QN => n4872);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => n6441
                           , QN => n4873);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n6728, QN => n4658);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n6727, QN => n4659);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n6726, QN => n4660);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n6725, QN => n4661);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n6724, QN => n4662);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n6723, QN => n4663);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n6722, QN => n4664);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n6721, QN => n4665);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n6720, QN => n4666);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n6719, QN => n4667);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n6718, QN => n4668);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n6717, QN => n4669);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n6716, QN => n4670);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n6715, QN => n4671);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => n6714
                           , QN => n4672);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => n6713
                           , QN => n4673);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => n6480
                           , QN => n4674);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n6479
                           , QN => n4675);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => n6478
                           , QN => n4676);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n6477
                           , QN => n4677);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => n6476
                           , QN => n4678);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n6475
                           , QN => n4679);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => n6474
                           , QN => n4680);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n6473
                           , QN => n4681);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n6824, QN => n4466);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n6823, QN => n4467);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n6822, QN => n4468);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n6821, QN => n4469);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n6820, QN => n4470);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n6819, QN => n4471);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n6818, QN => n4472);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n6817, QN => n4473);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n6816, QN => n4474);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n6815, QN => n4475);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n6814, QN => n4476);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n6813, QN => n4477);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n6812, QN => n4478);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n6811, QN => n4479);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => n6810
                           , QN => n4480);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => n6809
                           , QN => n4481);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n6512
                           , QN => n4482);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n6511
                           , QN => n4483);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n6510
                           , QN => n4484);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n6509
                           , QN => n4485);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n6508
                           , QN => n4486);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n6507
                           , QN => n4487);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n6506
                           , QN => n4488);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n6505
                           , QN => n4489);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n6920
                           , QN => n4274);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n6919
                           , QN => n4275);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n6918
                           , QN => n4276);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n6917
                           , QN => n4277);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n6916
                           , QN => n4278);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n6915
                           , QN => n4279);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n6914
                           , QN => n4280);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n6913
                           , QN => n4281);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n6912
                           , QN => n4282);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n6911
                           , QN => n4283);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n6910
                           , QN => n4284);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n6909
                           , QN => n4285);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n6908
                           , QN => n4286);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n6907
                           , QN => n4287);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n6906,
                           QN => n4288);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n6905,
                           QN => n4289);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n6544,
                           QN => n4290);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n6543,
                           QN => n4291);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n6542,
                           QN => n4292);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n6541,
                           QN => n4293);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n6540,
                           QN => n4294);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n6539,
                           QN => n4295);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n6538,
                           QN => n4296);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n6537,
                           QN => n4297);
   U5877 : INV_X1 port map( A => n7577, ZN => n7570);
   U5878 : INV_X1 port map( A => n7214, ZN => n7207);
   U5879 : INV_X1 port map( A => n7259, ZN => n7252);
   U5880 : INV_X1 port map( A => n7268, ZN => n7261);
   U5881 : INV_X1 port map( A => n7277, ZN => n7270);
   U5882 : INV_X1 port map( A => n7286, ZN => n7279);
   U5883 : INV_X1 port map( A => n7331, ZN => n7324);
   U5884 : INV_X1 port map( A => n7340, ZN => n7333);
   U5885 : INV_X1 port map( A => n7349, ZN => n7342);
   U5886 : INV_X1 port map( A => n7358, ZN => n7351);
   U5887 : INV_X1 port map( A => n7403, ZN => n7396);
   U5888 : INV_X1 port map( A => n7412, ZN => n7405);
   U5889 : INV_X1 port map( A => n7421, ZN => n7414);
   U5890 : INV_X1 port map( A => n7430, ZN => n7423);
   U5891 : INV_X1 port map( A => n7475, ZN => n7468);
   U5892 : INV_X1 port map( A => n7223, ZN => n7216);
   U5893 : INV_X1 port map( A => n7232, ZN => n7225);
   U5894 : INV_X1 port map( A => n7241, ZN => n7234);
   U5895 : INV_X1 port map( A => n7250, ZN => n7243);
   U5896 : INV_X1 port map( A => n7295, ZN => n7288);
   U5897 : INV_X1 port map( A => n7304, ZN => n7297);
   U5898 : INV_X1 port map( A => n7313, ZN => n7306);
   U5899 : INV_X1 port map( A => n7322, ZN => n7315);
   U5900 : INV_X1 port map( A => n7367, ZN => n7360);
   U5901 : INV_X1 port map( A => n7376, ZN => n7369);
   U5902 : INV_X1 port map( A => n7385, ZN => n7378);
   U5903 : INV_X1 port map( A => n7394, ZN => n7387);
   U5904 : INV_X1 port map( A => n7439, ZN => n7432);
   U5905 : INV_X1 port map( A => n7448, ZN => n7441);
   U5906 : INV_X1 port map( A => n7457, ZN => n7450);
   U5907 : INV_X1 port map( A => n7466, ZN => n7459);
   U5908 : BUF_X1 port map( A => n7578, Z => n7571);
   U5909 : BUF_X1 port map( A => n7578, Z => n7572);
   U5910 : BUF_X1 port map( A => n7578, Z => n7573);
   U5911 : BUF_X1 port map( A => n7578, Z => n7574);
   U5912 : BUF_X1 port map( A => n7578, Z => n7575);
   U5913 : BUF_X1 port map( A => n7578, Z => n7576);
   U5914 : BUF_X1 port map( A => n7578, Z => n7577);
   U5915 : BUF_X1 port map( A => n7206, Z => n7198);
   U5916 : BUF_X1 port map( A => n7206, Z => n7199);
   U5917 : BUF_X1 port map( A => n7206, Z => n7200);
   U5918 : BUF_X1 port map( A => n7206, Z => n7201);
   U5919 : BUF_X1 port map( A => n7206, Z => n7202);
   U5920 : BUF_X1 port map( A => n7206, Z => n7203);
   U5921 : BUF_X1 port map( A => n7203, Z => n7204);
   U5922 : BUF_X1 port map( A => n7198, Z => n7205);
   U5923 : BUF_X1 port map( A => n5775, Z => n7080);
   U5924 : BUF_X1 port map( A => n5785, Z => n7056);
   U5925 : BUF_X1 port map( A => n5780, Z => n7068);
   U5926 : BUF_X1 port map( A => n5790, Z => n7044);
   U5927 : BUF_X1 port map( A => n5799, Z => n7032);
   U5928 : BUF_X1 port map( A => n5809, Z => n7008);
   U5929 : BUF_X1 port map( A => n5804, Z => n7020);
   U5930 : BUF_X1 port map( A => n5814, Z => n6996);
   U5931 : BUF_X1 port map( A => n5775, Z => n7081);
   U5932 : BUF_X1 port map( A => n5785, Z => n7057);
   U5933 : BUF_X1 port map( A => n5780, Z => n7069);
   U5934 : BUF_X1 port map( A => n5790, Z => n7045);
   U5935 : BUF_X1 port map( A => n5799, Z => n7033);
   U5936 : BUF_X1 port map( A => n5809, Z => n7009);
   U5937 : BUF_X1 port map( A => n5804, Z => n7021);
   U5938 : BUF_X1 port map( A => n5814, Z => n6997);
   U5939 : BUF_X1 port map( A => n5122, Z => n7182);
   U5940 : BUF_X1 port map( A => n5132, Z => n7158);
   U5941 : BUF_X1 port map( A => n5127, Z => n7170);
   U5942 : BUF_X1 port map( A => n5137, Z => n7146);
   U5943 : BUF_X1 port map( A => n5146, Z => n7134);
   U5944 : BUF_X1 port map( A => n5156, Z => n7110);
   U5945 : BUF_X1 port map( A => n5151, Z => n7122);
   U5946 : BUF_X1 port map( A => n5161, Z => n7098);
   U5947 : BUF_X1 port map( A => n5122, Z => n7183);
   U5948 : BUF_X1 port map( A => n5132, Z => n7159);
   U5949 : BUF_X1 port map( A => n5127, Z => n7171);
   U5950 : BUF_X1 port map( A => n5137, Z => n7147);
   U5951 : BUF_X1 port map( A => n5146, Z => n7135);
   U5952 : BUF_X1 port map( A => n5156, Z => n7111);
   U5953 : BUF_X1 port map( A => n5151, Z => n7123);
   U5954 : BUF_X1 port map( A => n5161, Z => n7099);
   U5955 : BUF_X1 port map( A => n5776, Z => n7077);
   U5956 : BUF_X1 port map( A => n5786, Z => n7053);
   U5957 : BUF_X1 port map( A => n5781, Z => n7065);
   U5958 : BUF_X1 port map( A => n5791, Z => n7041);
   U5959 : BUF_X1 port map( A => n5800, Z => n7029);
   U5960 : BUF_X1 port map( A => n5810, Z => n7005);
   U5961 : BUF_X1 port map( A => n5805, Z => n7017);
   U5962 : BUF_X1 port map( A => n5815, Z => n6993);
   U5963 : BUF_X1 port map( A => n5776, Z => n7078);
   U5964 : BUF_X1 port map( A => n5786, Z => n7054);
   U5965 : BUF_X1 port map( A => n5781, Z => n7066);
   U5966 : BUF_X1 port map( A => n5791, Z => n7042);
   U5967 : BUF_X1 port map( A => n5800, Z => n7030);
   U5968 : BUF_X1 port map( A => n5810, Z => n7006);
   U5969 : BUF_X1 port map( A => n5805, Z => n7018);
   U5970 : BUF_X1 port map( A => n5815, Z => n6994);
   U5971 : BUF_X1 port map( A => n5123, Z => n7179);
   U5972 : BUF_X1 port map( A => n5133, Z => n7155);
   U5973 : BUF_X1 port map( A => n5128, Z => n7167);
   U5974 : BUF_X1 port map( A => n5138, Z => n7143);
   U5975 : BUF_X1 port map( A => n5147, Z => n7131);
   U5976 : BUF_X1 port map( A => n5157, Z => n7107);
   U5977 : BUF_X1 port map( A => n5152, Z => n7119);
   U5978 : BUF_X1 port map( A => n5162, Z => n7095);
   U5979 : BUF_X1 port map( A => n5123, Z => n7180);
   U5980 : BUF_X1 port map( A => n5133, Z => n7156);
   U5981 : BUF_X1 port map( A => n5128, Z => n7168);
   U5982 : BUF_X1 port map( A => n5138, Z => n7144);
   U5983 : BUF_X1 port map( A => n5147, Z => n7132);
   U5984 : BUF_X1 port map( A => n5157, Z => n7108);
   U5985 : BUF_X1 port map( A => n5152, Z => n7120);
   U5986 : BUF_X1 port map( A => n5162, Z => n7096);
   U5987 : BUF_X1 port map( A => n5772, Z => n7086);
   U5988 : BUF_X1 port map( A => n5782, Z => n7062);
   U5989 : BUF_X1 port map( A => n5777, Z => n7074);
   U5990 : BUF_X1 port map( A => n5787, Z => n7050);
   U5991 : BUF_X1 port map( A => n5796, Z => n7038);
   U5992 : BUF_X1 port map( A => n5806, Z => n7014);
   U5993 : BUF_X1 port map( A => n5801, Z => n7026);
   U5994 : BUF_X1 port map( A => n5811, Z => n7002);
   U5995 : BUF_X1 port map( A => n5772, Z => n7087);
   U5996 : BUF_X1 port map( A => n5782, Z => n7063);
   U5997 : BUF_X1 port map( A => n5777, Z => n7075);
   U5998 : BUF_X1 port map( A => n5787, Z => n7051);
   U5999 : BUF_X1 port map( A => n5796, Z => n7039);
   U6000 : BUF_X1 port map( A => n5806, Z => n7015);
   U6001 : BUF_X1 port map( A => n5801, Z => n7027);
   U6002 : BUF_X1 port map( A => n5811, Z => n7003);
   U6003 : BUF_X1 port map( A => n5119, Z => n7188);
   U6004 : BUF_X1 port map( A => n5129, Z => n7164);
   U6005 : BUF_X1 port map( A => n5124, Z => n7176);
   U6006 : BUF_X1 port map( A => n5134, Z => n7152);
   U6007 : BUF_X1 port map( A => n5143, Z => n7140);
   U6008 : BUF_X1 port map( A => n5153, Z => n7116);
   U6009 : BUF_X1 port map( A => n5148, Z => n7128);
   U6010 : BUF_X1 port map( A => n5158, Z => n7104);
   U6011 : BUF_X1 port map( A => n5119, Z => n7189);
   U6012 : BUF_X1 port map( A => n5129, Z => n7165);
   U6013 : BUF_X1 port map( A => n5124, Z => n7177);
   U6014 : BUF_X1 port map( A => n5134, Z => n7153);
   U6015 : BUF_X1 port map( A => n5143, Z => n7141);
   U6016 : BUF_X1 port map( A => n5153, Z => n7117);
   U6017 : BUF_X1 port map( A => n5148, Z => n7129);
   U6018 : BUF_X1 port map( A => n5158, Z => n7105);
   U6019 : BUF_X1 port map( A => n5773, Z => n7083);
   U6020 : BUF_X1 port map( A => n5783, Z => n7059);
   U6021 : BUF_X1 port map( A => n5778, Z => n7071);
   U6022 : BUF_X1 port map( A => n5788, Z => n7047);
   U6023 : BUF_X1 port map( A => n5797, Z => n7035);
   U6024 : BUF_X1 port map( A => n5807, Z => n7011);
   U6025 : BUF_X1 port map( A => n5802, Z => n7023);
   U6026 : BUF_X1 port map( A => n5812, Z => n6999);
   U6027 : BUF_X1 port map( A => n5773, Z => n7084);
   U6028 : BUF_X1 port map( A => n5783, Z => n7060);
   U6029 : BUF_X1 port map( A => n5778, Z => n7072);
   U6030 : BUF_X1 port map( A => n5788, Z => n7048);
   U6031 : BUF_X1 port map( A => n5797, Z => n7036);
   U6032 : BUF_X1 port map( A => n5807, Z => n7012);
   U6033 : BUF_X1 port map( A => n5802, Z => n7024);
   U6034 : BUF_X1 port map( A => n5812, Z => n7000);
   U6035 : BUF_X1 port map( A => n5120, Z => n7185);
   U6036 : BUF_X1 port map( A => n5130, Z => n7161);
   U6037 : BUF_X1 port map( A => n5125, Z => n7173);
   U6038 : BUF_X1 port map( A => n5135, Z => n7149);
   U6039 : BUF_X1 port map( A => n5144, Z => n7137);
   U6040 : BUF_X1 port map( A => n5154, Z => n7113);
   U6041 : BUF_X1 port map( A => n5149, Z => n7125);
   U6042 : BUF_X1 port map( A => n5159, Z => n7101);
   U6043 : BUF_X1 port map( A => n5120, Z => n7186);
   U6044 : BUF_X1 port map( A => n5130, Z => n7162);
   U6045 : BUF_X1 port map( A => n5125, Z => n7174);
   U6046 : BUF_X1 port map( A => n5135, Z => n7150);
   U6047 : BUF_X1 port map( A => n5144, Z => n7138);
   U6048 : BUF_X1 port map( A => n5154, Z => n7114);
   U6049 : BUF_X1 port map( A => n5149, Z => n7126);
   U6050 : BUF_X1 port map( A => n5159, Z => n7102);
   U6051 : BUF_X1 port map( A => n5775, Z => n7082);
   U6052 : BUF_X1 port map( A => n5785, Z => n7058);
   U6053 : BUF_X1 port map( A => n5780, Z => n7070);
   U6054 : BUF_X1 port map( A => n5790, Z => n7046);
   U6055 : BUF_X1 port map( A => n5799, Z => n7034);
   U6056 : BUF_X1 port map( A => n5809, Z => n7010);
   U6057 : BUF_X1 port map( A => n5804, Z => n7022);
   U6058 : BUF_X1 port map( A => n5814, Z => n6998);
   U6059 : BUF_X1 port map( A => n5122, Z => n7184);
   U6060 : BUF_X1 port map( A => n5132, Z => n7160);
   U6061 : BUF_X1 port map( A => n5127, Z => n7172);
   U6062 : BUF_X1 port map( A => n5137, Z => n7148);
   U6063 : BUF_X1 port map( A => n5146, Z => n7136);
   U6064 : BUF_X1 port map( A => n5156, Z => n7112);
   U6065 : BUF_X1 port map( A => n5151, Z => n7124);
   U6066 : BUF_X1 port map( A => n5161, Z => n7100);
   U6067 : BUF_X1 port map( A => n5776, Z => n7079);
   U6068 : BUF_X1 port map( A => n5786, Z => n7055);
   U6069 : BUF_X1 port map( A => n5781, Z => n7067);
   U6070 : BUF_X1 port map( A => n5791, Z => n7043);
   U6071 : BUF_X1 port map( A => n5800, Z => n7031);
   U6072 : BUF_X1 port map( A => n5810, Z => n7007);
   U6073 : BUF_X1 port map( A => n5805, Z => n7019);
   U6074 : BUF_X1 port map( A => n5815, Z => n6995);
   U6075 : BUF_X1 port map( A => n5123, Z => n7181);
   U6076 : BUF_X1 port map( A => n5133, Z => n7157);
   U6077 : BUF_X1 port map( A => n5128, Z => n7169);
   U6078 : BUF_X1 port map( A => n5138, Z => n7145);
   U6079 : BUF_X1 port map( A => n5147, Z => n7133);
   U6080 : BUF_X1 port map( A => n5157, Z => n7109);
   U6081 : BUF_X1 port map( A => n5152, Z => n7121);
   U6082 : BUF_X1 port map( A => n5162, Z => n7097);
   U6083 : BUF_X1 port map( A => n5772, Z => n7088);
   U6084 : BUF_X1 port map( A => n5782, Z => n7064);
   U6085 : BUF_X1 port map( A => n5777, Z => n7076);
   U6086 : BUF_X1 port map( A => n5787, Z => n7052);
   U6087 : BUF_X1 port map( A => n5796, Z => n7040);
   U6088 : BUF_X1 port map( A => n5806, Z => n7016);
   U6089 : BUF_X1 port map( A => n5801, Z => n7028);
   U6090 : BUF_X1 port map( A => n5811, Z => n7004);
   U6091 : BUF_X1 port map( A => n5119, Z => n7190);
   U6092 : BUF_X1 port map( A => n5129, Z => n7166);
   U6093 : BUF_X1 port map( A => n5124, Z => n7178);
   U6094 : BUF_X1 port map( A => n5134, Z => n7154);
   U6095 : BUF_X1 port map( A => n5143, Z => n7142);
   U6096 : BUF_X1 port map( A => n5153, Z => n7118);
   U6097 : BUF_X1 port map( A => n5148, Z => n7130);
   U6098 : BUF_X1 port map( A => n5158, Z => n7106);
   U6099 : BUF_X1 port map( A => n5773, Z => n7085);
   U6100 : BUF_X1 port map( A => n5783, Z => n7061);
   U6101 : BUF_X1 port map( A => n5778, Z => n7073);
   U6102 : BUF_X1 port map( A => n5788, Z => n7049);
   U6103 : BUF_X1 port map( A => n5797, Z => n7037);
   U6104 : BUF_X1 port map( A => n5807, Z => n7013);
   U6105 : BUF_X1 port map( A => n5802, Z => n7025);
   U6106 : BUF_X1 port map( A => n5812, Z => n7001);
   U6107 : BUF_X1 port map( A => n5120, Z => n7187);
   U6108 : BUF_X1 port map( A => n5130, Z => n7163);
   U6109 : BUF_X1 port map( A => n5125, Z => n7175);
   U6110 : BUF_X1 port map( A => n5135, Z => n7151);
   U6111 : BUF_X1 port map( A => n5144, Z => n7139);
   U6112 : BUF_X1 port map( A => n5154, Z => n7115);
   U6113 : BUF_X1 port map( A => n5149, Z => n7127);
   U6114 : BUF_X1 port map( A => n5159, Z => n7103);
   U6115 : BUF_X1 port map( A => n7215, Z => n7208);
   U6116 : BUF_X1 port map( A => n7215, Z => n7209);
   U6117 : BUF_X1 port map( A => n7215, Z => n7210);
   U6118 : BUF_X1 port map( A => n7215, Z => n7211);
   U6119 : BUF_X1 port map( A => n7215, Z => n7212);
   U6120 : BUF_X1 port map( A => n7215, Z => n7213);
   U6121 : BUF_X1 port map( A => n7224, Z => n7217);
   U6122 : BUF_X1 port map( A => n7224, Z => n7218);
   U6123 : BUF_X1 port map( A => n7224, Z => n7219);
   U6124 : BUF_X1 port map( A => n7224, Z => n7220);
   U6125 : BUF_X1 port map( A => n7224, Z => n7221);
   U6126 : BUF_X1 port map( A => n7224, Z => n7222);
   U6127 : BUF_X1 port map( A => n7233, Z => n7226);
   U6128 : BUF_X1 port map( A => n7233, Z => n7227);
   U6129 : BUF_X1 port map( A => n7233, Z => n7228);
   U6130 : BUF_X1 port map( A => n7233, Z => n7229);
   U6131 : BUF_X1 port map( A => n7233, Z => n7230);
   U6132 : BUF_X1 port map( A => n7233, Z => n7231);
   U6133 : BUF_X1 port map( A => n7242, Z => n7235);
   U6134 : BUF_X1 port map( A => n7242, Z => n7236);
   U6135 : BUF_X1 port map( A => n7242, Z => n7237);
   U6136 : BUF_X1 port map( A => n7242, Z => n7238);
   U6137 : BUF_X1 port map( A => n7242, Z => n7239);
   U6138 : BUF_X1 port map( A => n7242, Z => n7240);
   U6139 : BUF_X1 port map( A => n7251, Z => n7244);
   U6140 : BUF_X1 port map( A => n7251, Z => n7245);
   U6141 : BUF_X1 port map( A => n7251, Z => n7246);
   U6142 : BUF_X1 port map( A => n7251, Z => n7247);
   U6143 : BUF_X1 port map( A => n7251, Z => n7248);
   U6144 : BUF_X1 port map( A => n7251, Z => n7249);
   U6145 : BUF_X1 port map( A => n7260, Z => n7253);
   U6146 : BUF_X1 port map( A => n7260, Z => n7254);
   U6147 : BUF_X1 port map( A => n7260, Z => n7255);
   U6148 : BUF_X1 port map( A => n7260, Z => n7256);
   U6149 : BUF_X1 port map( A => n7260, Z => n7257);
   U6150 : BUF_X1 port map( A => n7260, Z => n7258);
   U6151 : BUF_X1 port map( A => n7269, Z => n7262);
   U6152 : BUF_X1 port map( A => n7269, Z => n7263);
   U6153 : BUF_X1 port map( A => n7269, Z => n7264);
   U6154 : BUF_X1 port map( A => n7269, Z => n7265);
   U6155 : BUF_X1 port map( A => n7269, Z => n7266);
   U6156 : BUF_X1 port map( A => n7269, Z => n7267);
   U6157 : BUF_X1 port map( A => n7278, Z => n7271);
   U6158 : BUF_X1 port map( A => n7278, Z => n7272);
   U6159 : BUF_X1 port map( A => n7278, Z => n7273);
   U6160 : BUF_X1 port map( A => n7278, Z => n7274);
   U6161 : BUF_X1 port map( A => n7278, Z => n7275);
   U6162 : BUF_X1 port map( A => n7278, Z => n7276);
   U6163 : BUF_X1 port map( A => n7287, Z => n7280);
   U6164 : BUF_X1 port map( A => n7287, Z => n7281);
   U6165 : BUF_X1 port map( A => n7287, Z => n7282);
   U6166 : BUF_X1 port map( A => n7287, Z => n7283);
   U6167 : BUF_X1 port map( A => n7287, Z => n7284);
   U6168 : BUF_X1 port map( A => n7287, Z => n7285);
   U6169 : BUF_X1 port map( A => n7296, Z => n7289);
   U6170 : BUF_X1 port map( A => n7296, Z => n7290);
   U6171 : BUF_X1 port map( A => n7296, Z => n7291);
   U6172 : BUF_X1 port map( A => n7296, Z => n7292);
   U6173 : BUF_X1 port map( A => n7296, Z => n7293);
   U6174 : BUF_X1 port map( A => n7296, Z => n7294);
   U6175 : BUF_X1 port map( A => n7305, Z => n7298);
   U6176 : BUF_X1 port map( A => n7305, Z => n7299);
   U6177 : BUF_X1 port map( A => n7305, Z => n7300);
   U6178 : BUF_X1 port map( A => n7305, Z => n7301);
   U6179 : BUF_X1 port map( A => n7305, Z => n7302);
   U6180 : BUF_X1 port map( A => n7305, Z => n7303);
   U6181 : BUF_X1 port map( A => n7314, Z => n7307);
   U6182 : BUF_X1 port map( A => n7314, Z => n7308);
   U6183 : BUF_X1 port map( A => n7314, Z => n7309);
   U6184 : BUF_X1 port map( A => n7314, Z => n7310);
   U6185 : BUF_X1 port map( A => n7314, Z => n7311);
   U6186 : BUF_X1 port map( A => n7314, Z => n7312);
   U6187 : BUF_X1 port map( A => n7323, Z => n7316);
   U6188 : BUF_X1 port map( A => n7323, Z => n7317);
   U6189 : BUF_X1 port map( A => n7323, Z => n7318);
   U6190 : BUF_X1 port map( A => n7323, Z => n7319);
   U6191 : BUF_X1 port map( A => n7323, Z => n7320);
   U6192 : BUF_X1 port map( A => n7323, Z => n7321);
   U6193 : BUF_X1 port map( A => n7332, Z => n7325);
   U6194 : BUF_X1 port map( A => n7332, Z => n7326);
   U6195 : BUF_X1 port map( A => n7332, Z => n7327);
   U6196 : BUF_X1 port map( A => n7332, Z => n7328);
   U6197 : BUF_X1 port map( A => n7332, Z => n7329);
   U6198 : BUF_X1 port map( A => n7332, Z => n7330);
   U6199 : BUF_X1 port map( A => n7341, Z => n7334);
   U6200 : BUF_X1 port map( A => n7341, Z => n7335);
   U6201 : BUF_X1 port map( A => n7341, Z => n7336);
   U6202 : BUF_X1 port map( A => n7341, Z => n7337);
   U6203 : BUF_X1 port map( A => n7341, Z => n7338);
   U6204 : BUF_X1 port map( A => n7341, Z => n7339);
   U6205 : BUF_X1 port map( A => n7350, Z => n7343);
   U6206 : BUF_X1 port map( A => n7350, Z => n7344);
   U6207 : BUF_X1 port map( A => n7350, Z => n7345);
   U6208 : BUF_X1 port map( A => n7350, Z => n7346);
   U6209 : BUF_X1 port map( A => n7350, Z => n7347);
   U6210 : BUF_X1 port map( A => n7350, Z => n7348);
   U6211 : BUF_X1 port map( A => n7359, Z => n7352);
   U6212 : BUF_X1 port map( A => n7359, Z => n7353);
   U6213 : BUF_X1 port map( A => n7359, Z => n7354);
   U6214 : BUF_X1 port map( A => n7359, Z => n7355);
   U6215 : BUF_X1 port map( A => n7359, Z => n7356);
   U6216 : BUF_X1 port map( A => n7359, Z => n7357);
   U6217 : BUF_X1 port map( A => n7368, Z => n7361);
   U6218 : BUF_X1 port map( A => n7368, Z => n7362);
   U6219 : BUF_X1 port map( A => n7368, Z => n7363);
   U6220 : BUF_X1 port map( A => n7368, Z => n7364);
   U6221 : BUF_X1 port map( A => n7368, Z => n7365);
   U6222 : BUF_X1 port map( A => n7368, Z => n7366);
   U6223 : BUF_X1 port map( A => n7377, Z => n7370);
   U6224 : BUF_X1 port map( A => n7377, Z => n7371);
   U6225 : BUF_X1 port map( A => n7377, Z => n7372);
   U6226 : BUF_X1 port map( A => n7377, Z => n7373);
   U6227 : BUF_X1 port map( A => n7377, Z => n7374);
   U6228 : BUF_X1 port map( A => n7377, Z => n7375);
   U6229 : BUF_X1 port map( A => n7386, Z => n7379);
   U6230 : BUF_X1 port map( A => n7386, Z => n7380);
   U6231 : BUF_X1 port map( A => n7386, Z => n7381);
   U6232 : BUF_X1 port map( A => n7386, Z => n7382);
   U6233 : BUF_X1 port map( A => n7386, Z => n7383);
   U6234 : BUF_X1 port map( A => n7386, Z => n7384);
   U6235 : BUF_X1 port map( A => n7395, Z => n7388);
   U6236 : BUF_X1 port map( A => n7395, Z => n7389);
   U6237 : BUF_X1 port map( A => n7395, Z => n7390);
   U6238 : BUF_X1 port map( A => n7395, Z => n7391);
   U6239 : BUF_X1 port map( A => n7395, Z => n7392);
   U6240 : BUF_X1 port map( A => n7395, Z => n7393);
   U6241 : BUF_X1 port map( A => n7404, Z => n7397);
   U6242 : BUF_X1 port map( A => n7404, Z => n7398);
   U6243 : BUF_X1 port map( A => n7404, Z => n7399);
   U6244 : BUF_X1 port map( A => n7404, Z => n7400);
   U6245 : BUF_X1 port map( A => n7404, Z => n7401);
   U6246 : BUF_X1 port map( A => n7404, Z => n7402);
   U6247 : BUF_X1 port map( A => n7413, Z => n7406);
   U6248 : BUF_X1 port map( A => n7413, Z => n7407);
   U6249 : BUF_X1 port map( A => n7413, Z => n7408);
   U6250 : BUF_X1 port map( A => n7413, Z => n7409);
   U6251 : BUF_X1 port map( A => n7413, Z => n7410);
   U6252 : BUF_X1 port map( A => n7413, Z => n7411);
   U6253 : BUF_X1 port map( A => n7422, Z => n7415);
   U6254 : BUF_X1 port map( A => n7422, Z => n7416);
   U6255 : BUF_X1 port map( A => n7422, Z => n7417);
   U6256 : BUF_X1 port map( A => n7422, Z => n7418);
   U6257 : BUF_X1 port map( A => n7422, Z => n7419);
   U6258 : BUF_X1 port map( A => n7422, Z => n7420);
   U6259 : BUF_X1 port map( A => n7431, Z => n7424);
   U6260 : BUF_X1 port map( A => n7431, Z => n7425);
   U6261 : BUF_X1 port map( A => n7431, Z => n7426);
   U6262 : BUF_X1 port map( A => n7431, Z => n7427);
   U6263 : BUF_X1 port map( A => n7431, Z => n7428);
   U6264 : BUF_X1 port map( A => n7431, Z => n7429);
   U6265 : BUF_X1 port map( A => n7440, Z => n7433);
   U6266 : BUF_X1 port map( A => n7440, Z => n7434);
   U6267 : BUF_X1 port map( A => n7440, Z => n7435);
   U6268 : BUF_X1 port map( A => n7440, Z => n7436);
   U6269 : BUF_X1 port map( A => n7440, Z => n7437);
   U6270 : BUF_X1 port map( A => n7440, Z => n7438);
   U6271 : BUF_X1 port map( A => n7449, Z => n7442);
   U6272 : BUF_X1 port map( A => n7449, Z => n7443);
   U6273 : BUF_X1 port map( A => n7449, Z => n7444);
   U6274 : BUF_X1 port map( A => n7449, Z => n7445);
   U6275 : BUF_X1 port map( A => n7449, Z => n7446);
   U6276 : BUF_X1 port map( A => n7449, Z => n7447);
   U6277 : BUF_X1 port map( A => n7458, Z => n7451);
   U6278 : BUF_X1 port map( A => n7458, Z => n7452);
   U6279 : BUF_X1 port map( A => n7458, Z => n7453);
   U6280 : BUF_X1 port map( A => n7458, Z => n7454);
   U6281 : BUF_X1 port map( A => n7458, Z => n7455);
   U6282 : BUF_X1 port map( A => n7458, Z => n7456);
   U6283 : BUF_X1 port map( A => n7467, Z => n7460);
   U6284 : BUF_X1 port map( A => n7467, Z => n7461);
   U6285 : BUF_X1 port map( A => n7467, Z => n7462);
   U6286 : BUF_X1 port map( A => n7467, Z => n7463);
   U6287 : BUF_X1 port map( A => n7467, Z => n7464);
   U6288 : BUF_X1 port map( A => n7467, Z => n7465);
   U6289 : BUF_X1 port map( A => n7476, Z => n7469);
   U6290 : BUF_X1 port map( A => n7476, Z => n7470);
   U6291 : BUF_X1 port map( A => n7476, Z => n7471);
   U6292 : BUF_X1 port map( A => n7476, Z => n7472);
   U6293 : BUF_X1 port map( A => n7476, Z => n7473);
   U6294 : BUF_X1 port map( A => n7476, Z => n7474);
   U6295 : BUF_X1 port map( A => n7215, Z => n7214);
   U6296 : BUF_X1 port map( A => n7224, Z => n7223);
   U6297 : BUF_X1 port map( A => n7233, Z => n7232);
   U6298 : BUF_X1 port map( A => n7242, Z => n7241);
   U6299 : BUF_X1 port map( A => n7251, Z => n7250);
   U6300 : BUF_X1 port map( A => n7260, Z => n7259);
   U6301 : BUF_X1 port map( A => n7269, Z => n7268);
   U6302 : BUF_X1 port map( A => n7278, Z => n7277);
   U6303 : BUF_X1 port map( A => n7287, Z => n7286);
   U6304 : BUF_X1 port map( A => n7296, Z => n7295);
   U6305 : BUF_X1 port map( A => n7305, Z => n7304);
   U6306 : BUF_X1 port map( A => n7314, Z => n7313);
   U6307 : BUF_X1 port map( A => n7323, Z => n7322);
   U6308 : BUF_X1 port map( A => n7332, Z => n7331);
   U6309 : BUF_X1 port map( A => n7341, Z => n7340);
   U6310 : BUF_X1 port map( A => n7350, Z => n7349);
   U6311 : BUF_X1 port map( A => n7359, Z => n7358);
   U6312 : BUF_X1 port map( A => n7368, Z => n7367);
   U6313 : BUF_X1 port map( A => n7377, Z => n7376);
   U6314 : BUF_X1 port map( A => n7386, Z => n7385);
   U6315 : BUF_X1 port map( A => n7395, Z => n7394);
   U6316 : BUF_X1 port map( A => n7404, Z => n7403);
   U6317 : BUF_X1 port map( A => n7413, Z => n7412);
   U6318 : BUF_X1 port map( A => n7422, Z => n7421);
   U6319 : BUF_X1 port map( A => n7431, Z => n7430);
   U6320 : BUF_X1 port map( A => n7440, Z => n7439);
   U6321 : BUF_X1 port map( A => n7449, Z => n7448);
   U6322 : BUF_X1 port map( A => n7458, Z => n7457);
   U6323 : BUF_X1 port map( A => n7467, Z => n7466);
   U6324 : BUF_X1 port map( A => n7476, Z => n7475);
   U6325 : INV_X1 port map( A => n5035, ZN => n7578);
   U6326 : OAI21_X1 port map( B1 => n5067, B2 => n5068, A => n7584, ZN => n5035
                           );
   U6327 : INV_X1 port map( A => n7197, ZN => n7206);
   U6328 : AOI221_X1 port map( B1 => n7086, B2 => n5001, C1 => n7083, C2 => 
                           n5033, A => n6393, ZN => n6392);
   U6329 : OAI22_X1 port map( A1 => n4937, A2 => n7080, B1 => n4969, B2 => 
                           n7077, ZN => n6393);
   U6330 : AOI221_X1 port map( B1 => n7038, B2 => n4617, C1 => n7035, C2 => 
                           n4649, A => n6411, ZN => n6410);
   U6331 : OAI22_X1 port map( A1 => n4553, A2 => n7032, B1 => n4585, B2 => 
                           n7029, ZN => n6411);
   U6332 : AOI221_X1 port map( B1 => n7086, B2 => n5000, C1 => n7083, C2 => 
                           n5032, A => n6374, ZN => n6373);
   U6333 : OAI22_X1 port map( A1 => n4936, A2 => n7080, B1 => n4968, B2 => 
                           n7077, ZN => n6374);
   U6334 : AOI221_X1 port map( B1 => n7038, B2 => n4616, C1 => n7035, C2 => 
                           n4648, A => n6382, ZN => n6381);
   U6335 : OAI22_X1 port map( A1 => n4552, A2 => n7032, B1 => n4584, B2 => 
                           n7029, ZN => n6382);
   U6336 : AOI221_X1 port map( B1 => n7086, B2 => n4999, C1 => n7083, C2 => 
                           n5031, A => n6355, ZN => n6354);
   U6337 : OAI22_X1 port map( A1 => n4935, A2 => n7080, B1 => n4967, B2 => 
                           n7077, ZN => n6355);
   U6338 : AOI221_X1 port map( B1 => n7038, B2 => n4615, C1 => n7035, C2 => 
                           n4647, A => n6363, ZN => n6362);
   U6339 : OAI22_X1 port map( A1 => n4551, A2 => n7032, B1 => n4583, B2 => 
                           n7029, ZN => n6363);
   U6340 : AOI221_X1 port map( B1 => n7086, B2 => n4998, C1 => n7083, C2 => 
                           n5030, A => n6336, ZN => n6335);
   U6341 : OAI22_X1 port map( A1 => n4934, A2 => n7080, B1 => n4966, B2 => 
                           n7077, ZN => n6336);
   U6342 : AOI221_X1 port map( B1 => n7038, B2 => n4614, C1 => n7035, C2 => 
                           n4646, A => n6344, ZN => n6343);
   U6343 : OAI22_X1 port map( A1 => n4550, A2 => n7032, B1 => n4582, B2 => 
                           n7029, ZN => n6344);
   U6344 : AOI221_X1 port map( B1 => n7086, B2 => n4997, C1 => n7083, C2 => 
                           n5029, A => n6317, ZN => n6316);
   U6345 : OAI22_X1 port map( A1 => n4933, A2 => n7080, B1 => n4965, B2 => 
                           n7077, ZN => n6317);
   U6346 : AOI221_X1 port map( B1 => n7038, B2 => n4613, C1 => n7035, C2 => 
                           n4645, A => n6325, ZN => n6324);
   U6347 : OAI22_X1 port map( A1 => n4549, A2 => n7032, B1 => n4581, B2 => 
                           n7029, ZN => n6325);
   U6348 : AOI221_X1 port map( B1 => n7086, B2 => n4996, C1 => n7083, C2 => 
                           n5028, A => n6298, ZN => n6297);
   U6349 : OAI22_X1 port map( A1 => n4932, A2 => n7080, B1 => n4964, B2 => 
                           n7077, ZN => n6298);
   U6350 : AOI221_X1 port map( B1 => n7038, B2 => n4612, C1 => n7035, C2 => 
                           n4644, A => n6306, ZN => n6305);
   U6351 : OAI22_X1 port map( A1 => n4548, A2 => n7032, B1 => n4580, B2 => 
                           n7029, ZN => n6306);
   U6352 : AOI221_X1 port map( B1 => n7086, B2 => n4995, C1 => n7083, C2 => 
                           n5027, A => n6279, ZN => n6278);
   U6353 : OAI22_X1 port map( A1 => n4931, A2 => n7080, B1 => n4963, B2 => 
                           n7077, ZN => n6279);
   U6354 : AOI221_X1 port map( B1 => n7038, B2 => n4611, C1 => n7035, C2 => 
                           n4643, A => n6287, ZN => n6286);
   U6355 : OAI22_X1 port map( A1 => n4547, A2 => n7032, B1 => n4579, B2 => 
                           n7029, ZN => n6287);
   U6356 : AOI221_X1 port map( B1 => n7086, B2 => n4994, C1 => n7083, C2 => 
                           n5026, A => n6260, ZN => n6259);
   U6357 : OAI22_X1 port map( A1 => n4930, A2 => n7080, B1 => n4962, B2 => 
                           n7077, ZN => n6260);
   U6358 : AOI221_X1 port map( B1 => n7038, B2 => n4610, C1 => n7035, C2 => 
                           n4642, A => n6268, ZN => n6267);
   U6359 : OAI22_X1 port map( A1 => n4546, A2 => n7032, B1 => n4578, B2 => 
                           n7029, ZN => n6268);
   U6360 : AOI221_X1 port map( B1 => n7086, B2 => n4993, C1 => n7083, C2 => 
                           n5025, A => n6241, ZN => n6240);
   U6361 : OAI22_X1 port map( A1 => n4929, A2 => n7080, B1 => n4961, B2 => 
                           n7077, ZN => n6241);
   U6362 : AOI221_X1 port map( B1 => n7038, B2 => n4609, C1 => n7035, C2 => 
                           n4641, A => n6249, ZN => n6248);
   U6363 : OAI22_X1 port map( A1 => n4545, A2 => n7032, B1 => n4577, B2 => 
                           n7029, ZN => n6249);
   U6364 : AOI221_X1 port map( B1 => n7086, B2 => n4992, C1 => n7083, C2 => 
                           n5024, A => n6222, ZN => n6221);
   U6365 : OAI22_X1 port map( A1 => n4928, A2 => n7080, B1 => n4960, B2 => 
                           n7077, ZN => n6222);
   U6366 : AOI221_X1 port map( B1 => n7038, B2 => n4608, C1 => n7035, C2 => 
                           n4640, A => n6230, ZN => n6229);
   U6367 : OAI22_X1 port map( A1 => n4544, A2 => n7032, B1 => n4576, B2 => 
                           n7029, ZN => n6230);
   U6368 : AOI221_X1 port map( B1 => n7086, B2 => n4991, C1 => n7083, C2 => 
                           n5023, A => n6203, ZN => n6202);
   U6369 : OAI22_X1 port map( A1 => n4927, A2 => n7080, B1 => n4959, B2 => 
                           n7077, ZN => n6203);
   U6370 : AOI221_X1 port map( B1 => n7038, B2 => n4607, C1 => n7035, C2 => 
                           n4639, A => n6211, ZN => n6210);
   U6371 : OAI22_X1 port map( A1 => n4543, A2 => n7032, B1 => n4575, B2 => 
                           n7029, ZN => n6211);
   U6372 : AOI221_X1 port map( B1 => n7086, B2 => n4990, C1 => n7083, C2 => 
                           n5022, A => n6184, ZN => n6183);
   U6373 : OAI22_X1 port map( A1 => n4926, A2 => n7080, B1 => n4958, B2 => 
                           n7077, ZN => n6184);
   U6374 : AOI221_X1 port map( B1 => n7038, B2 => n4606, C1 => n7035, C2 => 
                           n4638, A => n6192, ZN => n6191);
   U6375 : OAI22_X1 port map( A1 => n4542, A2 => n7032, B1 => n4574, B2 => 
                           n7029, ZN => n6192);
   U6376 : AOI221_X1 port map( B1 => n7087, B2 => n4989, C1 => n7084, C2 => 
                           n5021, A => n6165, ZN => n6164);
   U6377 : OAI22_X1 port map( A1 => n4925, A2 => n7081, B1 => n4957, B2 => 
                           n7078, ZN => n6165);
   U6378 : AOI221_X1 port map( B1 => n7039, B2 => n4605, C1 => n7036, C2 => 
                           n4637, A => n6173, ZN => n6172);
   U6379 : OAI22_X1 port map( A1 => n4541, A2 => n7033, B1 => n4573, B2 => 
                           n7030, ZN => n6173);
   U6380 : AOI221_X1 port map( B1 => n7087, B2 => n4988, C1 => n7084, C2 => 
                           n5020, A => n6146, ZN => n6145);
   U6381 : OAI22_X1 port map( A1 => n4924, A2 => n7081, B1 => n4956, B2 => 
                           n7078, ZN => n6146);
   U6382 : AOI221_X1 port map( B1 => n7039, B2 => n4604, C1 => n7036, C2 => 
                           n4636, A => n6154, ZN => n6153);
   U6383 : OAI22_X1 port map( A1 => n4540, A2 => n7033, B1 => n4572, B2 => 
                           n7030, ZN => n6154);
   U6384 : AOI221_X1 port map( B1 => n7087, B2 => n4987, C1 => n7084, C2 => 
                           n5019, A => n6127, ZN => n6126);
   U6385 : OAI22_X1 port map( A1 => n4923, A2 => n7081, B1 => n4955, B2 => 
                           n7078, ZN => n6127);
   U6386 : AOI221_X1 port map( B1 => n7039, B2 => n4603, C1 => n7036, C2 => 
                           n4635, A => n6135, ZN => n6134);
   U6387 : OAI22_X1 port map( A1 => n4539, A2 => n7033, B1 => n4571, B2 => 
                           n7030, ZN => n6135);
   U6388 : AOI221_X1 port map( B1 => n7087, B2 => n4986, C1 => n7084, C2 => 
                           n5018, A => n6108, ZN => n6107);
   U6389 : OAI22_X1 port map( A1 => n4922, A2 => n7081, B1 => n4954, B2 => 
                           n7078, ZN => n6108);
   U6390 : AOI221_X1 port map( B1 => n7039, B2 => n4602, C1 => n7036, C2 => 
                           n4634, A => n6116, ZN => n6115);
   U6391 : OAI22_X1 port map( A1 => n4538, A2 => n7033, B1 => n4570, B2 => 
                           n7030, ZN => n6116);
   U6392 : AOI221_X1 port map( B1 => n7087, B2 => n4985, C1 => n7084, C2 => 
                           n5017, A => n6089, ZN => n6088);
   U6393 : OAI22_X1 port map( A1 => n4921, A2 => n7081, B1 => n4953, B2 => 
                           n7078, ZN => n6089);
   U6394 : AOI221_X1 port map( B1 => n7039, B2 => n4601, C1 => n7036, C2 => 
                           n4633, A => n6097, ZN => n6096);
   U6395 : OAI22_X1 port map( A1 => n4537, A2 => n7033, B1 => n4569, B2 => 
                           n7030, ZN => n6097);
   U6396 : AOI221_X1 port map( B1 => n7087, B2 => n4984, C1 => n7084, C2 => 
                           n5016, A => n6070, ZN => n6069);
   U6397 : OAI22_X1 port map( A1 => n4920, A2 => n7081, B1 => n4952, B2 => 
                           n7078, ZN => n6070);
   U6398 : AOI221_X1 port map( B1 => n7039, B2 => n4600, C1 => n7036, C2 => 
                           n4632, A => n6078, ZN => n6077);
   U6399 : OAI22_X1 port map( A1 => n4536, A2 => n7033, B1 => n4568, B2 => 
                           n7030, ZN => n6078);
   U6400 : AOI221_X1 port map( B1 => n7087, B2 => n4983, C1 => n7084, C2 => 
                           n5015, A => n6051, ZN => n6050);
   U6401 : OAI22_X1 port map( A1 => n4919, A2 => n7081, B1 => n4951, B2 => 
                           n7078, ZN => n6051);
   U6402 : AOI221_X1 port map( B1 => n7039, B2 => n4599, C1 => n7036, C2 => 
                           n4631, A => n6059, ZN => n6058);
   U6403 : OAI22_X1 port map( A1 => n4535, A2 => n7033, B1 => n4567, B2 => 
                           n7030, ZN => n6059);
   U6404 : AOI221_X1 port map( B1 => n7087, B2 => n4982, C1 => n7084, C2 => 
                           n5014, A => n6032, ZN => n6031);
   U6405 : OAI22_X1 port map( A1 => n4918, A2 => n7081, B1 => n4950, B2 => 
                           n7078, ZN => n6032);
   U6406 : AOI221_X1 port map( B1 => n7039, B2 => n4598, C1 => n7036, C2 => 
                           n4630, A => n6040, ZN => n6039);
   U6407 : OAI22_X1 port map( A1 => n4534, A2 => n7033, B1 => n4566, B2 => 
                           n7030, ZN => n6040);
   U6408 : AOI221_X1 port map( B1 => n7087, B2 => n4981, C1 => n7084, C2 => 
                           n5013, A => n6013, ZN => n6012);
   U6409 : OAI22_X1 port map( A1 => n4917, A2 => n7081, B1 => n4949, B2 => 
                           n7078, ZN => n6013);
   U6410 : AOI221_X1 port map( B1 => n7039, B2 => n4597, C1 => n7036, C2 => 
                           n4629, A => n6021, ZN => n6020);
   U6411 : OAI22_X1 port map( A1 => n4533, A2 => n7033, B1 => n4565, B2 => 
                           n7030, ZN => n6021);
   U6412 : AOI221_X1 port map( B1 => n7087, B2 => n4980, C1 => n7084, C2 => 
                           n5012, A => n5994, ZN => n5993);
   U6413 : OAI22_X1 port map( A1 => n4916, A2 => n7081, B1 => n4948, B2 => 
                           n7078, ZN => n5994);
   U6414 : AOI221_X1 port map( B1 => n7039, B2 => n4596, C1 => n7036, C2 => 
                           n4628, A => n6002, ZN => n6001);
   U6415 : OAI22_X1 port map( A1 => n4532, A2 => n7033, B1 => n4564, B2 => 
                           n7030, ZN => n6002);
   U6416 : AOI221_X1 port map( B1 => n7087, B2 => n4979, C1 => n7084, C2 => 
                           n5011, A => n5975, ZN => n5974);
   U6417 : OAI22_X1 port map( A1 => n4915, A2 => n7081, B1 => n4947, B2 => 
                           n7078, ZN => n5975);
   U6418 : AOI221_X1 port map( B1 => n7039, B2 => n4595, C1 => n7036, C2 => 
                           n4627, A => n5983, ZN => n5982);
   U6419 : OAI22_X1 port map( A1 => n4531, A2 => n7033, B1 => n4563, B2 => 
                           n7030, ZN => n5983);
   U6420 : AOI221_X1 port map( B1 => n7087, B2 => n4978, C1 => n7084, C2 => 
                           n5010, A => n5956, ZN => n5955);
   U6421 : OAI22_X1 port map( A1 => n4914, A2 => n7081, B1 => n4946, B2 => 
                           n7078, ZN => n5956);
   U6422 : AOI221_X1 port map( B1 => n7039, B2 => n4594, C1 => n7036, C2 => 
                           n4626, A => n5964, ZN => n5963);
   U6423 : OAI22_X1 port map( A1 => n4530, A2 => n7033, B1 => n4562, B2 => 
                           n7030, ZN => n5964);
   U6424 : AOI221_X1 port map( B1 => n7088, B2 => n4977, C1 => n7085, C2 => 
                           n5009, A => n5937, ZN => n5936);
   U6425 : OAI22_X1 port map( A1 => n4913, A2 => n7082, B1 => n4945, B2 => 
                           n7079, ZN => n5937);
   U6426 : AOI221_X1 port map( B1 => n7040, B2 => n4593, C1 => n7037, C2 => 
                           n4625, A => n5945, ZN => n5944);
   U6427 : OAI22_X1 port map( A1 => n4529, A2 => n7034, B1 => n4561, B2 => 
                           n7031, ZN => n5945);
   U6428 : AOI221_X1 port map( B1 => n7088, B2 => n4976, C1 => n7085, C2 => 
                           n5008, A => n5918, ZN => n5917);
   U6429 : OAI22_X1 port map( A1 => n4912, A2 => n7082, B1 => n4944, B2 => 
                           n7079, ZN => n5918);
   U6430 : AOI221_X1 port map( B1 => n7040, B2 => n4592, C1 => n7037, C2 => 
                           n4624, A => n5926, ZN => n5925);
   U6431 : OAI22_X1 port map( A1 => n4528, A2 => n7034, B1 => n4560, B2 => 
                           n7031, ZN => n5926);
   U6432 : AOI221_X1 port map( B1 => n7088, B2 => n4975, C1 => n7085, C2 => 
                           n5007, A => n5899, ZN => n5898);
   U6433 : OAI22_X1 port map( A1 => n4911, A2 => n7082, B1 => n4943, B2 => 
                           n7079, ZN => n5899);
   U6434 : AOI221_X1 port map( B1 => n7040, B2 => n4591, C1 => n7037, C2 => 
                           n4623, A => n5907, ZN => n5906);
   U6435 : OAI22_X1 port map( A1 => n4527, A2 => n7034, B1 => n4559, B2 => 
                           n7031, ZN => n5907);
   U6436 : AOI221_X1 port map( B1 => n7088, B2 => n4974, C1 => n7085, C2 => 
                           n5006, A => n5880, ZN => n5879);
   U6437 : OAI22_X1 port map( A1 => n4910, A2 => n7082, B1 => n4942, B2 => 
                           n7079, ZN => n5880);
   U6438 : AOI221_X1 port map( B1 => n7040, B2 => n4590, C1 => n7037, C2 => 
                           n4622, A => n5888, ZN => n5887);
   U6439 : OAI22_X1 port map( A1 => n4526, A2 => n7034, B1 => n4558, B2 => 
                           n7031, ZN => n5888);
   U6440 : AOI221_X1 port map( B1 => n7088, B2 => n4973, C1 => n7085, C2 => 
                           n5005, A => n5861, ZN => n5860);
   U6441 : OAI22_X1 port map( A1 => n4909, A2 => n7082, B1 => n4941, B2 => 
                           n7079, ZN => n5861);
   U6442 : AOI221_X1 port map( B1 => n7040, B2 => n4589, C1 => n7037, C2 => 
                           n4621, A => n5869, ZN => n5868);
   U6443 : OAI22_X1 port map( A1 => n4525, A2 => n7034, B1 => n4557, B2 => 
                           n7031, ZN => n5869);
   U6444 : AOI221_X1 port map( B1 => n7088, B2 => n4972, C1 => n7085, C2 => 
                           n5004, A => n5842, ZN => n5841);
   U6445 : OAI22_X1 port map( A1 => n4908, A2 => n7082, B1 => n4940, B2 => 
                           n7079, ZN => n5842);
   U6446 : AOI221_X1 port map( B1 => n7040, B2 => n4588, C1 => n7037, C2 => 
                           n4620, A => n5850, ZN => n5849);
   U6447 : OAI22_X1 port map( A1 => n4524, A2 => n7034, B1 => n4556, B2 => 
                           n7031, ZN => n5850);
   U6448 : AOI221_X1 port map( B1 => n7088, B2 => n4971, C1 => n7085, C2 => 
                           n5003, A => n5823, ZN => n5822);
   U6449 : OAI22_X1 port map( A1 => n4907, A2 => n7082, B1 => n4939, B2 => 
                           n7079, ZN => n5823);
   U6450 : AOI221_X1 port map( B1 => n7040, B2 => n4587, C1 => n7037, C2 => 
                           n4619, A => n5831, ZN => n5830);
   U6451 : OAI22_X1 port map( A1 => n4523, A2 => n7034, B1 => n4555, B2 => 
                           n7031, ZN => n5831);
   U6452 : AOI221_X1 port map( B1 => n7088, B2 => n4970, C1 => n7085, C2 => 
                           n5002, A => n5774, ZN => n5771);
   U6453 : OAI22_X1 port map( A1 => n4906, A2 => n7082, B1 => n4938, B2 => 
                           n7079, ZN => n5774);
   U6454 : AOI221_X1 port map( B1 => n7040, B2 => n4586, C1 => n7037, C2 => 
                           n4618, A => n5798, ZN => n5795);
   U6455 : OAI22_X1 port map( A1 => n4522, A2 => n7034, B1 => n4554, B2 => 
                           n7031, ZN => n5798);
   U6456 : AOI221_X1 port map( B1 => n7188, B2 => n5001, C1 => n7185, C2 => 
                           n5033, A => n5740, ZN => n5739);
   U6457 : OAI22_X1 port map( A1 => n4937, A2 => n7182, B1 => n4969, B2 => 
                           n7179, ZN => n5740);
   U6458 : AOI221_X1 port map( B1 => n7140, B2 => n4617, C1 => n7137, C2 => 
                           n4649, A => n5758, ZN => n5757);
   U6459 : OAI22_X1 port map( A1 => n4553, A2 => n7134, B1 => n4585, B2 => 
                           n7131, ZN => n5758);
   U6460 : AOI221_X1 port map( B1 => n7188, B2 => n5000, C1 => n7185, C2 => 
                           n5032, A => n5721, ZN => n5720);
   U6461 : OAI22_X1 port map( A1 => n4936, A2 => n7182, B1 => n4968, B2 => 
                           n7179, ZN => n5721);
   U6462 : AOI221_X1 port map( B1 => n7140, B2 => n4616, C1 => n7137, C2 => 
                           n4648, A => n5729, ZN => n5728);
   U6463 : OAI22_X1 port map( A1 => n4552, A2 => n7134, B1 => n4584, B2 => 
                           n7131, ZN => n5729);
   U6464 : AOI221_X1 port map( B1 => n7188, B2 => n4999, C1 => n7185, C2 => 
                           n5031, A => n5702, ZN => n5701);
   U6465 : OAI22_X1 port map( A1 => n4935, A2 => n7182, B1 => n4967, B2 => 
                           n7179, ZN => n5702);
   U6466 : AOI221_X1 port map( B1 => n7140, B2 => n4615, C1 => n7137, C2 => 
                           n4647, A => n5710, ZN => n5709);
   U6467 : OAI22_X1 port map( A1 => n4551, A2 => n7134, B1 => n4583, B2 => 
                           n7131, ZN => n5710);
   U6468 : AOI221_X1 port map( B1 => n7188, B2 => n4998, C1 => n7185, C2 => 
                           n5030, A => n5683, ZN => n5682);
   U6469 : OAI22_X1 port map( A1 => n4934, A2 => n7182, B1 => n4966, B2 => 
                           n7179, ZN => n5683);
   U6470 : AOI221_X1 port map( B1 => n7140, B2 => n4614, C1 => n7137, C2 => 
                           n4646, A => n5691, ZN => n5690);
   U6471 : OAI22_X1 port map( A1 => n4550, A2 => n7134, B1 => n4582, B2 => 
                           n7131, ZN => n5691);
   U6472 : AOI221_X1 port map( B1 => n7188, B2 => n4997, C1 => n7185, C2 => 
                           n5029, A => n5664, ZN => n5663);
   U6473 : OAI22_X1 port map( A1 => n4933, A2 => n7182, B1 => n4965, B2 => 
                           n7179, ZN => n5664);
   U6474 : AOI221_X1 port map( B1 => n7140, B2 => n4613, C1 => n7137, C2 => 
                           n4645, A => n5672, ZN => n5671);
   U6475 : OAI22_X1 port map( A1 => n4549, A2 => n7134, B1 => n4581, B2 => 
                           n7131, ZN => n5672);
   U6476 : AOI221_X1 port map( B1 => n7188, B2 => n4996, C1 => n7185, C2 => 
                           n5028, A => n5645, ZN => n5644);
   U6477 : OAI22_X1 port map( A1 => n4932, A2 => n7182, B1 => n4964, B2 => 
                           n7179, ZN => n5645);
   U6478 : AOI221_X1 port map( B1 => n7140, B2 => n4612, C1 => n7137, C2 => 
                           n4644, A => n5653, ZN => n5652);
   U6479 : OAI22_X1 port map( A1 => n4548, A2 => n7134, B1 => n4580, B2 => 
                           n7131, ZN => n5653);
   U6480 : AOI221_X1 port map( B1 => n7188, B2 => n4995, C1 => n7185, C2 => 
                           n5027, A => n5626, ZN => n5625);
   U6481 : OAI22_X1 port map( A1 => n4931, A2 => n7182, B1 => n4963, B2 => 
                           n7179, ZN => n5626);
   U6482 : AOI221_X1 port map( B1 => n7140, B2 => n4611, C1 => n7137, C2 => 
                           n4643, A => n5634, ZN => n5633);
   U6483 : OAI22_X1 port map( A1 => n4547, A2 => n7134, B1 => n4579, B2 => 
                           n7131, ZN => n5634);
   U6484 : AOI221_X1 port map( B1 => n7188, B2 => n4994, C1 => n7185, C2 => 
                           n5026, A => n5607, ZN => n5606);
   U6485 : OAI22_X1 port map( A1 => n4930, A2 => n7182, B1 => n4962, B2 => 
                           n7179, ZN => n5607);
   U6486 : AOI221_X1 port map( B1 => n7140, B2 => n4610, C1 => n7137, C2 => 
                           n4642, A => n5615, ZN => n5614);
   U6487 : OAI22_X1 port map( A1 => n4546, A2 => n7134, B1 => n4578, B2 => 
                           n7131, ZN => n5615);
   U6488 : AOI221_X1 port map( B1 => n7188, B2 => n4993, C1 => n7185, C2 => 
                           n5025, A => n5588, ZN => n5587);
   U6489 : OAI22_X1 port map( A1 => n4929, A2 => n7182, B1 => n4961, B2 => 
                           n7179, ZN => n5588);
   U6490 : AOI221_X1 port map( B1 => n7140, B2 => n4609, C1 => n7137, C2 => 
                           n4641, A => n5596, ZN => n5595);
   U6491 : OAI22_X1 port map( A1 => n4545, A2 => n7134, B1 => n4577, B2 => 
                           n7131, ZN => n5596);
   U6492 : AOI221_X1 port map( B1 => n7188, B2 => n4992, C1 => n7185, C2 => 
                           n5024, A => n5569, ZN => n5568);
   U6493 : OAI22_X1 port map( A1 => n4928, A2 => n7182, B1 => n4960, B2 => 
                           n7179, ZN => n5569);
   U6494 : AOI221_X1 port map( B1 => n7140, B2 => n4608, C1 => n7137, C2 => 
                           n4640, A => n5577, ZN => n5576);
   U6495 : OAI22_X1 port map( A1 => n4544, A2 => n7134, B1 => n4576, B2 => 
                           n7131, ZN => n5577);
   U6496 : AOI221_X1 port map( B1 => n7188, B2 => n4991, C1 => n7185, C2 => 
                           n5023, A => n5550, ZN => n5549);
   U6497 : OAI22_X1 port map( A1 => n4927, A2 => n7182, B1 => n4959, B2 => 
                           n7179, ZN => n5550);
   U6498 : AOI221_X1 port map( B1 => n7140, B2 => n4607, C1 => n7137, C2 => 
                           n4639, A => n5558, ZN => n5557);
   U6499 : OAI22_X1 port map( A1 => n4543, A2 => n7134, B1 => n4575, B2 => 
                           n7131, ZN => n5558);
   U6500 : AOI221_X1 port map( B1 => n7188, B2 => n4990, C1 => n7185, C2 => 
                           n5022, A => n5531, ZN => n5530);
   U6501 : OAI22_X1 port map( A1 => n4926, A2 => n7182, B1 => n4958, B2 => 
                           n7179, ZN => n5531);
   U6502 : AOI221_X1 port map( B1 => n7140, B2 => n4606, C1 => n7137, C2 => 
                           n4638, A => n5539, ZN => n5538);
   U6503 : OAI22_X1 port map( A1 => n4542, A2 => n7134, B1 => n4574, B2 => 
                           n7131, ZN => n5539);
   U6504 : AOI221_X1 port map( B1 => n7189, B2 => n4989, C1 => n7186, C2 => 
                           n5021, A => n5512, ZN => n5511);
   U6505 : OAI22_X1 port map( A1 => n4925, A2 => n7183, B1 => n4957, B2 => 
                           n7180, ZN => n5512);
   U6506 : AOI221_X1 port map( B1 => n7141, B2 => n4605, C1 => n7138, C2 => 
                           n4637, A => n5520, ZN => n5519);
   U6507 : OAI22_X1 port map( A1 => n4541, A2 => n7135, B1 => n4573, B2 => 
                           n7132, ZN => n5520);
   U6508 : AOI221_X1 port map( B1 => n7189, B2 => n4988, C1 => n7186, C2 => 
                           n5020, A => n5493, ZN => n5492);
   U6509 : OAI22_X1 port map( A1 => n4924, A2 => n7183, B1 => n4956, B2 => 
                           n7180, ZN => n5493);
   U6510 : AOI221_X1 port map( B1 => n7141, B2 => n4604, C1 => n7138, C2 => 
                           n4636, A => n5501, ZN => n5500);
   U6511 : OAI22_X1 port map( A1 => n4540, A2 => n7135, B1 => n4572, B2 => 
                           n7132, ZN => n5501);
   U6512 : AOI221_X1 port map( B1 => n7189, B2 => n4987, C1 => n7186, C2 => 
                           n5019, A => n5474, ZN => n5473);
   U6513 : OAI22_X1 port map( A1 => n4923, A2 => n7183, B1 => n4955, B2 => 
                           n7180, ZN => n5474);
   U6514 : AOI221_X1 port map( B1 => n7141, B2 => n4603, C1 => n7138, C2 => 
                           n4635, A => n5482, ZN => n5481);
   U6515 : OAI22_X1 port map( A1 => n4539, A2 => n7135, B1 => n4571, B2 => 
                           n7132, ZN => n5482);
   U6516 : AOI221_X1 port map( B1 => n7189, B2 => n4986, C1 => n7186, C2 => 
                           n5018, A => n5455, ZN => n5454);
   U6517 : OAI22_X1 port map( A1 => n4922, A2 => n7183, B1 => n4954, B2 => 
                           n7180, ZN => n5455);
   U6518 : AOI221_X1 port map( B1 => n7141, B2 => n4602, C1 => n7138, C2 => 
                           n4634, A => n5463, ZN => n5462);
   U6519 : OAI22_X1 port map( A1 => n4538, A2 => n7135, B1 => n4570, B2 => 
                           n7132, ZN => n5463);
   U6520 : AOI221_X1 port map( B1 => n7189, B2 => n4985, C1 => n7186, C2 => 
                           n5017, A => n5436, ZN => n5435);
   U6521 : OAI22_X1 port map( A1 => n4921, A2 => n7183, B1 => n4953, B2 => 
                           n7180, ZN => n5436);
   U6522 : AOI221_X1 port map( B1 => n7141, B2 => n4601, C1 => n7138, C2 => 
                           n4633, A => n5444, ZN => n5443);
   U6523 : OAI22_X1 port map( A1 => n4537, A2 => n7135, B1 => n4569, B2 => 
                           n7132, ZN => n5444);
   U6524 : AOI221_X1 port map( B1 => n7189, B2 => n4984, C1 => n7186, C2 => 
                           n5016, A => n5417, ZN => n5416);
   U6525 : OAI22_X1 port map( A1 => n4920, A2 => n7183, B1 => n4952, B2 => 
                           n7180, ZN => n5417);
   U6526 : AOI221_X1 port map( B1 => n7141, B2 => n4600, C1 => n7138, C2 => 
                           n4632, A => n5425, ZN => n5424);
   U6527 : OAI22_X1 port map( A1 => n4536, A2 => n7135, B1 => n4568, B2 => 
                           n7132, ZN => n5425);
   U6528 : AOI221_X1 port map( B1 => n7189, B2 => n4983, C1 => n7186, C2 => 
                           n5015, A => n5398, ZN => n5397);
   U6529 : OAI22_X1 port map( A1 => n4919, A2 => n7183, B1 => n4951, B2 => 
                           n7180, ZN => n5398);
   U6530 : AOI221_X1 port map( B1 => n7141, B2 => n4599, C1 => n7138, C2 => 
                           n4631, A => n5406, ZN => n5405);
   U6531 : OAI22_X1 port map( A1 => n4535, A2 => n7135, B1 => n4567, B2 => 
                           n7132, ZN => n5406);
   U6532 : AOI221_X1 port map( B1 => n7189, B2 => n4982, C1 => n7186, C2 => 
                           n5014, A => n5379, ZN => n5378);
   U6533 : OAI22_X1 port map( A1 => n4918, A2 => n7183, B1 => n4950, B2 => 
                           n7180, ZN => n5379);
   U6534 : AOI221_X1 port map( B1 => n7141, B2 => n4598, C1 => n7138, C2 => 
                           n4630, A => n5387, ZN => n5386);
   U6535 : OAI22_X1 port map( A1 => n4534, A2 => n7135, B1 => n4566, B2 => 
                           n7132, ZN => n5387);
   U6536 : AOI221_X1 port map( B1 => n7189, B2 => n4981, C1 => n7186, C2 => 
                           n5013, A => n5360, ZN => n5359);
   U6537 : OAI22_X1 port map( A1 => n4917, A2 => n7183, B1 => n4949, B2 => 
                           n7180, ZN => n5360);
   U6538 : AOI221_X1 port map( B1 => n7141, B2 => n4597, C1 => n7138, C2 => 
                           n4629, A => n5368, ZN => n5367);
   U6539 : OAI22_X1 port map( A1 => n4533, A2 => n7135, B1 => n4565, B2 => 
                           n7132, ZN => n5368);
   U6540 : AOI221_X1 port map( B1 => n7189, B2 => n4980, C1 => n7186, C2 => 
                           n5012, A => n5341, ZN => n5340);
   U6541 : OAI22_X1 port map( A1 => n4916, A2 => n7183, B1 => n4948, B2 => 
                           n7180, ZN => n5341);
   U6542 : AOI221_X1 port map( B1 => n7141, B2 => n4596, C1 => n7138, C2 => 
                           n4628, A => n5349, ZN => n5348);
   U6543 : OAI22_X1 port map( A1 => n4532, A2 => n7135, B1 => n4564, B2 => 
                           n7132, ZN => n5349);
   U6544 : AOI221_X1 port map( B1 => n7189, B2 => n4979, C1 => n7186, C2 => 
                           n5011, A => n5322, ZN => n5321);
   U6545 : OAI22_X1 port map( A1 => n4915, A2 => n7183, B1 => n4947, B2 => 
                           n7180, ZN => n5322);
   U6546 : AOI221_X1 port map( B1 => n7141, B2 => n4595, C1 => n7138, C2 => 
                           n4627, A => n5330, ZN => n5329);
   U6547 : OAI22_X1 port map( A1 => n4531, A2 => n7135, B1 => n4563, B2 => 
                           n7132, ZN => n5330);
   U6548 : AOI221_X1 port map( B1 => n7189, B2 => n4978, C1 => n7186, C2 => 
                           n5010, A => n5303, ZN => n5302);
   U6549 : OAI22_X1 port map( A1 => n4914, A2 => n7183, B1 => n4946, B2 => 
                           n7180, ZN => n5303);
   U6550 : AOI221_X1 port map( B1 => n7141, B2 => n4594, C1 => n7138, C2 => 
                           n4626, A => n5311, ZN => n5310);
   U6551 : OAI22_X1 port map( A1 => n4530, A2 => n7135, B1 => n4562, B2 => 
                           n7132, ZN => n5311);
   U6552 : AOI221_X1 port map( B1 => n7190, B2 => n4977, C1 => n7187, C2 => 
                           n5009, A => n5284, ZN => n5283);
   U6553 : OAI22_X1 port map( A1 => n4913, A2 => n7184, B1 => n4945, B2 => 
                           n7181, ZN => n5284);
   U6554 : AOI221_X1 port map( B1 => n7142, B2 => n4593, C1 => n7139, C2 => 
                           n4625, A => n5292, ZN => n5291);
   U6555 : OAI22_X1 port map( A1 => n4529, A2 => n7136, B1 => n4561, B2 => 
                           n7133, ZN => n5292);
   U6556 : AOI221_X1 port map( B1 => n7190, B2 => n4976, C1 => n7187, C2 => 
                           n5008, A => n5265, ZN => n5264);
   U6557 : OAI22_X1 port map( A1 => n4912, A2 => n7184, B1 => n4944, B2 => 
                           n7181, ZN => n5265);
   U6558 : AOI221_X1 port map( B1 => n7142, B2 => n4592, C1 => n7139, C2 => 
                           n4624, A => n5273, ZN => n5272);
   U6559 : OAI22_X1 port map( A1 => n4528, A2 => n7136, B1 => n4560, B2 => 
                           n7133, ZN => n5273);
   U6560 : AOI221_X1 port map( B1 => n7190, B2 => n4975, C1 => n7187, C2 => 
                           n5007, A => n5246, ZN => n5245);
   U6561 : OAI22_X1 port map( A1 => n4911, A2 => n7184, B1 => n4943, B2 => 
                           n7181, ZN => n5246);
   U6562 : AOI221_X1 port map( B1 => n7142, B2 => n4591, C1 => n7139, C2 => 
                           n4623, A => n5254, ZN => n5253);
   U6563 : OAI22_X1 port map( A1 => n4527, A2 => n7136, B1 => n4559, B2 => 
                           n7133, ZN => n5254);
   U6564 : AOI221_X1 port map( B1 => n7190, B2 => n4974, C1 => n7187, C2 => 
                           n5006, A => n5227, ZN => n5226);
   U6565 : OAI22_X1 port map( A1 => n4910, A2 => n7184, B1 => n4942, B2 => 
                           n7181, ZN => n5227);
   U6566 : AOI221_X1 port map( B1 => n7142, B2 => n4590, C1 => n7139, C2 => 
                           n4622, A => n5235, ZN => n5234);
   U6567 : OAI22_X1 port map( A1 => n4526, A2 => n7136, B1 => n4558, B2 => 
                           n7133, ZN => n5235);
   U6568 : AOI221_X1 port map( B1 => n7190, B2 => n4973, C1 => n7187, C2 => 
                           n5005, A => n5208, ZN => n5207);
   U6569 : OAI22_X1 port map( A1 => n4909, A2 => n7184, B1 => n4941, B2 => 
                           n7181, ZN => n5208);
   U6570 : AOI221_X1 port map( B1 => n7142, B2 => n4589, C1 => n7139, C2 => 
                           n4621, A => n5216, ZN => n5215);
   U6571 : OAI22_X1 port map( A1 => n4525, A2 => n7136, B1 => n4557, B2 => 
                           n7133, ZN => n5216);
   U6572 : AOI221_X1 port map( B1 => n7190, B2 => n4972, C1 => n7187, C2 => 
                           n5004, A => n5189, ZN => n5188);
   U6573 : OAI22_X1 port map( A1 => n4908, A2 => n7184, B1 => n4940, B2 => 
                           n7181, ZN => n5189);
   U6574 : AOI221_X1 port map( B1 => n7142, B2 => n4588, C1 => n7139, C2 => 
                           n4620, A => n5197, ZN => n5196);
   U6575 : OAI22_X1 port map( A1 => n4524, A2 => n7136, B1 => n4556, B2 => 
                           n7133, ZN => n5197);
   U6576 : AOI221_X1 port map( B1 => n7190, B2 => n4971, C1 => n7187, C2 => 
                           n5003, A => n5170, ZN => n5169);
   U6577 : OAI22_X1 port map( A1 => n4907, A2 => n7184, B1 => n4939, B2 => 
                           n7181, ZN => n5170);
   U6578 : AOI221_X1 port map( B1 => n7142, B2 => n4587, C1 => n7139, C2 => 
                           n4619, A => n5178, ZN => n5177);
   U6579 : OAI22_X1 port map( A1 => n4523, A2 => n7136, B1 => n4555, B2 => 
                           n7133, ZN => n5178);
   U6580 : AOI221_X1 port map( B1 => n7190, B2 => n4970, C1 => n7187, C2 => 
                           n5002, A => n5121, ZN => n5118);
   U6581 : OAI22_X1 port map( A1 => n4906, A2 => n7184, B1 => n4938, B2 => 
                           n7181, ZN => n5121);
   U6582 : AOI221_X1 port map( B1 => n7142, B2 => n4586, C1 => n7139, C2 => 
                           n4618, A => n5145, ZN => n5142);
   U6583 : OAI22_X1 port map( A1 => n4522, A2 => n7136, B1 => n4554, B2 => 
                           n7133, ZN => n5145);
   U6584 : AOI221_X1 port map( B1 => n7062, B2 => n4809, C1 => n7059, C2 => 
                           n4841, A => n6404, ZN => n6390);
   U6585 : OAI22_X1 port map( A1 => n4745, A2 => n7056, B1 => n4777, B2 => 
                           n7053, ZN => n6404);
   U6586 : AOI221_X1 port map( B1 => n7014, B2 => n4425, C1 => n7011, C2 => 
                           n4457, A => n6414, ZN => n6408);
   U6587 : OAI22_X1 port map( A1 => n4361, A2 => n7008, B1 => n4393, B2 => 
                           n7005, ZN => n6414);
   U6588 : AOI221_X1 port map( B1 => n7062, B2 => n4808, C1 => n7059, C2 => 
                           n4840, A => n6376, ZN => n6371);
   U6589 : OAI22_X1 port map( A1 => n4744, A2 => n7056, B1 => n4776, B2 => 
                           n7053, ZN => n6376);
   U6590 : AOI221_X1 port map( B1 => n7014, B2 => n4424, C1 => n7011, C2 => 
                           n4456, A => n6384, ZN => n6379);
   U6591 : OAI22_X1 port map( A1 => n4360, A2 => n7008, B1 => n4392, B2 => 
                           n7005, ZN => n6384);
   U6592 : AOI221_X1 port map( B1 => n7062, B2 => n4807, C1 => n7059, C2 => 
                           n4839, A => n6357, ZN => n6352);
   U6593 : OAI22_X1 port map( A1 => n4743, A2 => n7056, B1 => n4775, B2 => 
                           n7053, ZN => n6357);
   U6594 : AOI221_X1 port map( B1 => n7014, B2 => n4423, C1 => n7011, C2 => 
                           n4455, A => n6365, ZN => n6360);
   U6595 : OAI22_X1 port map( A1 => n4359, A2 => n7008, B1 => n4391, B2 => 
                           n7005, ZN => n6365);
   U6596 : AOI221_X1 port map( B1 => n7062, B2 => n4806, C1 => n7059, C2 => 
                           n4838, A => n6338, ZN => n6333);
   U6597 : OAI22_X1 port map( A1 => n4742, A2 => n7056, B1 => n4774, B2 => 
                           n7053, ZN => n6338);
   U6598 : AOI221_X1 port map( B1 => n7014, B2 => n4422, C1 => n7011, C2 => 
                           n4454, A => n6346, ZN => n6341);
   U6599 : OAI22_X1 port map( A1 => n4358, A2 => n7008, B1 => n4390, B2 => 
                           n7005, ZN => n6346);
   U6600 : AOI221_X1 port map( B1 => n7062, B2 => n4805, C1 => n7059, C2 => 
                           n4837, A => n6319, ZN => n6314);
   U6601 : OAI22_X1 port map( A1 => n4741, A2 => n7056, B1 => n4773, B2 => 
                           n7053, ZN => n6319);
   U6602 : AOI221_X1 port map( B1 => n7014, B2 => n4421, C1 => n7011, C2 => 
                           n4453, A => n6327, ZN => n6322);
   U6603 : OAI22_X1 port map( A1 => n4357, A2 => n7008, B1 => n4389, B2 => 
                           n7005, ZN => n6327);
   U6604 : AOI221_X1 port map( B1 => n7062, B2 => n4804, C1 => n7059, C2 => 
                           n4836, A => n6300, ZN => n6295);
   U6605 : OAI22_X1 port map( A1 => n4740, A2 => n7056, B1 => n4772, B2 => 
                           n7053, ZN => n6300);
   U6606 : AOI221_X1 port map( B1 => n7014, B2 => n4420, C1 => n7011, C2 => 
                           n4452, A => n6308, ZN => n6303);
   U6607 : OAI22_X1 port map( A1 => n4356, A2 => n7008, B1 => n4388, B2 => 
                           n7005, ZN => n6308);
   U6608 : AOI221_X1 port map( B1 => n7062, B2 => n4803, C1 => n7059, C2 => 
                           n4835, A => n6281, ZN => n6276);
   U6609 : OAI22_X1 port map( A1 => n4739, A2 => n7056, B1 => n4771, B2 => 
                           n7053, ZN => n6281);
   U6610 : AOI221_X1 port map( B1 => n7014, B2 => n4419, C1 => n7011, C2 => 
                           n4451, A => n6289, ZN => n6284);
   U6611 : OAI22_X1 port map( A1 => n4355, A2 => n7008, B1 => n4387, B2 => 
                           n7005, ZN => n6289);
   U6612 : AOI221_X1 port map( B1 => n7062, B2 => n4802, C1 => n7059, C2 => 
                           n4834, A => n6262, ZN => n6257);
   U6613 : OAI22_X1 port map( A1 => n4738, A2 => n7056, B1 => n4770, B2 => 
                           n7053, ZN => n6262);
   U6614 : AOI221_X1 port map( B1 => n7014, B2 => n4418, C1 => n7011, C2 => 
                           n4450, A => n6270, ZN => n6265);
   U6615 : OAI22_X1 port map( A1 => n4354, A2 => n7008, B1 => n4386, B2 => 
                           n7005, ZN => n6270);
   U6616 : AOI221_X1 port map( B1 => n7062, B2 => n4801, C1 => n7059, C2 => 
                           n4833, A => n6243, ZN => n6238);
   U6617 : OAI22_X1 port map( A1 => n4737, A2 => n7056, B1 => n4769, B2 => 
                           n7053, ZN => n6243);
   U6618 : AOI221_X1 port map( B1 => n7014, B2 => n4417, C1 => n7011, C2 => 
                           n4449, A => n6251, ZN => n6246);
   U6619 : OAI22_X1 port map( A1 => n4353, A2 => n7008, B1 => n4385, B2 => 
                           n7005, ZN => n6251);
   U6620 : AOI221_X1 port map( B1 => n7062, B2 => n4800, C1 => n7059, C2 => 
                           n4832, A => n6224, ZN => n6219);
   U6621 : OAI22_X1 port map( A1 => n4736, A2 => n7056, B1 => n4768, B2 => 
                           n7053, ZN => n6224);
   U6622 : AOI221_X1 port map( B1 => n7014, B2 => n4416, C1 => n7011, C2 => 
                           n4448, A => n6232, ZN => n6227);
   U6623 : OAI22_X1 port map( A1 => n4352, A2 => n7008, B1 => n4384, B2 => 
                           n7005, ZN => n6232);
   U6624 : AOI221_X1 port map( B1 => n7062, B2 => n4799, C1 => n7059, C2 => 
                           n4831, A => n6205, ZN => n6200);
   U6625 : OAI22_X1 port map( A1 => n4735, A2 => n7056, B1 => n4767, B2 => 
                           n7053, ZN => n6205);
   U6626 : AOI221_X1 port map( B1 => n7014, B2 => n4415, C1 => n7011, C2 => 
                           n4447, A => n6213, ZN => n6208);
   U6627 : OAI22_X1 port map( A1 => n4351, A2 => n7008, B1 => n4383, B2 => 
                           n7005, ZN => n6213);
   U6628 : AOI221_X1 port map( B1 => n7062, B2 => n4798, C1 => n7059, C2 => 
                           n4830, A => n6186, ZN => n6181);
   U6629 : OAI22_X1 port map( A1 => n4734, A2 => n7056, B1 => n4766, B2 => 
                           n7053, ZN => n6186);
   U6630 : AOI221_X1 port map( B1 => n7014, B2 => n4414, C1 => n7011, C2 => 
                           n4446, A => n6194, ZN => n6189);
   U6631 : OAI22_X1 port map( A1 => n4350, A2 => n7008, B1 => n4382, B2 => 
                           n7005, ZN => n6194);
   U6632 : AOI221_X1 port map( B1 => n7063, B2 => n4797, C1 => n7060, C2 => 
                           n4829, A => n6167, ZN => n6162);
   U6633 : OAI22_X1 port map( A1 => n4733, A2 => n7057, B1 => n4765, B2 => 
                           n7054, ZN => n6167);
   U6634 : AOI221_X1 port map( B1 => n7015, B2 => n4413, C1 => n7012, C2 => 
                           n4445, A => n6175, ZN => n6170);
   U6635 : OAI22_X1 port map( A1 => n4349, A2 => n7009, B1 => n4381, B2 => 
                           n7006, ZN => n6175);
   U6636 : AOI221_X1 port map( B1 => n7063, B2 => n4796, C1 => n7060, C2 => 
                           n4828, A => n6148, ZN => n6143);
   U6637 : OAI22_X1 port map( A1 => n4732, A2 => n7057, B1 => n4764, B2 => 
                           n7054, ZN => n6148);
   U6638 : AOI221_X1 port map( B1 => n7015, B2 => n4412, C1 => n7012, C2 => 
                           n4444, A => n6156, ZN => n6151);
   U6639 : OAI22_X1 port map( A1 => n4348, A2 => n7009, B1 => n4380, B2 => 
                           n7006, ZN => n6156);
   U6640 : AOI221_X1 port map( B1 => n7063, B2 => n4795, C1 => n7060, C2 => 
                           n4827, A => n6129, ZN => n6124);
   U6641 : OAI22_X1 port map( A1 => n4731, A2 => n7057, B1 => n4763, B2 => 
                           n7054, ZN => n6129);
   U6642 : AOI221_X1 port map( B1 => n7015, B2 => n4411, C1 => n7012, C2 => 
                           n4443, A => n6137, ZN => n6132);
   U6643 : OAI22_X1 port map( A1 => n4347, A2 => n7009, B1 => n4379, B2 => 
                           n7006, ZN => n6137);
   U6644 : AOI221_X1 port map( B1 => n7063, B2 => n4794, C1 => n7060, C2 => 
                           n4826, A => n6110, ZN => n6105);
   U6645 : OAI22_X1 port map( A1 => n4730, A2 => n7057, B1 => n4762, B2 => 
                           n7054, ZN => n6110);
   U6646 : AOI221_X1 port map( B1 => n7015, B2 => n4410, C1 => n7012, C2 => 
                           n4442, A => n6118, ZN => n6113);
   U6647 : OAI22_X1 port map( A1 => n4346, A2 => n7009, B1 => n4378, B2 => 
                           n7006, ZN => n6118);
   U6648 : AOI221_X1 port map( B1 => n7063, B2 => n4793, C1 => n7060, C2 => 
                           n4825, A => n6091, ZN => n6086);
   U6649 : OAI22_X1 port map( A1 => n4729, A2 => n7057, B1 => n4761, B2 => 
                           n7054, ZN => n6091);
   U6650 : AOI221_X1 port map( B1 => n7015, B2 => n4409, C1 => n7012, C2 => 
                           n4441, A => n6099, ZN => n6094);
   U6651 : OAI22_X1 port map( A1 => n4345, A2 => n7009, B1 => n4377, B2 => 
                           n7006, ZN => n6099);
   U6652 : AOI221_X1 port map( B1 => n7063, B2 => n4792, C1 => n7060, C2 => 
                           n4824, A => n6072, ZN => n6067);
   U6653 : OAI22_X1 port map( A1 => n4728, A2 => n7057, B1 => n4760, B2 => 
                           n7054, ZN => n6072);
   U6654 : AOI221_X1 port map( B1 => n7015, B2 => n4408, C1 => n7012, C2 => 
                           n4440, A => n6080, ZN => n6075);
   U6655 : OAI22_X1 port map( A1 => n4344, A2 => n7009, B1 => n4376, B2 => 
                           n7006, ZN => n6080);
   U6656 : AOI221_X1 port map( B1 => n7063, B2 => n4791, C1 => n7060, C2 => 
                           n4823, A => n6053, ZN => n6048);
   U6657 : OAI22_X1 port map( A1 => n4727, A2 => n7057, B1 => n4759, B2 => 
                           n7054, ZN => n6053);
   U6658 : AOI221_X1 port map( B1 => n7015, B2 => n4407, C1 => n7012, C2 => 
                           n4439, A => n6061, ZN => n6056);
   U6659 : OAI22_X1 port map( A1 => n4343, A2 => n7009, B1 => n4375, B2 => 
                           n7006, ZN => n6061);
   U6660 : AOI221_X1 port map( B1 => n7063, B2 => n4790, C1 => n7060, C2 => 
                           n4822, A => n6034, ZN => n6029);
   U6661 : OAI22_X1 port map( A1 => n4726, A2 => n7057, B1 => n4758, B2 => 
                           n7054, ZN => n6034);
   U6662 : AOI221_X1 port map( B1 => n7015, B2 => n4406, C1 => n7012, C2 => 
                           n4438, A => n6042, ZN => n6037);
   U6663 : OAI22_X1 port map( A1 => n4342, A2 => n7009, B1 => n4374, B2 => 
                           n7006, ZN => n6042);
   U6664 : AOI221_X1 port map( B1 => n7063, B2 => n4789, C1 => n7060, C2 => 
                           n4821, A => n6015, ZN => n6010);
   U6665 : OAI22_X1 port map( A1 => n4725, A2 => n7057, B1 => n4757, B2 => 
                           n7054, ZN => n6015);
   U6666 : AOI221_X1 port map( B1 => n7015, B2 => n4405, C1 => n7012, C2 => 
                           n4437, A => n6023, ZN => n6018);
   U6667 : OAI22_X1 port map( A1 => n4341, A2 => n7009, B1 => n4373, B2 => 
                           n7006, ZN => n6023);
   U6668 : AOI221_X1 port map( B1 => n7063, B2 => n4788, C1 => n7060, C2 => 
                           n4820, A => n5996, ZN => n5991);
   U6669 : OAI22_X1 port map( A1 => n4724, A2 => n7057, B1 => n4756, B2 => 
                           n7054, ZN => n5996);
   U6670 : AOI221_X1 port map( B1 => n7015, B2 => n4404, C1 => n7012, C2 => 
                           n4436, A => n6004, ZN => n5999);
   U6671 : OAI22_X1 port map( A1 => n4340, A2 => n7009, B1 => n4372, B2 => 
                           n7006, ZN => n6004);
   U6672 : AOI221_X1 port map( B1 => n7063, B2 => n4787, C1 => n7060, C2 => 
                           n4819, A => n5977, ZN => n5972);
   U6673 : OAI22_X1 port map( A1 => n4723, A2 => n7057, B1 => n4755, B2 => 
                           n7054, ZN => n5977);
   U6674 : AOI221_X1 port map( B1 => n7015, B2 => n4403, C1 => n7012, C2 => 
                           n4435, A => n5985, ZN => n5980);
   U6675 : OAI22_X1 port map( A1 => n4339, A2 => n7009, B1 => n4371, B2 => 
                           n7006, ZN => n5985);
   U6676 : AOI221_X1 port map( B1 => n7063, B2 => n4786, C1 => n7060, C2 => 
                           n4818, A => n5958, ZN => n5953);
   U6677 : OAI22_X1 port map( A1 => n4722, A2 => n7057, B1 => n4754, B2 => 
                           n7054, ZN => n5958);
   U6678 : AOI221_X1 port map( B1 => n7015, B2 => n4402, C1 => n7012, C2 => 
                           n4434, A => n5966, ZN => n5961);
   U6679 : OAI22_X1 port map( A1 => n4338, A2 => n7009, B1 => n4370, B2 => 
                           n7006, ZN => n5966);
   U6680 : AOI221_X1 port map( B1 => n7064, B2 => n4785, C1 => n7061, C2 => 
                           n4817, A => n5939, ZN => n5934);
   U6681 : OAI22_X1 port map( A1 => n4721, A2 => n7058, B1 => n4753, B2 => 
                           n7055, ZN => n5939);
   U6682 : AOI221_X1 port map( B1 => n7016, B2 => n4401, C1 => n7013, C2 => 
                           n4433, A => n5947, ZN => n5942);
   U6683 : OAI22_X1 port map( A1 => n4337, A2 => n7010, B1 => n4369, B2 => 
                           n7007, ZN => n5947);
   U6684 : AOI221_X1 port map( B1 => n7064, B2 => n4784, C1 => n7061, C2 => 
                           n4816, A => n5920, ZN => n5915);
   U6685 : OAI22_X1 port map( A1 => n4720, A2 => n7058, B1 => n4752, B2 => 
                           n7055, ZN => n5920);
   U6686 : AOI221_X1 port map( B1 => n7016, B2 => n4400, C1 => n7013, C2 => 
                           n4432, A => n5928, ZN => n5923);
   U6687 : OAI22_X1 port map( A1 => n4336, A2 => n7010, B1 => n4368, B2 => 
                           n7007, ZN => n5928);
   U6688 : AOI221_X1 port map( B1 => n7064, B2 => n4783, C1 => n7061, C2 => 
                           n4815, A => n5901, ZN => n5896);
   U6689 : OAI22_X1 port map( A1 => n4719, A2 => n7058, B1 => n4751, B2 => 
                           n7055, ZN => n5901);
   U6690 : AOI221_X1 port map( B1 => n7016, B2 => n4399, C1 => n7013, C2 => 
                           n4431, A => n5909, ZN => n5904);
   U6691 : OAI22_X1 port map( A1 => n4335, A2 => n7010, B1 => n4367, B2 => 
                           n7007, ZN => n5909);
   U6692 : AOI221_X1 port map( B1 => n7064, B2 => n4782, C1 => n7061, C2 => 
                           n4814, A => n5882, ZN => n5877);
   U6693 : OAI22_X1 port map( A1 => n4718, A2 => n7058, B1 => n4750, B2 => 
                           n7055, ZN => n5882);
   U6694 : AOI221_X1 port map( B1 => n7016, B2 => n4398, C1 => n7013, C2 => 
                           n4430, A => n5890, ZN => n5885);
   U6695 : OAI22_X1 port map( A1 => n4334, A2 => n7010, B1 => n4366, B2 => 
                           n7007, ZN => n5890);
   U6696 : AOI221_X1 port map( B1 => n7064, B2 => n4781, C1 => n7061, C2 => 
                           n4813, A => n5863, ZN => n5858);
   U6697 : OAI22_X1 port map( A1 => n4717, A2 => n7058, B1 => n4749, B2 => 
                           n7055, ZN => n5863);
   U6698 : AOI221_X1 port map( B1 => n7016, B2 => n4397, C1 => n7013, C2 => 
                           n4429, A => n5871, ZN => n5866);
   U6699 : OAI22_X1 port map( A1 => n4333, A2 => n7010, B1 => n4365, B2 => 
                           n7007, ZN => n5871);
   U6700 : AOI221_X1 port map( B1 => n7064, B2 => n4780, C1 => n7061, C2 => 
                           n4812, A => n5844, ZN => n5839);
   U6701 : OAI22_X1 port map( A1 => n4716, A2 => n7058, B1 => n4748, B2 => 
                           n7055, ZN => n5844);
   U6702 : AOI221_X1 port map( B1 => n7016, B2 => n4396, C1 => n7013, C2 => 
                           n4428, A => n5852, ZN => n5847);
   U6703 : OAI22_X1 port map( A1 => n4332, A2 => n7010, B1 => n4364, B2 => 
                           n7007, ZN => n5852);
   U6704 : AOI221_X1 port map( B1 => n7064, B2 => n4779, C1 => n7061, C2 => 
                           n4811, A => n5825, ZN => n5820);
   U6705 : OAI22_X1 port map( A1 => n4715, A2 => n7058, B1 => n4747, B2 => 
                           n7055, ZN => n5825);
   U6706 : AOI221_X1 port map( B1 => n7016, B2 => n4395, C1 => n7013, C2 => 
                           n4427, A => n5833, ZN => n5828);
   U6707 : OAI22_X1 port map( A1 => n4331, A2 => n7010, B1 => n4363, B2 => 
                           n7007, ZN => n5833);
   U6708 : AOI221_X1 port map( B1 => n7064, B2 => n4778, C1 => n7061, C2 => 
                           n4810, A => n5784, ZN => n5769);
   U6709 : OAI22_X1 port map( A1 => n4714, A2 => n7058, B1 => n4746, B2 => 
                           n7055, ZN => n5784);
   U6710 : AOI221_X1 port map( B1 => n7016, B2 => n4394, C1 => n7013, C2 => 
                           n4426, A => n5808, ZN => n5793);
   U6711 : OAI22_X1 port map( A1 => n4330, A2 => n7010, B1 => n4362, B2 => 
                           n7007, ZN => n5808);
   U6712 : AOI221_X1 port map( B1 => n7164, B2 => n4809, C1 => n7161, C2 => 
                           n4841, A => n5751, ZN => n5737);
   U6713 : OAI22_X1 port map( A1 => n4745, A2 => n7158, B1 => n4777, B2 => 
                           n7155, ZN => n5751);
   U6714 : AOI221_X1 port map( B1 => n7116, B2 => n4425, C1 => n7113, C2 => 
                           n4457, A => n5761, ZN => n5755);
   U6715 : OAI22_X1 port map( A1 => n4361, A2 => n7110, B1 => n4393, B2 => 
                           n7107, ZN => n5761);
   U6716 : AOI221_X1 port map( B1 => n7164, B2 => n4808, C1 => n7161, C2 => 
                           n4840, A => n5723, ZN => n5718);
   U6717 : OAI22_X1 port map( A1 => n4744, A2 => n7158, B1 => n4776, B2 => 
                           n7155, ZN => n5723);
   U6718 : AOI221_X1 port map( B1 => n7116, B2 => n4424, C1 => n7113, C2 => 
                           n4456, A => n5731, ZN => n5726);
   U6719 : OAI22_X1 port map( A1 => n4360, A2 => n7110, B1 => n4392, B2 => 
                           n7107, ZN => n5731);
   U6720 : AOI221_X1 port map( B1 => n7164, B2 => n4807, C1 => n7161, C2 => 
                           n4839, A => n5704, ZN => n5699);
   U6721 : OAI22_X1 port map( A1 => n4743, A2 => n7158, B1 => n4775, B2 => 
                           n7155, ZN => n5704);
   U6722 : AOI221_X1 port map( B1 => n7116, B2 => n4423, C1 => n7113, C2 => 
                           n4455, A => n5712, ZN => n5707);
   U6723 : OAI22_X1 port map( A1 => n4359, A2 => n7110, B1 => n4391, B2 => 
                           n7107, ZN => n5712);
   U6724 : AOI221_X1 port map( B1 => n7164, B2 => n4806, C1 => n7161, C2 => 
                           n4838, A => n5685, ZN => n5680);
   U6725 : OAI22_X1 port map( A1 => n4742, A2 => n7158, B1 => n4774, B2 => 
                           n7155, ZN => n5685);
   U6726 : AOI221_X1 port map( B1 => n7116, B2 => n4422, C1 => n7113, C2 => 
                           n4454, A => n5693, ZN => n5688);
   U6727 : OAI22_X1 port map( A1 => n4358, A2 => n7110, B1 => n4390, B2 => 
                           n7107, ZN => n5693);
   U6728 : AOI221_X1 port map( B1 => n7164, B2 => n4805, C1 => n7161, C2 => 
                           n4837, A => n5666, ZN => n5661);
   U6729 : OAI22_X1 port map( A1 => n4741, A2 => n7158, B1 => n4773, B2 => 
                           n7155, ZN => n5666);
   U6730 : AOI221_X1 port map( B1 => n7116, B2 => n4421, C1 => n7113, C2 => 
                           n4453, A => n5674, ZN => n5669);
   U6731 : OAI22_X1 port map( A1 => n4357, A2 => n7110, B1 => n4389, B2 => 
                           n7107, ZN => n5674);
   U6732 : AOI221_X1 port map( B1 => n7164, B2 => n4804, C1 => n7161, C2 => 
                           n4836, A => n5647, ZN => n5642);
   U6733 : OAI22_X1 port map( A1 => n4740, A2 => n7158, B1 => n4772, B2 => 
                           n7155, ZN => n5647);
   U6734 : AOI221_X1 port map( B1 => n7116, B2 => n4420, C1 => n7113, C2 => 
                           n4452, A => n5655, ZN => n5650);
   U6735 : OAI22_X1 port map( A1 => n4356, A2 => n7110, B1 => n4388, B2 => 
                           n7107, ZN => n5655);
   U6736 : AOI221_X1 port map( B1 => n7164, B2 => n4803, C1 => n7161, C2 => 
                           n4835, A => n5628, ZN => n5623);
   U6737 : OAI22_X1 port map( A1 => n4739, A2 => n7158, B1 => n4771, B2 => 
                           n7155, ZN => n5628);
   U6738 : AOI221_X1 port map( B1 => n7116, B2 => n4419, C1 => n7113, C2 => 
                           n4451, A => n5636, ZN => n5631);
   U6739 : OAI22_X1 port map( A1 => n4355, A2 => n7110, B1 => n4387, B2 => 
                           n7107, ZN => n5636);
   U6740 : AOI221_X1 port map( B1 => n7164, B2 => n4802, C1 => n7161, C2 => 
                           n4834, A => n5609, ZN => n5604);
   U6741 : OAI22_X1 port map( A1 => n4738, A2 => n7158, B1 => n4770, B2 => 
                           n7155, ZN => n5609);
   U6742 : AOI221_X1 port map( B1 => n7116, B2 => n4418, C1 => n7113, C2 => 
                           n4450, A => n5617, ZN => n5612);
   U6743 : OAI22_X1 port map( A1 => n4354, A2 => n7110, B1 => n4386, B2 => 
                           n7107, ZN => n5617);
   U6744 : AOI221_X1 port map( B1 => n7164, B2 => n4801, C1 => n7161, C2 => 
                           n4833, A => n5590, ZN => n5585);
   U6745 : OAI22_X1 port map( A1 => n4737, A2 => n7158, B1 => n4769, B2 => 
                           n7155, ZN => n5590);
   U6746 : AOI221_X1 port map( B1 => n7116, B2 => n4417, C1 => n7113, C2 => 
                           n4449, A => n5598, ZN => n5593);
   U6747 : OAI22_X1 port map( A1 => n4353, A2 => n7110, B1 => n4385, B2 => 
                           n7107, ZN => n5598);
   U6748 : AOI221_X1 port map( B1 => n7164, B2 => n4800, C1 => n7161, C2 => 
                           n4832, A => n5571, ZN => n5566);
   U6749 : OAI22_X1 port map( A1 => n4736, A2 => n7158, B1 => n4768, B2 => 
                           n7155, ZN => n5571);
   U6750 : AOI221_X1 port map( B1 => n7116, B2 => n4416, C1 => n7113, C2 => 
                           n4448, A => n5579, ZN => n5574);
   U6751 : OAI22_X1 port map( A1 => n4352, A2 => n7110, B1 => n4384, B2 => 
                           n7107, ZN => n5579);
   U6752 : AOI221_X1 port map( B1 => n7164, B2 => n4799, C1 => n7161, C2 => 
                           n4831, A => n5552, ZN => n5547);
   U6753 : OAI22_X1 port map( A1 => n4735, A2 => n7158, B1 => n4767, B2 => 
                           n7155, ZN => n5552);
   U6754 : AOI221_X1 port map( B1 => n7116, B2 => n4415, C1 => n7113, C2 => 
                           n4447, A => n5560, ZN => n5555);
   U6755 : OAI22_X1 port map( A1 => n4351, A2 => n7110, B1 => n4383, B2 => 
                           n7107, ZN => n5560);
   U6756 : AOI221_X1 port map( B1 => n7164, B2 => n4798, C1 => n7161, C2 => 
                           n4830, A => n5533, ZN => n5528);
   U6757 : OAI22_X1 port map( A1 => n4734, A2 => n7158, B1 => n4766, B2 => 
                           n7155, ZN => n5533);
   U6758 : AOI221_X1 port map( B1 => n7116, B2 => n4414, C1 => n7113, C2 => 
                           n4446, A => n5541, ZN => n5536);
   U6759 : OAI22_X1 port map( A1 => n4350, A2 => n7110, B1 => n4382, B2 => 
                           n7107, ZN => n5541);
   U6760 : AOI221_X1 port map( B1 => n7165, B2 => n4797, C1 => n7162, C2 => 
                           n4829, A => n5514, ZN => n5509);
   U6761 : OAI22_X1 port map( A1 => n4733, A2 => n7159, B1 => n4765, B2 => 
                           n7156, ZN => n5514);
   U6762 : AOI221_X1 port map( B1 => n7117, B2 => n4413, C1 => n7114, C2 => 
                           n4445, A => n5522, ZN => n5517);
   U6763 : OAI22_X1 port map( A1 => n4349, A2 => n7111, B1 => n4381, B2 => 
                           n7108, ZN => n5522);
   U6764 : AOI221_X1 port map( B1 => n7165, B2 => n4796, C1 => n7162, C2 => 
                           n4828, A => n5495, ZN => n5490);
   U6765 : OAI22_X1 port map( A1 => n4732, A2 => n7159, B1 => n4764, B2 => 
                           n7156, ZN => n5495);
   U6766 : AOI221_X1 port map( B1 => n7117, B2 => n4412, C1 => n7114, C2 => 
                           n4444, A => n5503, ZN => n5498);
   U6767 : OAI22_X1 port map( A1 => n4348, A2 => n7111, B1 => n4380, B2 => 
                           n7108, ZN => n5503);
   U6768 : AOI221_X1 port map( B1 => n7165, B2 => n4795, C1 => n7162, C2 => 
                           n4827, A => n5476, ZN => n5471);
   U6769 : OAI22_X1 port map( A1 => n4731, A2 => n7159, B1 => n4763, B2 => 
                           n7156, ZN => n5476);
   U6770 : AOI221_X1 port map( B1 => n7117, B2 => n4411, C1 => n7114, C2 => 
                           n4443, A => n5484, ZN => n5479);
   U6771 : OAI22_X1 port map( A1 => n4347, A2 => n7111, B1 => n4379, B2 => 
                           n7108, ZN => n5484);
   U6772 : AOI221_X1 port map( B1 => n7165, B2 => n4794, C1 => n7162, C2 => 
                           n4826, A => n5457, ZN => n5452);
   U6773 : OAI22_X1 port map( A1 => n4730, A2 => n7159, B1 => n4762, B2 => 
                           n7156, ZN => n5457);
   U6774 : AOI221_X1 port map( B1 => n7117, B2 => n4410, C1 => n7114, C2 => 
                           n4442, A => n5465, ZN => n5460);
   U6775 : OAI22_X1 port map( A1 => n4346, A2 => n7111, B1 => n4378, B2 => 
                           n7108, ZN => n5465);
   U6776 : AOI221_X1 port map( B1 => n7165, B2 => n4793, C1 => n7162, C2 => 
                           n4825, A => n5438, ZN => n5433);
   U6777 : OAI22_X1 port map( A1 => n4729, A2 => n7159, B1 => n4761, B2 => 
                           n7156, ZN => n5438);
   U6778 : AOI221_X1 port map( B1 => n7117, B2 => n4409, C1 => n7114, C2 => 
                           n4441, A => n5446, ZN => n5441);
   U6779 : OAI22_X1 port map( A1 => n4345, A2 => n7111, B1 => n4377, B2 => 
                           n7108, ZN => n5446);
   U6780 : AOI221_X1 port map( B1 => n7165, B2 => n4792, C1 => n7162, C2 => 
                           n4824, A => n5419, ZN => n5414);
   U6781 : OAI22_X1 port map( A1 => n4728, A2 => n7159, B1 => n4760, B2 => 
                           n7156, ZN => n5419);
   U6782 : AOI221_X1 port map( B1 => n7117, B2 => n4408, C1 => n7114, C2 => 
                           n4440, A => n5427, ZN => n5422);
   U6783 : OAI22_X1 port map( A1 => n4344, A2 => n7111, B1 => n4376, B2 => 
                           n7108, ZN => n5427);
   U6784 : AOI221_X1 port map( B1 => n7165, B2 => n4791, C1 => n7162, C2 => 
                           n4823, A => n5400, ZN => n5395);
   U6785 : OAI22_X1 port map( A1 => n4727, A2 => n7159, B1 => n4759, B2 => 
                           n7156, ZN => n5400);
   U6786 : AOI221_X1 port map( B1 => n7117, B2 => n4407, C1 => n7114, C2 => 
                           n4439, A => n5408, ZN => n5403);
   U6787 : OAI22_X1 port map( A1 => n4343, A2 => n7111, B1 => n4375, B2 => 
                           n7108, ZN => n5408);
   U6788 : AOI221_X1 port map( B1 => n7165, B2 => n4790, C1 => n7162, C2 => 
                           n4822, A => n5381, ZN => n5376);
   U6789 : OAI22_X1 port map( A1 => n4726, A2 => n7159, B1 => n4758, B2 => 
                           n7156, ZN => n5381);
   U6790 : AOI221_X1 port map( B1 => n7117, B2 => n4406, C1 => n7114, C2 => 
                           n4438, A => n5389, ZN => n5384);
   U6791 : OAI22_X1 port map( A1 => n4342, A2 => n7111, B1 => n4374, B2 => 
                           n7108, ZN => n5389);
   U6792 : AOI221_X1 port map( B1 => n7165, B2 => n4789, C1 => n7162, C2 => 
                           n4821, A => n5362, ZN => n5357);
   U6793 : OAI22_X1 port map( A1 => n4725, A2 => n7159, B1 => n4757, B2 => 
                           n7156, ZN => n5362);
   U6794 : AOI221_X1 port map( B1 => n7117, B2 => n4405, C1 => n7114, C2 => 
                           n4437, A => n5370, ZN => n5365);
   U6795 : OAI22_X1 port map( A1 => n4341, A2 => n7111, B1 => n4373, B2 => 
                           n7108, ZN => n5370);
   U6796 : AOI221_X1 port map( B1 => n7165, B2 => n4788, C1 => n7162, C2 => 
                           n4820, A => n5343, ZN => n5338);
   U6797 : OAI22_X1 port map( A1 => n4724, A2 => n7159, B1 => n4756, B2 => 
                           n7156, ZN => n5343);
   U6798 : AOI221_X1 port map( B1 => n7117, B2 => n4404, C1 => n7114, C2 => 
                           n4436, A => n5351, ZN => n5346);
   U6799 : OAI22_X1 port map( A1 => n4340, A2 => n7111, B1 => n4372, B2 => 
                           n7108, ZN => n5351);
   U6800 : AOI221_X1 port map( B1 => n7165, B2 => n4787, C1 => n7162, C2 => 
                           n4819, A => n5324, ZN => n5319);
   U6801 : OAI22_X1 port map( A1 => n4723, A2 => n7159, B1 => n4755, B2 => 
                           n7156, ZN => n5324);
   U6802 : AOI221_X1 port map( B1 => n7117, B2 => n4403, C1 => n7114, C2 => 
                           n4435, A => n5332, ZN => n5327);
   U6803 : OAI22_X1 port map( A1 => n4339, A2 => n7111, B1 => n4371, B2 => 
                           n7108, ZN => n5332);
   U6804 : AOI221_X1 port map( B1 => n7165, B2 => n4786, C1 => n7162, C2 => 
                           n4818, A => n5305, ZN => n5300);
   U6805 : OAI22_X1 port map( A1 => n4722, A2 => n7159, B1 => n4754, B2 => 
                           n7156, ZN => n5305);
   U6806 : AOI221_X1 port map( B1 => n7117, B2 => n4402, C1 => n7114, C2 => 
                           n4434, A => n5313, ZN => n5308);
   U6807 : OAI22_X1 port map( A1 => n4338, A2 => n7111, B1 => n4370, B2 => 
                           n7108, ZN => n5313);
   U6808 : AOI221_X1 port map( B1 => n7166, B2 => n4785, C1 => n7163, C2 => 
                           n4817, A => n5286, ZN => n5281);
   U6809 : OAI22_X1 port map( A1 => n4721, A2 => n7160, B1 => n4753, B2 => 
                           n7157, ZN => n5286);
   U6810 : AOI221_X1 port map( B1 => n7118, B2 => n4401, C1 => n7115, C2 => 
                           n4433, A => n5294, ZN => n5289);
   U6811 : OAI22_X1 port map( A1 => n4337, A2 => n7112, B1 => n4369, B2 => 
                           n7109, ZN => n5294);
   U6812 : AOI221_X1 port map( B1 => n7166, B2 => n4784, C1 => n7163, C2 => 
                           n4816, A => n5267, ZN => n5262);
   U6813 : OAI22_X1 port map( A1 => n4720, A2 => n7160, B1 => n4752, B2 => 
                           n7157, ZN => n5267);
   U6814 : AOI221_X1 port map( B1 => n7118, B2 => n4400, C1 => n7115, C2 => 
                           n4432, A => n5275, ZN => n5270);
   U6815 : OAI22_X1 port map( A1 => n4336, A2 => n7112, B1 => n4368, B2 => 
                           n7109, ZN => n5275);
   U6816 : AOI221_X1 port map( B1 => n7166, B2 => n4783, C1 => n7163, C2 => 
                           n4815, A => n5248, ZN => n5243);
   U6817 : OAI22_X1 port map( A1 => n4719, A2 => n7160, B1 => n4751, B2 => 
                           n7157, ZN => n5248);
   U6818 : AOI221_X1 port map( B1 => n7118, B2 => n4399, C1 => n7115, C2 => 
                           n4431, A => n5256, ZN => n5251);
   U6819 : OAI22_X1 port map( A1 => n4335, A2 => n7112, B1 => n4367, B2 => 
                           n7109, ZN => n5256);
   U6820 : AOI221_X1 port map( B1 => n7166, B2 => n4782, C1 => n7163, C2 => 
                           n4814, A => n5229, ZN => n5224);
   U6821 : OAI22_X1 port map( A1 => n4718, A2 => n7160, B1 => n4750, B2 => 
                           n7157, ZN => n5229);
   U6822 : AOI221_X1 port map( B1 => n7118, B2 => n4398, C1 => n7115, C2 => 
                           n4430, A => n5237, ZN => n5232);
   U6823 : OAI22_X1 port map( A1 => n4334, A2 => n7112, B1 => n4366, B2 => 
                           n7109, ZN => n5237);
   U6824 : AOI221_X1 port map( B1 => n7166, B2 => n4781, C1 => n7163, C2 => 
                           n4813, A => n5210, ZN => n5205);
   U6825 : OAI22_X1 port map( A1 => n4717, A2 => n7160, B1 => n4749, B2 => 
                           n7157, ZN => n5210);
   U6826 : AOI221_X1 port map( B1 => n7118, B2 => n4397, C1 => n7115, C2 => 
                           n4429, A => n5218, ZN => n5213);
   U6827 : OAI22_X1 port map( A1 => n4333, A2 => n7112, B1 => n4365, B2 => 
                           n7109, ZN => n5218);
   U6828 : AOI221_X1 port map( B1 => n7166, B2 => n4780, C1 => n7163, C2 => 
                           n4812, A => n5191, ZN => n5186);
   U6829 : OAI22_X1 port map( A1 => n4716, A2 => n7160, B1 => n4748, B2 => 
                           n7157, ZN => n5191);
   U6830 : AOI221_X1 port map( B1 => n7118, B2 => n4396, C1 => n7115, C2 => 
                           n4428, A => n5199, ZN => n5194);
   U6831 : OAI22_X1 port map( A1 => n4332, A2 => n7112, B1 => n4364, B2 => 
                           n7109, ZN => n5199);
   U6832 : AOI221_X1 port map( B1 => n7166, B2 => n4779, C1 => n7163, C2 => 
                           n4811, A => n5172, ZN => n5167);
   U6833 : OAI22_X1 port map( A1 => n4715, A2 => n7160, B1 => n4747, B2 => 
                           n7157, ZN => n5172);
   U6834 : AOI221_X1 port map( B1 => n7118, B2 => n4395, C1 => n7115, C2 => 
                           n4427, A => n5180, ZN => n5175);
   U6835 : OAI22_X1 port map( A1 => n4331, A2 => n7112, B1 => n4363, B2 => 
                           n7109, ZN => n5180);
   U6836 : AOI221_X1 port map( B1 => n7166, B2 => n4778, C1 => n7163, C2 => 
                           n4810, A => n5131, ZN => n5116);
   U6837 : OAI22_X1 port map( A1 => n4714, A2 => n7160, B1 => n4746, B2 => 
                           n7157, ZN => n5131);
   U6838 : AOI221_X1 port map( B1 => n7118, B2 => n4394, C1 => n7115, C2 => 
                           n4426, A => n5155, ZN => n5140);
   U6839 : OAI22_X1 port map( A1 => n4330, A2 => n7112, B1 => n4362, B2 => 
                           n7109, ZN => n5155);
   U6840 : OAI22_X1 port map( A1 => n7221, A2 => n7551, B1 => n5108, B2 => 
                           n4945, ZN => n2680);
   U6841 : OAI22_X1 port map( A1 => n7222, A2 => n7554, B1 => n5108, B2 => 
                           n4944, ZN => n2681);
   U6842 : OAI22_X1 port map( A1 => n7222, A2 => n7557, B1 => n5108, B2 => 
                           n4943, ZN => n2682);
   U6843 : OAI22_X1 port map( A1 => n7222, A2 => n7560, B1 => n5108, B2 => 
                           n4942, ZN => n2683);
   U6844 : OAI22_X1 port map( A1 => n7222, A2 => n7563, B1 => n5108, B2 => 
                           n4941, ZN => n2684);
   U6845 : OAI22_X1 port map( A1 => n7222, A2 => n7566, B1 => n5108, B2 => 
                           n4940, ZN => n2685);
   U6846 : OAI22_X1 port map( A1 => n7223, A2 => n7569, B1 => n5108, B2 => 
                           n4939, ZN => n2686);
   U6847 : OAI22_X1 port map( A1 => n7223, A2 => n7581, B1 => n5108, B2 => 
                           n4938, ZN => n2687);
   U6848 : OAI22_X1 port map( A1 => n7230, A2 => n7551, B1 => n5107, B2 => 
                           n4913, ZN => n2712);
   U6849 : OAI22_X1 port map( A1 => n7231, A2 => n7554, B1 => n5107, B2 => 
                           n4912, ZN => n2713);
   U6850 : OAI22_X1 port map( A1 => n7231, A2 => n7557, B1 => n5107, B2 => 
                           n4911, ZN => n2714);
   U6851 : OAI22_X1 port map( A1 => n7231, A2 => n7560, B1 => n5107, B2 => 
                           n4910, ZN => n2715);
   U6852 : OAI22_X1 port map( A1 => n7231, A2 => n7563, B1 => n5107, B2 => 
                           n4909, ZN => n2716);
   U6853 : OAI22_X1 port map( A1 => n7231, A2 => n7566, B1 => n5107, B2 => 
                           n4908, ZN => n2717);
   U6854 : OAI22_X1 port map( A1 => n7232, A2 => n7569, B1 => n5107, B2 => 
                           n4907, ZN => n2718);
   U6855 : OAI22_X1 port map( A1 => n7232, A2 => n7581, B1 => n5107, B2 => 
                           n4906, ZN => n2719);
   U6856 : OAI22_X1 port map( A1 => n7293, A2 => n7550, B1 => n5099, B2 => 
                           n4753, ZN => n2936);
   U6857 : OAI22_X1 port map( A1 => n7294, A2 => n7553, B1 => n5099, B2 => 
                           n4752, ZN => n2937);
   U6858 : OAI22_X1 port map( A1 => n7294, A2 => n7556, B1 => n5099, B2 => 
                           n4751, ZN => n2938);
   U6859 : OAI22_X1 port map( A1 => n7294, A2 => n7559, B1 => n5099, B2 => 
                           n4750, ZN => n2939);
   U6860 : OAI22_X1 port map( A1 => n7294, A2 => n7562, B1 => n5099, B2 => 
                           n4749, ZN => n2940);
   U6861 : OAI22_X1 port map( A1 => n7294, A2 => n7565, B1 => n5099, B2 => 
                           n4748, ZN => n2941);
   U6862 : OAI22_X1 port map( A1 => n7295, A2 => n7568, B1 => n5099, B2 => 
                           n4747, ZN => n2942);
   U6863 : OAI22_X1 port map( A1 => n7295, A2 => n7580, B1 => n5099, B2 => 
                           n4746, ZN => n2943);
   U6864 : OAI22_X1 port map( A1 => n7302, A2 => n7550, B1 => n5098, B2 => 
                           n4721, ZN => n2968);
   U6865 : OAI22_X1 port map( A1 => n7303, A2 => n7553, B1 => n5098, B2 => 
                           n4720, ZN => n2969);
   U6866 : OAI22_X1 port map( A1 => n7303, A2 => n7556, B1 => n5098, B2 => 
                           n4719, ZN => n2970);
   U6867 : OAI22_X1 port map( A1 => n7303, A2 => n7559, B1 => n5098, B2 => 
                           n4718, ZN => n2971);
   U6868 : OAI22_X1 port map( A1 => n7303, A2 => n7562, B1 => n5098, B2 => 
                           n4717, ZN => n2972);
   U6869 : OAI22_X1 port map( A1 => n7303, A2 => n7565, B1 => n5098, B2 => 
                           n4716, ZN => n2973);
   U6870 : OAI22_X1 port map( A1 => n7304, A2 => n7568, B1 => n5098, B2 => 
                           n4715, ZN => n2974);
   U6871 : OAI22_X1 port map( A1 => n7304, A2 => n7580, B1 => n5098, B2 => 
                           n4714, ZN => n2975);
   U6872 : OAI22_X1 port map( A1 => n7365, A2 => n7550, B1 => n5090, B2 => 
                           n4561, ZN => n3192);
   U6873 : OAI22_X1 port map( A1 => n7366, A2 => n7553, B1 => n5090, B2 => 
                           n4560, ZN => n3193);
   U6874 : OAI22_X1 port map( A1 => n7366, A2 => n7556, B1 => n5090, B2 => 
                           n4559, ZN => n3194);
   U6875 : OAI22_X1 port map( A1 => n7366, A2 => n7559, B1 => n5090, B2 => 
                           n4558, ZN => n3195);
   U6876 : OAI22_X1 port map( A1 => n7366, A2 => n7562, B1 => n5090, B2 => 
                           n4557, ZN => n3196);
   U6877 : OAI22_X1 port map( A1 => n7366, A2 => n7565, B1 => n5090, B2 => 
                           n4556, ZN => n3197);
   U6878 : OAI22_X1 port map( A1 => n7367, A2 => n7568, B1 => n5090, B2 => 
                           n4555, ZN => n3198);
   U6879 : OAI22_X1 port map( A1 => n7367, A2 => n7580, B1 => n5090, B2 => 
                           n4554, ZN => n3199);
   U6880 : OAI22_X1 port map( A1 => n7374, A2 => n7550, B1 => n5089, B2 => 
                           n4529, ZN => n3224);
   U6881 : OAI22_X1 port map( A1 => n7375, A2 => n7553, B1 => n5089, B2 => 
                           n4528, ZN => n3225);
   U6882 : OAI22_X1 port map( A1 => n7375, A2 => n7556, B1 => n5089, B2 => 
                           n4527, ZN => n3226);
   U6883 : OAI22_X1 port map( A1 => n7375, A2 => n7559, B1 => n5089, B2 => 
                           n4526, ZN => n3227);
   U6884 : OAI22_X1 port map( A1 => n7375, A2 => n7562, B1 => n5089, B2 => 
                           n4525, ZN => n3228);
   U6885 : OAI22_X1 port map( A1 => n7375, A2 => n7565, B1 => n5089, B2 => 
                           n4524, ZN => n3229);
   U6886 : OAI22_X1 port map( A1 => n7376, A2 => n7568, B1 => n5089, B2 => 
                           n4523, ZN => n3230);
   U6887 : OAI22_X1 port map( A1 => n7376, A2 => n7580, B1 => n5089, B2 => 
                           n4522, ZN => n3231);
   U6888 : OAI22_X1 port map( A1 => n7437, A2 => n7549, B1 => n5077, B2 => 
                           n4369, ZN => n3448);
   U6889 : OAI22_X1 port map( A1 => n7438, A2 => n7552, B1 => n5077, B2 => 
                           n4368, ZN => n3449);
   U6890 : OAI22_X1 port map( A1 => n7438, A2 => n7555, B1 => n5077, B2 => 
                           n4367, ZN => n3450);
   U6891 : OAI22_X1 port map( A1 => n7438, A2 => n7558, B1 => n5077, B2 => 
                           n4366, ZN => n3451);
   U6892 : OAI22_X1 port map( A1 => n7438, A2 => n7561, B1 => n5077, B2 => 
                           n4365, ZN => n3452);
   U6893 : OAI22_X1 port map( A1 => n7438, A2 => n7564, B1 => n5077, B2 => 
                           n4364, ZN => n3453);
   U6894 : OAI22_X1 port map( A1 => n7439, A2 => n7567, B1 => n5077, B2 => 
                           n4363, ZN => n3454);
   U6895 : OAI22_X1 port map( A1 => n7439, A2 => n7579, B1 => n5077, B2 => 
                           n4362, ZN => n3455);
   U6896 : OAI22_X1 port map( A1 => n7446, A2 => n7549, B1 => n5075, B2 => 
                           n4337, ZN => n3480);
   U6897 : OAI22_X1 port map( A1 => n7447, A2 => n7552, B1 => n5075, B2 => 
                           n4336, ZN => n3481);
   U6898 : OAI22_X1 port map( A1 => n7447, A2 => n7555, B1 => n5075, B2 => 
                           n4335, ZN => n3482);
   U6899 : OAI22_X1 port map( A1 => n7447, A2 => n7558, B1 => n5075, B2 => 
                           n4334, ZN => n3483);
   U6900 : OAI22_X1 port map( A1 => n7447, A2 => n7561, B1 => n5075, B2 => 
                           n4333, ZN => n3484);
   U6901 : OAI22_X1 port map( A1 => n7447, A2 => n7564, B1 => n5075, B2 => 
                           n4332, ZN => n3485);
   U6902 : OAI22_X1 port map( A1 => n7448, A2 => n7567, B1 => n5075, B2 => 
                           n4331, ZN => n3486);
   U6903 : OAI22_X1 port map( A1 => n7448, A2 => n7579, B1 => n5075, B2 => 
                           n4330, ZN => n3487);
   U6904 : OAI22_X1 port map( A1 => n7217, A2 => n7479, B1 => n7216, B2 => 
                           n4969, ZN => n2656);
   U6905 : OAI22_X1 port map( A1 => n7217, A2 => n7482, B1 => n7216, B2 => 
                           n4968, ZN => n2657);
   U6906 : OAI22_X1 port map( A1 => n7217, A2 => n7485, B1 => n7216, B2 => 
                           n4967, ZN => n2658);
   U6907 : OAI22_X1 port map( A1 => n7217, A2 => n7488, B1 => n7216, B2 => 
                           n4966, ZN => n2659);
   U6908 : OAI22_X1 port map( A1 => n7217, A2 => n7491, B1 => n7216, B2 => 
                           n4965, ZN => n2660);
   U6909 : OAI22_X1 port map( A1 => n7218, A2 => n7494, B1 => n7216, B2 => 
                           n4964, ZN => n2661);
   U6910 : OAI22_X1 port map( A1 => n7218, A2 => n7497, B1 => n7216, B2 => 
                           n4963, ZN => n2662);
   U6911 : OAI22_X1 port map( A1 => n7218, A2 => n7500, B1 => n7216, B2 => 
                           n4962, ZN => n2663);
   U6912 : OAI22_X1 port map( A1 => n7218, A2 => n7503, B1 => n7216, B2 => 
                           n4961, ZN => n2664);
   U6913 : OAI22_X1 port map( A1 => n7218, A2 => n7506, B1 => n7216, B2 => 
                           n4960, ZN => n2665);
   U6914 : OAI22_X1 port map( A1 => n7219, A2 => n7509, B1 => n7216, B2 => 
                           n4959, ZN => n2666);
   U6915 : OAI22_X1 port map( A1 => n7219, A2 => n7512, B1 => n7216, B2 => 
                           n4958, ZN => n2667);
   U6916 : OAI22_X1 port map( A1 => n7219, A2 => n7515, B1 => n5108, B2 => 
                           n4957, ZN => n2668);
   U6917 : OAI22_X1 port map( A1 => n7219, A2 => n7518, B1 => n5108, B2 => 
                           n4956, ZN => n2669);
   U6918 : OAI22_X1 port map( A1 => n7219, A2 => n7521, B1 => n5108, B2 => 
                           n4955, ZN => n2670);
   U6919 : OAI22_X1 port map( A1 => n7220, A2 => n7524, B1 => n7216, B2 => 
                           n4954, ZN => n2671);
   U6920 : OAI22_X1 port map( A1 => n7220, A2 => n7527, B1 => n7216, B2 => 
                           n4953, ZN => n2672);
   U6921 : OAI22_X1 port map( A1 => n7220, A2 => n7530, B1 => n7216, B2 => 
                           n4952, ZN => n2673);
   U6922 : OAI22_X1 port map( A1 => n7220, A2 => n7533, B1 => n7216, B2 => 
                           n4951, ZN => n2674);
   U6923 : OAI22_X1 port map( A1 => n7220, A2 => n7536, B1 => n7216, B2 => 
                           n4950, ZN => n2675);
   U6924 : OAI22_X1 port map( A1 => n7221, A2 => n7539, B1 => n7216, B2 => 
                           n4949, ZN => n2676);
   U6925 : OAI22_X1 port map( A1 => n7221, A2 => n7542, B1 => n7216, B2 => 
                           n4948, ZN => n2677);
   U6926 : OAI22_X1 port map( A1 => n7221, A2 => n7545, B1 => n7216, B2 => 
                           n4947, ZN => n2678);
   U6927 : OAI22_X1 port map( A1 => n7221, A2 => n7548, B1 => n7216, B2 => 
                           n4946, ZN => n2679);
   U6928 : OAI22_X1 port map( A1 => n7226, A2 => n7479, B1 => n7225, B2 => 
                           n4937, ZN => n2688);
   U6929 : OAI22_X1 port map( A1 => n7226, A2 => n7482, B1 => n7225, B2 => 
                           n4936, ZN => n2689);
   U6930 : OAI22_X1 port map( A1 => n7226, A2 => n7485, B1 => n7225, B2 => 
                           n4935, ZN => n2690);
   U6931 : OAI22_X1 port map( A1 => n7226, A2 => n7488, B1 => n7225, B2 => 
                           n4934, ZN => n2691);
   U6932 : OAI22_X1 port map( A1 => n7226, A2 => n7491, B1 => n7225, B2 => 
                           n4933, ZN => n2692);
   U6933 : OAI22_X1 port map( A1 => n7227, A2 => n7494, B1 => n7225, B2 => 
                           n4932, ZN => n2693);
   U6934 : OAI22_X1 port map( A1 => n7227, A2 => n7497, B1 => n7225, B2 => 
                           n4931, ZN => n2694);
   U6935 : OAI22_X1 port map( A1 => n7227, A2 => n7500, B1 => n7225, B2 => 
                           n4930, ZN => n2695);
   U6936 : OAI22_X1 port map( A1 => n7227, A2 => n7503, B1 => n7225, B2 => 
                           n4929, ZN => n2696);
   U6937 : OAI22_X1 port map( A1 => n7227, A2 => n7506, B1 => n7225, B2 => 
                           n4928, ZN => n2697);
   U6938 : OAI22_X1 port map( A1 => n7228, A2 => n7509, B1 => n7225, B2 => 
                           n4927, ZN => n2698);
   U6939 : OAI22_X1 port map( A1 => n7228, A2 => n7512, B1 => n7225, B2 => 
                           n4926, ZN => n2699);
   U6940 : OAI22_X1 port map( A1 => n7228, A2 => n7515, B1 => n5107, B2 => 
                           n4925, ZN => n2700);
   U6941 : OAI22_X1 port map( A1 => n7228, A2 => n7518, B1 => n5107, B2 => 
                           n4924, ZN => n2701);
   U6942 : OAI22_X1 port map( A1 => n7228, A2 => n7521, B1 => n5107, B2 => 
                           n4923, ZN => n2702);
   U6943 : OAI22_X1 port map( A1 => n7229, A2 => n7524, B1 => n7225, B2 => 
                           n4922, ZN => n2703);
   U6944 : OAI22_X1 port map( A1 => n7229, A2 => n7527, B1 => n7225, B2 => 
                           n4921, ZN => n2704);
   U6945 : OAI22_X1 port map( A1 => n7229, A2 => n7530, B1 => n7225, B2 => 
                           n4920, ZN => n2705);
   U6946 : OAI22_X1 port map( A1 => n7229, A2 => n7533, B1 => n7225, B2 => 
                           n4919, ZN => n2706);
   U6947 : OAI22_X1 port map( A1 => n7229, A2 => n7536, B1 => n7225, B2 => 
                           n4918, ZN => n2707);
   U6948 : OAI22_X1 port map( A1 => n7230, A2 => n7539, B1 => n7225, B2 => 
                           n4917, ZN => n2708);
   U6949 : OAI22_X1 port map( A1 => n7230, A2 => n7542, B1 => n7225, B2 => 
                           n4916, ZN => n2709);
   U6950 : OAI22_X1 port map( A1 => n7230, A2 => n7545, B1 => n7225, B2 => 
                           n4915, ZN => n2710);
   U6951 : OAI22_X1 port map( A1 => n7230, A2 => n7548, B1 => n7225, B2 => 
                           n4914, ZN => n2711);
   U6952 : OAI22_X1 port map( A1 => n7289, A2 => n7478, B1 => n7288, B2 => 
                           n4777, ZN => n2912);
   U6953 : OAI22_X1 port map( A1 => n7289, A2 => n7481, B1 => n7288, B2 => 
                           n4776, ZN => n2913);
   U6954 : OAI22_X1 port map( A1 => n7289, A2 => n7484, B1 => n7288, B2 => 
                           n4775, ZN => n2914);
   U6955 : OAI22_X1 port map( A1 => n7289, A2 => n7487, B1 => n7288, B2 => 
                           n4774, ZN => n2915);
   U6956 : OAI22_X1 port map( A1 => n7289, A2 => n7490, B1 => n7288, B2 => 
                           n4773, ZN => n2916);
   U6957 : OAI22_X1 port map( A1 => n7290, A2 => n7493, B1 => n7288, B2 => 
                           n4772, ZN => n2917);
   U6958 : OAI22_X1 port map( A1 => n7290, A2 => n7496, B1 => n7288, B2 => 
                           n4771, ZN => n2918);
   U6959 : OAI22_X1 port map( A1 => n7290, A2 => n7499, B1 => n7288, B2 => 
                           n4770, ZN => n2919);
   U6960 : OAI22_X1 port map( A1 => n7290, A2 => n7502, B1 => n7288, B2 => 
                           n4769, ZN => n2920);
   U6961 : OAI22_X1 port map( A1 => n7290, A2 => n7505, B1 => n7288, B2 => 
                           n4768, ZN => n2921);
   U6962 : OAI22_X1 port map( A1 => n7291, A2 => n7508, B1 => n7288, B2 => 
                           n4767, ZN => n2922);
   U6963 : OAI22_X1 port map( A1 => n7291, A2 => n7511, B1 => n7288, B2 => 
                           n4766, ZN => n2923);
   U6964 : OAI22_X1 port map( A1 => n7291, A2 => n7514, B1 => n5099, B2 => 
                           n4765, ZN => n2924);
   U6965 : OAI22_X1 port map( A1 => n7291, A2 => n7517, B1 => n5099, B2 => 
                           n4764, ZN => n2925);
   U6966 : OAI22_X1 port map( A1 => n7291, A2 => n7520, B1 => n5099, B2 => 
                           n4763, ZN => n2926);
   U6967 : OAI22_X1 port map( A1 => n7292, A2 => n7523, B1 => n7288, B2 => 
                           n4762, ZN => n2927);
   U6968 : OAI22_X1 port map( A1 => n7292, A2 => n7526, B1 => n7288, B2 => 
                           n4761, ZN => n2928);
   U6969 : OAI22_X1 port map( A1 => n7292, A2 => n7529, B1 => n7288, B2 => 
                           n4760, ZN => n2929);
   U6970 : OAI22_X1 port map( A1 => n7292, A2 => n7532, B1 => n7288, B2 => 
                           n4759, ZN => n2930);
   U6971 : OAI22_X1 port map( A1 => n7292, A2 => n7535, B1 => n7288, B2 => 
                           n4758, ZN => n2931);
   U6972 : OAI22_X1 port map( A1 => n7293, A2 => n7538, B1 => n7288, B2 => 
                           n4757, ZN => n2932);
   U6973 : OAI22_X1 port map( A1 => n7293, A2 => n7541, B1 => n7288, B2 => 
                           n4756, ZN => n2933);
   U6974 : OAI22_X1 port map( A1 => n7293, A2 => n7544, B1 => n7288, B2 => 
                           n4755, ZN => n2934);
   U6975 : OAI22_X1 port map( A1 => n7293, A2 => n7547, B1 => n7288, B2 => 
                           n4754, ZN => n2935);
   U6976 : OAI22_X1 port map( A1 => n7298, A2 => n7478, B1 => n7297, B2 => 
                           n4745, ZN => n2944);
   U6977 : OAI22_X1 port map( A1 => n7298, A2 => n7481, B1 => n7297, B2 => 
                           n4744, ZN => n2945);
   U6978 : OAI22_X1 port map( A1 => n7298, A2 => n7484, B1 => n7297, B2 => 
                           n4743, ZN => n2946);
   U6979 : OAI22_X1 port map( A1 => n7298, A2 => n7487, B1 => n7297, B2 => 
                           n4742, ZN => n2947);
   U6980 : OAI22_X1 port map( A1 => n7298, A2 => n7490, B1 => n7297, B2 => 
                           n4741, ZN => n2948);
   U6981 : OAI22_X1 port map( A1 => n7299, A2 => n7493, B1 => n7297, B2 => 
                           n4740, ZN => n2949);
   U6982 : OAI22_X1 port map( A1 => n7299, A2 => n7496, B1 => n7297, B2 => 
                           n4739, ZN => n2950);
   U6983 : OAI22_X1 port map( A1 => n7299, A2 => n7499, B1 => n7297, B2 => 
                           n4738, ZN => n2951);
   U6984 : OAI22_X1 port map( A1 => n7299, A2 => n7502, B1 => n7297, B2 => 
                           n4737, ZN => n2952);
   U6985 : OAI22_X1 port map( A1 => n7299, A2 => n7505, B1 => n7297, B2 => 
                           n4736, ZN => n2953);
   U6986 : OAI22_X1 port map( A1 => n7300, A2 => n7508, B1 => n7297, B2 => 
                           n4735, ZN => n2954);
   U6987 : OAI22_X1 port map( A1 => n7300, A2 => n7511, B1 => n7297, B2 => 
                           n4734, ZN => n2955);
   U6988 : OAI22_X1 port map( A1 => n7300, A2 => n7514, B1 => n5098, B2 => 
                           n4733, ZN => n2956);
   U6989 : OAI22_X1 port map( A1 => n7300, A2 => n7517, B1 => n5098, B2 => 
                           n4732, ZN => n2957);
   U6990 : OAI22_X1 port map( A1 => n7300, A2 => n7520, B1 => n5098, B2 => 
                           n4731, ZN => n2958);
   U6991 : OAI22_X1 port map( A1 => n7301, A2 => n7523, B1 => n7297, B2 => 
                           n4730, ZN => n2959);
   U6992 : OAI22_X1 port map( A1 => n7301, A2 => n7526, B1 => n7297, B2 => 
                           n4729, ZN => n2960);
   U6993 : OAI22_X1 port map( A1 => n7301, A2 => n7529, B1 => n7297, B2 => 
                           n4728, ZN => n2961);
   U6994 : OAI22_X1 port map( A1 => n7301, A2 => n7532, B1 => n7297, B2 => 
                           n4727, ZN => n2962);
   U6995 : OAI22_X1 port map( A1 => n7301, A2 => n7535, B1 => n7297, B2 => 
                           n4726, ZN => n2963);
   U6996 : OAI22_X1 port map( A1 => n7302, A2 => n7538, B1 => n7297, B2 => 
                           n4725, ZN => n2964);
   U6997 : OAI22_X1 port map( A1 => n7302, A2 => n7541, B1 => n7297, B2 => 
                           n4724, ZN => n2965);
   U6998 : OAI22_X1 port map( A1 => n7302, A2 => n7544, B1 => n7297, B2 => 
                           n4723, ZN => n2966);
   U6999 : OAI22_X1 port map( A1 => n7302, A2 => n7547, B1 => n7297, B2 => 
                           n4722, ZN => n2967);
   U7000 : OAI22_X1 port map( A1 => n7361, A2 => n7478, B1 => n7360, B2 => 
                           n4585, ZN => n3168);
   U7001 : OAI22_X1 port map( A1 => n7361, A2 => n7481, B1 => n7360, B2 => 
                           n4584, ZN => n3169);
   U7002 : OAI22_X1 port map( A1 => n7361, A2 => n7484, B1 => n7360, B2 => 
                           n4583, ZN => n3170);
   U7003 : OAI22_X1 port map( A1 => n7361, A2 => n7487, B1 => n7360, B2 => 
                           n4582, ZN => n3171);
   U7004 : OAI22_X1 port map( A1 => n7361, A2 => n7490, B1 => n7360, B2 => 
                           n4581, ZN => n3172);
   U7005 : OAI22_X1 port map( A1 => n7362, A2 => n7493, B1 => n7360, B2 => 
                           n4580, ZN => n3173);
   U7006 : OAI22_X1 port map( A1 => n7362, A2 => n7496, B1 => n7360, B2 => 
                           n4579, ZN => n3174);
   U7007 : OAI22_X1 port map( A1 => n7362, A2 => n7499, B1 => n7360, B2 => 
                           n4578, ZN => n3175);
   U7008 : OAI22_X1 port map( A1 => n7362, A2 => n7502, B1 => n7360, B2 => 
                           n4577, ZN => n3176);
   U7009 : OAI22_X1 port map( A1 => n7362, A2 => n7505, B1 => n7360, B2 => 
                           n4576, ZN => n3177);
   U7010 : OAI22_X1 port map( A1 => n7363, A2 => n7508, B1 => n7360, B2 => 
                           n4575, ZN => n3178);
   U7011 : OAI22_X1 port map( A1 => n7363, A2 => n7511, B1 => n7360, B2 => 
                           n4574, ZN => n3179);
   U7012 : OAI22_X1 port map( A1 => n7363, A2 => n7514, B1 => n5090, B2 => 
                           n4573, ZN => n3180);
   U7013 : OAI22_X1 port map( A1 => n7363, A2 => n7517, B1 => n5090, B2 => 
                           n4572, ZN => n3181);
   U7014 : OAI22_X1 port map( A1 => n7363, A2 => n7520, B1 => n5090, B2 => 
                           n4571, ZN => n3182);
   U7015 : OAI22_X1 port map( A1 => n7364, A2 => n7523, B1 => n7360, B2 => 
                           n4570, ZN => n3183);
   U7016 : OAI22_X1 port map( A1 => n7364, A2 => n7526, B1 => n7360, B2 => 
                           n4569, ZN => n3184);
   U7017 : OAI22_X1 port map( A1 => n7364, A2 => n7529, B1 => n7360, B2 => 
                           n4568, ZN => n3185);
   U7018 : OAI22_X1 port map( A1 => n7364, A2 => n7532, B1 => n7360, B2 => 
                           n4567, ZN => n3186);
   U7019 : OAI22_X1 port map( A1 => n7364, A2 => n7535, B1 => n7360, B2 => 
                           n4566, ZN => n3187);
   U7020 : OAI22_X1 port map( A1 => n7365, A2 => n7538, B1 => n7360, B2 => 
                           n4565, ZN => n3188);
   U7021 : OAI22_X1 port map( A1 => n7365, A2 => n7541, B1 => n7360, B2 => 
                           n4564, ZN => n3189);
   U7022 : OAI22_X1 port map( A1 => n7365, A2 => n7544, B1 => n7360, B2 => 
                           n4563, ZN => n3190);
   U7023 : OAI22_X1 port map( A1 => n7365, A2 => n7547, B1 => n7360, B2 => 
                           n4562, ZN => n3191);
   U7024 : OAI22_X1 port map( A1 => n7370, A2 => n7478, B1 => n7369, B2 => 
                           n4553, ZN => n3200);
   U7025 : OAI22_X1 port map( A1 => n7370, A2 => n7481, B1 => n7369, B2 => 
                           n4552, ZN => n3201);
   U7026 : OAI22_X1 port map( A1 => n7370, A2 => n7484, B1 => n7369, B2 => 
                           n4551, ZN => n3202);
   U7027 : OAI22_X1 port map( A1 => n7370, A2 => n7487, B1 => n7369, B2 => 
                           n4550, ZN => n3203);
   U7028 : OAI22_X1 port map( A1 => n7370, A2 => n7490, B1 => n7369, B2 => 
                           n4549, ZN => n3204);
   U7029 : OAI22_X1 port map( A1 => n7371, A2 => n7493, B1 => n7369, B2 => 
                           n4548, ZN => n3205);
   U7030 : OAI22_X1 port map( A1 => n7371, A2 => n7496, B1 => n7369, B2 => 
                           n4547, ZN => n3206);
   U7031 : OAI22_X1 port map( A1 => n7371, A2 => n7499, B1 => n7369, B2 => 
                           n4546, ZN => n3207);
   U7032 : OAI22_X1 port map( A1 => n7371, A2 => n7502, B1 => n7369, B2 => 
                           n4545, ZN => n3208);
   U7033 : OAI22_X1 port map( A1 => n7371, A2 => n7505, B1 => n7369, B2 => 
                           n4544, ZN => n3209);
   U7034 : OAI22_X1 port map( A1 => n7372, A2 => n7508, B1 => n7369, B2 => 
                           n4543, ZN => n3210);
   U7035 : OAI22_X1 port map( A1 => n7372, A2 => n7511, B1 => n7369, B2 => 
                           n4542, ZN => n3211);
   U7036 : OAI22_X1 port map( A1 => n7372, A2 => n7514, B1 => n5089, B2 => 
                           n4541, ZN => n3212);
   U7037 : OAI22_X1 port map( A1 => n7372, A2 => n7517, B1 => n5089, B2 => 
                           n4540, ZN => n3213);
   U7038 : OAI22_X1 port map( A1 => n7372, A2 => n7520, B1 => n5089, B2 => 
                           n4539, ZN => n3214);
   U7039 : OAI22_X1 port map( A1 => n7373, A2 => n7523, B1 => n7369, B2 => 
                           n4538, ZN => n3215);
   U7040 : OAI22_X1 port map( A1 => n7373, A2 => n7526, B1 => n7369, B2 => 
                           n4537, ZN => n3216);
   U7041 : OAI22_X1 port map( A1 => n7373, A2 => n7529, B1 => n7369, B2 => 
                           n4536, ZN => n3217);
   U7042 : OAI22_X1 port map( A1 => n7373, A2 => n7532, B1 => n7369, B2 => 
                           n4535, ZN => n3218);
   U7043 : OAI22_X1 port map( A1 => n7373, A2 => n7535, B1 => n7369, B2 => 
                           n4534, ZN => n3219);
   U7044 : OAI22_X1 port map( A1 => n7374, A2 => n7538, B1 => n7369, B2 => 
                           n4533, ZN => n3220);
   U7045 : OAI22_X1 port map( A1 => n7374, A2 => n7541, B1 => n7369, B2 => 
                           n4532, ZN => n3221);
   U7046 : OAI22_X1 port map( A1 => n7374, A2 => n7544, B1 => n7369, B2 => 
                           n4531, ZN => n3222);
   U7047 : OAI22_X1 port map( A1 => n7374, A2 => n7547, B1 => n7369, B2 => 
                           n4530, ZN => n3223);
   U7048 : OAI22_X1 port map( A1 => n7433, A2 => n7477, B1 => n7432, B2 => 
                           n4393, ZN => n3424);
   U7049 : OAI22_X1 port map( A1 => n7433, A2 => n7480, B1 => n7432, B2 => 
                           n4392, ZN => n3425);
   U7050 : OAI22_X1 port map( A1 => n7433, A2 => n7483, B1 => n7432, B2 => 
                           n4391, ZN => n3426);
   U7051 : OAI22_X1 port map( A1 => n7433, A2 => n7486, B1 => n7432, B2 => 
                           n4390, ZN => n3427);
   U7052 : OAI22_X1 port map( A1 => n7433, A2 => n7489, B1 => n7432, B2 => 
                           n4389, ZN => n3428);
   U7053 : OAI22_X1 port map( A1 => n7434, A2 => n7492, B1 => n7432, B2 => 
                           n4388, ZN => n3429);
   U7054 : OAI22_X1 port map( A1 => n7434, A2 => n7495, B1 => n7432, B2 => 
                           n4387, ZN => n3430);
   U7055 : OAI22_X1 port map( A1 => n7434, A2 => n7498, B1 => n7432, B2 => 
                           n4386, ZN => n3431);
   U7056 : OAI22_X1 port map( A1 => n7434, A2 => n7501, B1 => n7432, B2 => 
                           n4385, ZN => n3432);
   U7057 : OAI22_X1 port map( A1 => n7434, A2 => n7504, B1 => n7432, B2 => 
                           n4384, ZN => n3433);
   U7058 : OAI22_X1 port map( A1 => n7435, A2 => n7507, B1 => n7432, B2 => 
                           n4383, ZN => n3434);
   U7059 : OAI22_X1 port map( A1 => n7435, A2 => n7510, B1 => n7432, B2 => 
                           n4382, ZN => n3435);
   U7060 : OAI22_X1 port map( A1 => n7435, A2 => n7513, B1 => n5077, B2 => 
                           n4381, ZN => n3436);
   U7061 : OAI22_X1 port map( A1 => n7435, A2 => n7516, B1 => n5077, B2 => 
                           n4380, ZN => n3437);
   U7062 : OAI22_X1 port map( A1 => n7435, A2 => n7519, B1 => n5077, B2 => 
                           n4379, ZN => n3438);
   U7063 : OAI22_X1 port map( A1 => n7436, A2 => n7522, B1 => n7432, B2 => 
                           n4378, ZN => n3439);
   U7064 : OAI22_X1 port map( A1 => n7436, A2 => n7525, B1 => n7432, B2 => 
                           n4377, ZN => n3440);
   U7065 : OAI22_X1 port map( A1 => n7436, A2 => n7528, B1 => n7432, B2 => 
                           n4376, ZN => n3441);
   U7066 : OAI22_X1 port map( A1 => n7436, A2 => n7531, B1 => n7432, B2 => 
                           n4375, ZN => n3442);
   U7067 : OAI22_X1 port map( A1 => n7436, A2 => n7534, B1 => n7432, B2 => 
                           n4374, ZN => n3443);
   U7068 : OAI22_X1 port map( A1 => n7437, A2 => n7537, B1 => n7432, B2 => 
                           n4373, ZN => n3444);
   U7069 : OAI22_X1 port map( A1 => n7437, A2 => n7540, B1 => n7432, B2 => 
                           n4372, ZN => n3445);
   U7070 : OAI22_X1 port map( A1 => n7437, A2 => n7543, B1 => n7432, B2 => 
                           n4371, ZN => n3446);
   U7071 : OAI22_X1 port map( A1 => n7437, A2 => n7546, B1 => n7432, B2 => 
                           n4370, ZN => n3447);
   U7072 : OAI22_X1 port map( A1 => n7442, A2 => n7477, B1 => n7441, B2 => 
                           n4361, ZN => n3456);
   U7073 : OAI22_X1 port map( A1 => n7442, A2 => n7480, B1 => n7441, B2 => 
                           n4360, ZN => n3457);
   U7074 : OAI22_X1 port map( A1 => n7442, A2 => n7483, B1 => n7441, B2 => 
                           n4359, ZN => n3458);
   U7075 : OAI22_X1 port map( A1 => n7442, A2 => n7486, B1 => n7441, B2 => 
                           n4358, ZN => n3459);
   U7076 : OAI22_X1 port map( A1 => n7442, A2 => n7489, B1 => n7441, B2 => 
                           n4357, ZN => n3460);
   U7077 : OAI22_X1 port map( A1 => n7443, A2 => n7492, B1 => n7441, B2 => 
                           n4356, ZN => n3461);
   U7078 : OAI22_X1 port map( A1 => n7443, A2 => n7495, B1 => n7441, B2 => 
                           n4355, ZN => n3462);
   U7079 : OAI22_X1 port map( A1 => n7443, A2 => n7498, B1 => n7441, B2 => 
                           n4354, ZN => n3463);
   U7080 : OAI22_X1 port map( A1 => n7443, A2 => n7501, B1 => n7441, B2 => 
                           n4353, ZN => n3464);
   U7081 : OAI22_X1 port map( A1 => n7443, A2 => n7504, B1 => n7441, B2 => 
                           n4352, ZN => n3465);
   U7082 : OAI22_X1 port map( A1 => n7444, A2 => n7507, B1 => n7441, B2 => 
                           n4351, ZN => n3466);
   U7083 : OAI22_X1 port map( A1 => n7444, A2 => n7510, B1 => n7441, B2 => 
                           n4350, ZN => n3467);
   U7084 : OAI22_X1 port map( A1 => n7444, A2 => n7513, B1 => n5075, B2 => 
                           n4349, ZN => n3468);
   U7085 : OAI22_X1 port map( A1 => n7444, A2 => n7516, B1 => n5075, B2 => 
                           n4348, ZN => n3469);
   U7086 : OAI22_X1 port map( A1 => n7444, A2 => n7519, B1 => n5075, B2 => 
                           n4347, ZN => n3470);
   U7087 : OAI22_X1 port map( A1 => n7445, A2 => n7522, B1 => n7441, B2 => 
                           n4346, ZN => n3471);
   U7088 : OAI22_X1 port map( A1 => n7445, A2 => n7525, B1 => n7441, B2 => 
                           n4345, ZN => n3472);
   U7089 : OAI22_X1 port map( A1 => n7445, A2 => n7528, B1 => n7441, B2 => 
                           n4344, ZN => n3473);
   U7090 : OAI22_X1 port map( A1 => n7445, A2 => n7531, B1 => n7441, B2 => 
                           n4343, ZN => n3474);
   U7091 : OAI22_X1 port map( A1 => n7445, A2 => n7534, B1 => n7441, B2 => 
                           n4342, ZN => n3475);
   U7092 : OAI22_X1 port map( A1 => n7446, A2 => n7537, B1 => n7441, B2 => 
                           n4341, ZN => n3476);
   U7093 : OAI22_X1 port map( A1 => n7446, A2 => n7540, B1 => n7441, B2 => 
                           n4340, ZN => n3477);
   U7094 : OAI22_X1 port map( A1 => n7446, A2 => n7543, B1 => n7441, B2 => 
                           n4339, ZN => n3478);
   U7095 : OAI22_X1 port map( A1 => n7446, A2 => n7546, B1 => n7441, B2 => 
                           n4338, ZN => n3479);
   U7096 : BUF_X1 port map( A => n5764, Z => n7090);
   U7097 : BUF_X1 port map( A => n5111, Z => n7192);
   U7098 : BUF_X1 port map( A => n5764, Z => n7091);
   U7099 : BUF_X1 port map( A => n5111, Z => n7193);
   U7100 : BUF_X1 port map( A => n5764, Z => n7092);
   U7101 : BUF_X1 port map( A => n5764, Z => n7093);
   U7102 : BUF_X1 port map( A => n5111, Z => n7194);
   U7103 : BUF_X1 port map( A => n5111, Z => n7195);
   U7104 : BUF_X1 port map( A => n4254, Z => n7585);
   U7105 : BUF_X1 port map( A => n4254, Z => n7586);
   U7106 : BUF_X1 port map( A => n4254, Z => n7583);
   U7107 : BUF_X1 port map( A => n4254, Z => n7582);
   U7108 : BUF_X1 port map( A => n5066, Z => n7478);
   U7109 : BUF_X1 port map( A => n5065, Z => n7481);
   U7110 : BUF_X1 port map( A => n5064, Z => n7484);
   U7111 : BUF_X1 port map( A => n5063, Z => n7487);
   U7112 : BUF_X1 port map( A => n5062, Z => n7490);
   U7113 : BUF_X1 port map( A => n5061, Z => n7493);
   U7114 : BUF_X1 port map( A => n5060, Z => n7496);
   U7115 : BUF_X1 port map( A => n5059, Z => n7499);
   U7116 : BUF_X1 port map( A => n5058, Z => n7502);
   U7117 : BUF_X1 port map( A => n5057, Z => n7505);
   U7118 : BUF_X1 port map( A => n5056, Z => n7508);
   U7119 : BUF_X1 port map( A => n5055, Z => n7511);
   U7120 : BUF_X1 port map( A => n5054, Z => n7514);
   U7121 : BUF_X1 port map( A => n5053, Z => n7517);
   U7122 : BUF_X1 port map( A => n5052, Z => n7520);
   U7123 : BUF_X1 port map( A => n5051, Z => n7523);
   U7124 : BUF_X1 port map( A => n5050, Z => n7526);
   U7125 : BUF_X1 port map( A => n5049, Z => n7529);
   U7126 : BUF_X1 port map( A => n5048, Z => n7532);
   U7127 : BUF_X1 port map( A => n5047, Z => n7535);
   U7128 : BUF_X1 port map( A => n5046, Z => n7538);
   U7129 : BUF_X1 port map( A => n5045, Z => n7541);
   U7130 : BUF_X1 port map( A => n5044, Z => n7544);
   U7131 : BUF_X1 port map( A => n5043, Z => n7547);
   U7132 : BUF_X1 port map( A => n5042, Z => n7550);
   U7133 : BUF_X1 port map( A => n5041, Z => n7553);
   U7134 : BUF_X1 port map( A => n5040, Z => n7556);
   U7135 : BUF_X1 port map( A => n5039, Z => n7559);
   U7136 : BUF_X1 port map( A => n5038, Z => n7562);
   U7137 : BUF_X1 port map( A => n5037, Z => n7565);
   U7138 : BUF_X1 port map( A => n5036, Z => n7568);
   U7139 : BUF_X1 port map( A => n5034, Z => n7580);
   U7140 : BUF_X1 port map( A => n5066, Z => n7477);
   U7141 : BUF_X1 port map( A => n5065, Z => n7480);
   U7142 : BUF_X1 port map( A => n5064, Z => n7483);
   U7143 : BUF_X1 port map( A => n5063, Z => n7486);
   U7144 : BUF_X1 port map( A => n5062, Z => n7489);
   U7145 : BUF_X1 port map( A => n5061, Z => n7492);
   U7146 : BUF_X1 port map( A => n5060, Z => n7495);
   U7147 : BUF_X1 port map( A => n5059, Z => n7498);
   U7148 : BUF_X1 port map( A => n5058, Z => n7501);
   U7149 : BUF_X1 port map( A => n5057, Z => n7504);
   U7150 : BUF_X1 port map( A => n5056, Z => n7507);
   U7151 : BUF_X1 port map( A => n5055, Z => n7510);
   U7152 : BUF_X1 port map( A => n5054, Z => n7513);
   U7153 : BUF_X1 port map( A => n5053, Z => n7516);
   U7154 : BUF_X1 port map( A => n5052, Z => n7519);
   U7155 : BUF_X1 port map( A => n5051, Z => n7522);
   U7156 : BUF_X1 port map( A => n5050, Z => n7525);
   U7157 : BUF_X1 port map( A => n5049, Z => n7528);
   U7158 : BUF_X1 port map( A => n5048, Z => n7531);
   U7159 : BUF_X1 port map( A => n5047, Z => n7534);
   U7160 : BUF_X1 port map( A => n5046, Z => n7537);
   U7161 : BUF_X1 port map( A => n5045, Z => n7540);
   U7162 : BUF_X1 port map( A => n5044, Z => n7543);
   U7163 : BUF_X1 port map( A => n5043, Z => n7546);
   U7164 : BUF_X1 port map( A => n5042, Z => n7549);
   U7165 : BUF_X1 port map( A => n5041, Z => n7552);
   U7166 : BUF_X1 port map( A => n5040, Z => n7555);
   U7167 : BUF_X1 port map( A => n5039, Z => n7558);
   U7168 : BUF_X1 port map( A => n5038, Z => n7561);
   U7169 : BUF_X1 port map( A => n5037, Z => n7564);
   U7170 : BUF_X1 port map( A => n5036, Z => n7567);
   U7171 : BUF_X1 port map( A => n5034, Z => n7579);
   U7172 : BUF_X1 port map( A => n4254, Z => n7584);
   U7173 : BUF_X1 port map( A => n5764, Z => n7089);
   U7174 : BUF_X1 port map( A => n5111, Z => n7191);
   U7175 : BUF_X1 port map( A => n5066, Z => n7479);
   U7176 : BUF_X1 port map( A => n5065, Z => n7482);
   U7177 : BUF_X1 port map( A => n5064, Z => n7485);
   U7178 : BUF_X1 port map( A => n5063, Z => n7488);
   U7179 : BUF_X1 port map( A => n5062, Z => n7491);
   U7180 : BUF_X1 port map( A => n5061, Z => n7494);
   U7181 : BUF_X1 port map( A => n5060, Z => n7497);
   U7182 : BUF_X1 port map( A => n5059, Z => n7500);
   U7183 : BUF_X1 port map( A => n5058, Z => n7503);
   U7184 : BUF_X1 port map( A => n5057, Z => n7506);
   U7185 : BUF_X1 port map( A => n5056, Z => n7509);
   U7186 : BUF_X1 port map( A => n5055, Z => n7512);
   U7187 : BUF_X1 port map( A => n5054, Z => n7515);
   U7188 : BUF_X1 port map( A => n5053, Z => n7518);
   U7189 : BUF_X1 port map( A => n5052, Z => n7521);
   U7190 : BUF_X1 port map( A => n5051, Z => n7524);
   U7191 : BUF_X1 port map( A => n5050, Z => n7527);
   U7192 : BUF_X1 port map( A => n5049, Z => n7530);
   U7193 : BUF_X1 port map( A => n5048, Z => n7533);
   U7194 : BUF_X1 port map( A => n5047, Z => n7536);
   U7195 : BUF_X1 port map( A => n5046, Z => n7539);
   U7196 : BUF_X1 port map( A => n5045, Z => n7542);
   U7197 : BUF_X1 port map( A => n5044, Z => n7545);
   U7198 : BUF_X1 port map( A => n5043, Z => n7548);
   U7199 : BUF_X1 port map( A => n5042, Z => n7551);
   U7200 : BUF_X1 port map( A => n5041, Z => n7554);
   U7201 : BUF_X1 port map( A => n5040, Z => n7557);
   U7202 : BUF_X1 port map( A => n5039, Z => n7560);
   U7203 : BUF_X1 port map( A => n5038, Z => n7563);
   U7204 : BUF_X1 port map( A => n5037, Z => n7566);
   U7205 : BUF_X1 port map( A => n5036, Z => n7569);
   U7206 : BUF_X1 port map( A => n5034, Z => n7581);
   U7207 : NAND2_X1 port map( A1 => n6400, A2 => n6412, ZN => n5805);
   U7208 : NAND2_X1 port map( A1 => n5747, A2 => n5759, ZN => n5152);
   U7209 : NAND2_X1 port map( A1 => n6401, A2 => n6412, ZN => n5804);
   U7210 : NAND2_X1 port map( A1 => n5748, A2 => n5759, ZN => n5151);
   U7211 : NAND2_X1 port map( A1 => n6415, A2 => n6396, ZN => n5809);
   U7212 : NAND2_X1 port map( A1 => n6415, A2 => n6395, ZN => n5810);
   U7213 : NAND2_X1 port map( A1 => n6415, A2 => n6401, ZN => n5814);
   U7214 : NAND2_X1 port map( A1 => n6415, A2 => n6400, ZN => n5815);
   U7215 : NAND2_X1 port map( A1 => n5762, A2 => n5743, ZN => n5156);
   U7216 : NAND2_X1 port map( A1 => n5762, A2 => n5742, ZN => n5157);
   U7217 : NAND2_X1 port map( A1 => n5762, A2 => n5748, ZN => n5161);
   U7218 : NAND2_X1 port map( A1 => n5762, A2 => n5747, ZN => n5162);
   U7219 : NAND2_X1 port map( A1 => n6394, A2 => n6400, ZN => n5781);
   U7220 : NAND2_X1 port map( A1 => n6405, A2 => n6400, ZN => n5791);
   U7221 : NAND2_X1 port map( A1 => n5741, A2 => n5747, ZN => n5128);
   U7222 : NAND2_X1 port map( A1 => n5752, A2 => n5747, ZN => n5138);
   U7223 : NAND2_X1 port map( A1 => n6394, A2 => n6401, ZN => n5780);
   U7224 : NAND2_X1 port map( A1 => n6405, A2 => n6401, ZN => n5790);
   U7225 : NAND2_X1 port map( A1 => n5741, A2 => n5748, ZN => n5127);
   U7226 : NAND2_X1 port map( A1 => n5752, A2 => n5748, ZN => n5137);
   U7227 : NAND2_X1 port map( A1 => n6396, A2 => n6412, ZN => n5799);
   U7228 : NAND2_X1 port map( A1 => n6395, A2 => n6412, ZN => n5800);
   U7229 : NAND2_X1 port map( A1 => n5743, A2 => n5759, ZN => n5146);
   U7230 : NAND2_X1 port map( A1 => n5742, A2 => n5759, ZN => n5147);
   U7231 : NAND2_X1 port map( A1 => n6394, A2 => n6396, ZN => n5775);
   U7232 : NAND2_X1 port map( A1 => n6394, A2 => n6395, ZN => n5776);
   U7233 : NAND2_X1 port map( A1 => n6405, A2 => n6396, ZN => n5785);
   U7234 : NAND2_X1 port map( A1 => n6405, A2 => n6395, ZN => n5786);
   U7235 : NAND2_X1 port map( A1 => n5741, A2 => n5743, ZN => n5122);
   U7236 : NAND2_X1 port map( A1 => n5741, A2 => n5742, ZN => n5123);
   U7237 : NAND2_X1 port map( A1 => n5752, A2 => n5743, ZN => n5132);
   U7238 : NAND2_X1 port map( A1 => n5752, A2 => n5742, ZN => n5133);
   U7239 : AND2_X1 port map( A1 => n6415, A2 => n6398, ZN => n5806);
   U7240 : AND2_X1 port map( A1 => n6415, A2 => n6397, ZN => n5807);
   U7241 : AND2_X1 port map( A1 => n6415, A2 => n6403, ZN => n5811);
   U7242 : AND2_X1 port map( A1 => n6415, A2 => n6402, ZN => n5812);
   U7243 : AND2_X1 port map( A1 => n5762, A2 => n5745, ZN => n5153);
   U7244 : AND2_X1 port map( A1 => n5762, A2 => n5744, ZN => n5154);
   U7245 : AND2_X1 port map( A1 => n5762, A2 => n5750, ZN => n5158);
   U7246 : AND2_X1 port map( A1 => n5762, A2 => n5749, ZN => n5159);
   U7247 : AND2_X1 port map( A1 => n6398, A2 => n6412, ZN => n5796);
   U7248 : AND2_X1 port map( A1 => n6397, A2 => n6412, ZN => n5797);
   U7249 : AND2_X1 port map( A1 => n6403, A2 => n6412, ZN => n5801);
   U7250 : AND2_X1 port map( A1 => n6402, A2 => n6412, ZN => n5802);
   U7251 : AND2_X1 port map( A1 => n5745, A2 => n5759, ZN => n5143);
   U7252 : AND2_X1 port map( A1 => n5744, A2 => n5759, ZN => n5144);
   U7253 : AND2_X1 port map( A1 => n5750, A2 => n5759, ZN => n5148);
   U7254 : AND2_X1 port map( A1 => n5749, A2 => n5759, ZN => n5149);
   U7255 : AND2_X1 port map( A1 => n6394, A2 => n6403, ZN => n5777);
   U7256 : AND2_X1 port map( A1 => n6394, A2 => n6402, ZN => n5778);
   U7257 : AND2_X1 port map( A1 => n6405, A2 => n6403, ZN => n5787);
   U7258 : AND2_X1 port map( A1 => n6405, A2 => n6402, ZN => n5788);
   U7259 : AND2_X1 port map( A1 => n5741, A2 => n5750, ZN => n5124);
   U7260 : AND2_X1 port map( A1 => n5741, A2 => n5749, ZN => n5125);
   U7261 : AND2_X1 port map( A1 => n5752, A2 => n5750, ZN => n5134);
   U7262 : AND2_X1 port map( A1 => n5752, A2 => n5749, ZN => n5135);
   U7263 : AND2_X1 port map( A1 => n6394, A2 => n6398, ZN => n5772);
   U7264 : AND2_X1 port map( A1 => n6394, A2 => n6397, ZN => n5773);
   U7265 : AND2_X1 port map( A1 => n6405, A2 => n6398, ZN => n5782);
   U7266 : AND2_X1 port map( A1 => n6405, A2 => n6397, ZN => n5783);
   U7267 : AND2_X1 port map( A1 => n5741, A2 => n5745, ZN => n5119);
   U7268 : AND2_X1 port map( A1 => n5741, A2 => n5744, ZN => n5120);
   U7269 : AND2_X1 port map( A1 => n5752, A2 => n5745, ZN => n5129);
   U7270 : AND2_X1 port map( A1 => n5752, A2 => n5744, ZN => n5130);
   U7271 : BUF_X1 port map( A => n5110, Z => n7197);
   U7272 : OAI21_X1 port map( B1 => n5082, B2 => n5103, A => n7587, ZN => n5110
                           );
   U7273 : INV_X1 port map( A => n5109, ZN => n7215);
   U7274 : OAI21_X1 port map( B1 => n5080, B2 => n5103, A => n7584, ZN => n5109
                           );
   U7275 : INV_X1 port map( A => n5108, ZN => n7224);
   U7276 : OAI21_X1 port map( B1 => n5078, B2 => n5103, A => n7584, ZN => n5108
                           );
   U7277 : INV_X1 port map( A => n5107, ZN => n7233);
   U7278 : OAI21_X1 port map( B1 => n5076, B2 => n5103, A => n7584, ZN => n5107
                           );
   U7279 : INV_X1 port map( A => n5106, ZN => n7242);
   U7280 : OAI21_X1 port map( B1 => n5074, B2 => n5103, A => n7585, ZN => n5106
                           );
   U7281 : INV_X1 port map( A => n5105, ZN => n7251);
   U7282 : OAI21_X1 port map( B1 => n5072, B2 => n5103, A => n7585, ZN => n5105
                           );
   U7283 : INV_X1 port map( A => n5104, ZN => n7260);
   U7284 : OAI21_X1 port map( B1 => n5070, B2 => n5103, A => n7585, ZN => n5104
                           );
   U7285 : INV_X1 port map( A => n5102, ZN => n7269);
   U7286 : OAI21_X1 port map( B1 => n5068, B2 => n5103, A => n7585, ZN => n5102
                           );
   U7287 : INV_X1 port map( A => n5101, ZN => n7278);
   U7288 : OAI21_X1 port map( B1 => n5082, B2 => n5094, A => n7585, ZN => n5101
                           );
   U7289 : INV_X1 port map( A => n5100, ZN => n7287);
   U7290 : OAI21_X1 port map( B1 => n5080, B2 => n5094, A => n7585, ZN => n5100
                           );
   U7291 : INV_X1 port map( A => n5099, ZN => n7296);
   U7292 : OAI21_X1 port map( B1 => n5078, B2 => n5094, A => n7585, ZN => n5099
                           );
   U7293 : INV_X1 port map( A => n5098, ZN => n7305);
   U7294 : OAI21_X1 port map( B1 => n5076, B2 => n5094, A => n7585, ZN => n5098
                           );
   U7295 : INV_X1 port map( A => n5097, ZN => n7314);
   U7296 : OAI21_X1 port map( B1 => n5074, B2 => n5094, A => n7585, ZN => n5097
                           );
   U7297 : INV_X1 port map( A => n5096, ZN => n7323);
   U7298 : OAI21_X1 port map( B1 => n5072, B2 => n5094, A => n7585, ZN => n5096
                           );
   U7299 : INV_X1 port map( A => n5095, ZN => n7332);
   U7300 : OAI21_X1 port map( B1 => n5070, B2 => n5094, A => n7585, ZN => n5095
                           );
   U7301 : INV_X1 port map( A => n5093, ZN => n7341);
   U7302 : OAI21_X1 port map( B1 => n5068, B2 => n5094, A => n7585, ZN => n5093
                           );
   U7303 : INV_X1 port map( A => n5092, ZN => n7350);
   U7304 : OAI21_X1 port map( B1 => n5082, B2 => n5085, A => n7585, ZN => n5092
                           );
   U7305 : INV_X1 port map( A => n5091, ZN => n7359);
   U7306 : OAI21_X1 port map( B1 => n5080, B2 => n5085, A => n7586, ZN => n5091
                           );
   U7307 : INV_X1 port map( A => n5090, ZN => n7368);
   U7308 : OAI21_X1 port map( B1 => n5078, B2 => n5085, A => n7586, ZN => n5090
                           );
   U7309 : INV_X1 port map( A => n5089, ZN => n7377);
   U7310 : OAI21_X1 port map( B1 => n5076, B2 => n5085, A => n7586, ZN => n5089
                           );
   U7311 : INV_X1 port map( A => n5088, ZN => n7386);
   U7312 : OAI21_X1 port map( B1 => n5074, B2 => n5085, A => n7586, ZN => n5088
                           );
   U7313 : INV_X1 port map( A => n5087, ZN => n7395);
   U7314 : OAI21_X1 port map( B1 => n5072, B2 => n5085, A => n7586, ZN => n5087
                           );
   U7315 : INV_X1 port map( A => n5086, ZN => n7404);
   U7316 : OAI21_X1 port map( B1 => n5070, B2 => n5085, A => n7586, ZN => n5086
                           );
   U7317 : INV_X1 port map( A => n5084, ZN => n7413);
   U7318 : OAI21_X1 port map( B1 => n5068, B2 => n5085, A => n7586, ZN => n5084
                           );
   U7319 : INV_X1 port map( A => n5081, ZN => n7422);
   U7320 : OAI21_X1 port map( B1 => n5067, B2 => n5082, A => n7586, ZN => n5081
                           );
   U7321 : INV_X1 port map( A => n5079, ZN => n7431);
   U7322 : OAI21_X1 port map( B1 => n5067, B2 => n5080, A => n7586, ZN => n5079
                           );
   U7323 : INV_X1 port map( A => n5077, ZN => n7440);
   U7324 : OAI21_X1 port map( B1 => n5067, B2 => n5078, A => n7586, ZN => n5077
                           );
   U7325 : INV_X1 port map( A => n5075, ZN => n7449);
   U7326 : OAI21_X1 port map( B1 => n5067, B2 => n5076, A => n7586, ZN => n5075
                           );
   U7327 : INV_X1 port map( A => n5073, ZN => n7458);
   U7328 : OAI21_X1 port map( B1 => n5067, B2 => n5074, A => n7586, ZN => n5073
                           );
   U7329 : INV_X1 port map( A => n5071, ZN => n7467);
   U7330 : OAI21_X1 port map( B1 => n5067, B2 => n5072, A => n7586, ZN => n5071
                           );
   U7331 : INV_X1 port map( A => n5069, ZN => n7476);
   U7332 : OAI21_X1 port map( B1 => n5067, B2 => n5070, A => n7587, ZN => n5069
                           );
   U7333 : AOI221_X1 port map( B1 => n7074, B2 => n6433, C1 => n7071, C2 => 
                           n6441, A => n6399, ZN => n6391);
   U7334 : OAI22_X1 port map( A1 => n832, A2 => n7068, B1 => n800, B2 => n7065,
                           ZN => n6399);
   U7335 : AOI221_X1 port map( B1 => n7026, B2 => n6497, C1 => n7023, C2 => 
                           n6505, A => n6413, ZN => n6409);
   U7336 : OAI22_X1 port map( A1 => n320, A2 => n7020, B1 => n288, B2 => n7017,
                           ZN => n6413);
   U7337 : AOI221_X1 port map( B1 => n7074, B2 => n6434, C1 => n7071, C2 => 
                           n6442, A => n6375, ZN => n6372);
   U7338 : OAI22_X1 port map( A1 => n831, A2 => n7068, B1 => n799, B2 => n7065,
                           ZN => n6375);
   U7339 : AOI221_X1 port map( B1 => n7026, B2 => n6498, C1 => n7023, C2 => 
                           n6506, A => n6383, ZN => n6380);
   U7340 : OAI22_X1 port map( A1 => n319, A2 => n7020, B1 => n287, B2 => n7017,
                           ZN => n6383);
   U7341 : AOI221_X1 port map( B1 => n7074, B2 => n6435, C1 => n7071, C2 => 
                           n6443, A => n6356, ZN => n6353);
   U7342 : OAI22_X1 port map( A1 => n830, A2 => n7068, B1 => n798, B2 => n7065,
                           ZN => n6356);
   U7343 : AOI221_X1 port map( B1 => n7026, B2 => n6499, C1 => n7023, C2 => 
                           n6507, A => n6364, ZN => n6361);
   U7344 : OAI22_X1 port map( A1 => n318, A2 => n7020, B1 => n286, B2 => n7017,
                           ZN => n6364);
   U7345 : AOI221_X1 port map( B1 => n7074, B2 => n6436, C1 => n7071, C2 => 
                           n6444, A => n6337, ZN => n6334);
   U7346 : OAI22_X1 port map( A1 => n829, A2 => n7068, B1 => n797, B2 => n7065,
                           ZN => n6337);
   U7347 : AOI221_X1 port map( B1 => n7026, B2 => n6500, C1 => n7023, C2 => 
                           n6508, A => n6345, ZN => n6342);
   U7348 : OAI22_X1 port map( A1 => n317, A2 => n7020, B1 => n285, B2 => n7017,
                           ZN => n6345);
   U7349 : AOI221_X1 port map( B1 => n7074, B2 => n6437, C1 => n7071, C2 => 
                           n6445, A => n6318, ZN => n6315);
   U7350 : OAI22_X1 port map( A1 => n828, A2 => n7068, B1 => n796, B2 => n7065,
                           ZN => n6318);
   U7351 : AOI221_X1 port map( B1 => n7026, B2 => n6501, C1 => n7023, C2 => 
                           n6509, A => n6326, ZN => n6323);
   U7352 : OAI22_X1 port map( A1 => n316, A2 => n7020, B1 => n284, B2 => n7017,
                           ZN => n6326);
   U7353 : AOI221_X1 port map( B1 => n7074, B2 => n6438, C1 => n7071, C2 => 
                           n6446, A => n6299, ZN => n6296);
   U7354 : OAI22_X1 port map( A1 => n827, A2 => n7068, B1 => n795, B2 => n7065,
                           ZN => n6299);
   U7355 : AOI221_X1 port map( B1 => n7026, B2 => n6502, C1 => n7023, C2 => 
                           n6510, A => n6307, ZN => n6304);
   U7356 : OAI22_X1 port map( A1 => n315, A2 => n7020, B1 => n283, B2 => n7017,
                           ZN => n6307);
   U7357 : AOI221_X1 port map( B1 => n7074, B2 => n6439, C1 => n7071, C2 => 
                           n6447, A => n6280, ZN => n6277);
   U7358 : OAI22_X1 port map( A1 => n826, A2 => n7068, B1 => n794, B2 => n7065,
                           ZN => n6280);
   U7359 : AOI221_X1 port map( B1 => n7026, B2 => n6503, C1 => n7023, C2 => 
                           n6511, A => n6288, ZN => n6285);
   U7360 : OAI22_X1 port map( A1 => n314, A2 => n7020, B1 => n282, B2 => n7017,
                           ZN => n6288);
   U7361 : AOI221_X1 port map( B1 => n7074, B2 => n6440, C1 => n7071, C2 => 
                           n6448, A => n6261, ZN => n6258);
   U7362 : OAI22_X1 port map( A1 => n825, A2 => n7068, B1 => n793, B2 => n7065,
                           ZN => n6261);
   U7363 : AOI221_X1 port map( B1 => n7026, B2 => n6504, C1 => n7023, C2 => 
                           n6512, A => n6269, ZN => n6266);
   U7364 : OAI22_X1 port map( A1 => n313, A2 => n7020, B1 => n281, B2 => n7017,
                           ZN => n6269);
   U7365 : AOI221_X1 port map( B1 => n7074, B2 => n6593, C1 => n7071, C2 => 
                           n6617, A => n6242, ZN => n6239);
   U7366 : OAI22_X1 port map( A1 => n824, A2 => n7068, B1 => n792, B2 => n7065,
                           ZN => n6242);
   U7367 : AOI221_X1 port map( B1 => n7026, B2 => n6785, C1 => n7023, C2 => 
                           n6809, A => n6250, ZN => n6247);
   U7368 : OAI22_X1 port map( A1 => n312, A2 => n7020, B1 => n280, B2 => n7017,
                           ZN => n6250);
   U7369 : AOI221_X1 port map( B1 => n7074, B2 => n6594, C1 => n7071, C2 => 
                           n6618, A => n6223, ZN => n6220);
   U7370 : OAI22_X1 port map( A1 => n823, A2 => n7068, B1 => n791, B2 => n7065,
                           ZN => n6223);
   U7371 : AOI221_X1 port map( B1 => n7026, B2 => n6786, C1 => n7023, C2 => 
                           n6810, A => n6231, ZN => n6228);
   U7372 : OAI22_X1 port map( A1 => n311, A2 => n7020, B1 => n279, B2 => n7017,
                           ZN => n6231);
   U7373 : AOI221_X1 port map( B1 => n7074, B2 => n6595, C1 => n7071, C2 => 
                           n6619, A => n6204, ZN => n6201);
   U7374 : OAI22_X1 port map( A1 => n822, A2 => n7068, B1 => n790, B2 => n7065,
                           ZN => n6204);
   U7375 : AOI221_X1 port map( B1 => n7026, B2 => n6787, C1 => n7023, C2 => 
                           n6811, A => n6212, ZN => n6209);
   U7376 : OAI22_X1 port map( A1 => n310, A2 => n7020, B1 => n278, B2 => n7017,
                           ZN => n6212);
   U7377 : AOI221_X1 port map( B1 => n7074, B2 => n6596, C1 => n7071, C2 => 
                           n6620, A => n6185, ZN => n6182);
   U7378 : OAI22_X1 port map( A1 => n821, A2 => n7068, B1 => n789, B2 => n7065,
                           ZN => n6185);
   U7379 : AOI221_X1 port map( B1 => n7026, B2 => n6788, C1 => n7023, C2 => 
                           n6812, A => n6193, ZN => n6190);
   U7380 : OAI22_X1 port map( A1 => n309, A2 => n7020, B1 => n277, B2 => n7017,
                           ZN => n6193);
   U7381 : AOI221_X1 port map( B1 => n7075, B2 => n6597, C1 => n7072, C2 => 
                           n6621, A => n6166, ZN => n6163);
   U7382 : OAI22_X1 port map( A1 => n820, A2 => n7069, B1 => n788, B2 => n7066,
                           ZN => n6166);
   U7383 : AOI221_X1 port map( B1 => n7027, B2 => n6789, C1 => n7024, C2 => 
                           n6813, A => n6174, ZN => n6171);
   U7384 : OAI22_X1 port map( A1 => n308, A2 => n7021, B1 => n276, B2 => n7018,
                           ZN => n6174);
   U7385 : AOI221_X1 port map( B1 => n7075, B2 => n6598, C1 => n7072, C2 => 
                           n6622, A => n6147, ZN => n6144);
   U7386 : OAI22_X1 port map( A1 => n819, A2 => n7069, B1 => n787, B2 => n7066,
                           ZN => n6147);
   U7387 : AOI221_X1 port map( B1 => n7027, B2 => n6790, C1 => n7024, C2 => 
                           n6814, A => n6155, ZN => n6152);
   U7388 : OAI22_X1 port map( A1 => n307, A2 => n7021, B1 => n275, B2 => n7018,
                           ZN => n6155);
   U7389 : AOI221_X1 port map( B1 => n7075, B2 => n6599, C1 => n7072, C2 => 
                           n6623, A => n6128, ZN => n6125);
   U7390 : OAI22_X1 port map( A1 => n818, A2 => n7069, B1 => n786, B2 => n7066,
                           ZN => n6128);
   U7391 : AOI221_X1 port map( B1 => n7027, B2 => n6791, C1 => n7024, C2 => 
                           n6815, A => n6136, ZN => n6133);
   U7392 : OAI22_X1 port map( A1 => n306, A2 => n7021, B1 => n274, B2 => n7018,
                           ZN => n6136);
   U7393 : AOI221_X1 port map( B1 => n7075, B2 => n6600, C1 => n7072, C2 => 
                           n6624, A => n6109, ZN => n6106);
   U7394 : OAI22_X1 port map( A1 => n817, A2 => n7069, B1 => n785, B2 => n7066,
                           ZN => n6109);
   U7395 : AOI221_X1 port map( B1 => n7027, B2 => n6792, C1 => n7024, C2 => 
                           n6816, A => n6117, ZN => n6114);
   U7396 : OAI22_X1 port map( A1 => n305, A2 => n7021, B1 => n273, B2 => n7018,
                           ZN => n6117);
   U7397 : AOI221_X1 port map( B1 => n7075, B2 => n6601, C1 => n7072, C2 => 
                           n6625, A => n6090, ZN => n6087);
   U7398 : OAI22_X1 port map( A1 => n816, A2 => n7069, B1 => n784, B2 => n7066,
                           ZN => n6090);
   U7399 : AOI221_X1 port map( B1 => n7027, B2 => n6793, C1 => n7024, C2 => 
                           n6817, A => n6098, ZN => n6095);
   U7400 : OAI22_X1 port map( A1 => n304, A2 => n7021, B1 => n272, B2 => n7018,
                           ZN => n6098);
   U7401 : AOI221_X1 port map( B1 => n7075, B2 => n6602, C1 => n7072, C2 => 
                           n6626, A => n6071, ZN => n6068);
   U7402 : OAI22_X1 port map( A1 => n815, A2 => n7069, B1 => n783, B2 => n7066,
                           ZN => n6071);
   U7403 : AOI221_X1 port map( B1 => n7027, B2 => n6794, C1 => n7024, C2 => 
                           n6818, A => n6079, ZN => n6076);
   U7404 : OAI22_X1 port map( A1 => n303, A2 => n7021, B1 => n271, B2 => n7018,
                           ZN => n6079);
   U7405 : AOI221_X1 port map( B1 => n7075, B2 => n6603, C1 => n7072, C2 => 
                           n6627, A => n6052, ZN => n6049);
   U7406 : OAI22_X1 port map( A1 => n814, A2 => n7069, B1 => n782, B2 => n7066,
                           ZN => n6052);
   U7407 : AOI221_X1 port map( B1 => n7027, B2 => n6795, C1 => n7024, C2 => 
                           n6819, A => n6060, ZN => n6057);
   U7408 : OAI22_X1 port map( A1 => n302, A2 => n7021, B1 => n270, B2 => n7018,
                           ZN => n6060);
   U7409 : AOI221_X1 port map( B1 => n7075, B2 => n6604, C1 => n7072, C2 => 
                           n6628, A => n6033, ZN => n6030);
   U7410 : OAI22_X1 port map( A1 => n813, A2 => n7069, B1 => n781, B2 => n7066,
                           ZN => n6033);
   U7411 : AOI221_X1 port map( B1 => n7027, B2 => n6796, C1 => n7024, C2 => 
                           n6820, A => n6041, ZN => n6038);
   U7412 : OAI22_X1 port map( A1 => n301, A2 => n7021, B1 => n269, B2 => n7018,
                           ZN => n6041);
   U7413 : AOI221_X1 port map( B1 => n7075, B2 => n6605, C1 => n7072, C2 => 
                           n6629, A => n6014, ZN => n6011);
   U7414 : OAI22_X1 port map( A1 => n812, A2 => n7069, B1 => n780, B2 => n7066,
                           ZN => n6014);
   U7415 : AOI221_X1 port map( B1 => n7027, B2 => n6797, C1 => n7024, C2 => 
                           n6821, A => n6022, ZN => n6019);
   U7416 : OAI22_X1 port map( A1 => n300, A2 => n7021, B1 => n268, B2 => n7018,
                           ZN => n6022);
   U7417 : AOI221_X1 port map( B1 => n7075, B2 => n6606, C1 => n7072, C2 => 
                           n6630, A => n5995, ZN => n5992);
   U7418 : OAI22_X1 port map( A1 => n811, A2 => n7069, B1 => n779, B2 => n7066,
                           ZN => n5995);
   U7419 : AOI221_X1 port map( B1 => n7027, B2 => n6798, C1 => n7024, C2 => 
                           n6822, A => n6003, ZN => n6000);
   U7420 : OAI22_X1 port map( A1 => n299, A2 => n7021, B1 => n267, B2 => n7018,
                           ZN => n6003);
   U7421 : AOI221_X1 port map( B1 => n7075, B2 => n6607, C1 => n7072, C2 => 
                           n6631, A => n5976, ZN => n5973);
   U7422 : OAI22_X1 port map( A1 => n810, A2 => n7069, B1 => n778, B2 => n7066,
                           ZN => n5976);
   U7423 : AOI221_X1 port map( B1 => n7027, B2 => n6799, C1 => n7024, C2 => 
                           n6823, A => n5984, ZN => n5981);
   U7424 : OAI22_X1 port map( A1 => n298, A2 => n7021, B1 => n266, B2 => n7018,
                           ZN => n5984);
   U7425 : AOI221_X1 port map( B1 => n7075, B2 => n6608, C1 => n7072, C2 => 
                           n6632, A => n5957, ZN => n5954);
   U7426 : OAI22_X1 port map( A1 => n809, A2 => n7069, B1 => n777, B2 => n7066,
                           ZN => n5957);
   U7427 : AOI221_X1 port map( B1 => n7027, B2 => n6800, C1 => n7024, C2 => 
                           n6824, A => n5965, ZN => n5962);
   U7428 : OAI22_X1 port map( A1 => n297, A2 => n7021, B1 => n265, B2 => n7018,
                           ZN => n5965);
   U7429 : AOI221_X1 port map( B1 => n7076, B2 => n6609, C1 => n7073, C2 => 
                           n6633, A => n5938, ZN => n5935);
   U7430 : OAI22_X1 port map( A1 => n808, A2 => n7070, B1 => n776, B2 => n7067,
                           ZN => n5938);
   U7431 : AOI221_X1 port map( B1 => n7028, B2 => n6801, C1 => n7025, C2 => 
                           n6825, A => n5946, ZN => n5943);
   U7432 : OAI22_X1 port map( A1 => n296, A2 => n7022, B1 => n264, B2 => n7019,
                           ZN => n5946);
   U7433 : AOI221_X1 port map( B1 => n7076, B2 => n6610, C1 => n7073, C2 => 
                           n6634, A => n5919, ZN => n5916);
   U7434 : OAI22_X1 port map( A1 => n807, A2 => n7070, B1 => n775, B2 => n7067,
                           ZN => n5919);
   U7435 : AOI221_X1 port map( B1 => n7028, B2 => n6802, C1 => n7025, C2 => 
                           n6826, A => n5927, ZN => n5924);
   U7436 : OAI22_X1 port map( A1 => n295, A2 => n7022, B1 => n263, B2 => n7019,
                           ZN => n5927);
   U7437 : AOI221_X1 port map( B1 => n7076, B2 => n6611, C1 => n7073, C2 => 
                           n6635, A => n5900, ZN => n5897);
   U7438 : OAI22_X1 port map( A1 => n806, A2 => n7070, B1 => n774, B2 => n7067,
                           ZN => n5900);
   U7439 : AOI221_X1 port map( B1 => n7028, B2 => n6803, C1 => n7025, C2 => 
                           n6827, A => n5908, ZN => n5905);
   U7440 : OAI22_X1 port map( A1 => n294, A2 => n7022, B1 => n262, B2 => n7019,
                           ZN => n5908);
   U7441 : AOI221_X1 port map( B1 => n7076, B2 => n6612, C1 => n7073, C2 => 
                           n6636, A => n5881, ZN => n5878);
   U7442 : OAI22_X1 port map( A1 => n805, A2 => n7070, B1 => n773, B2 => n7067,
                           ZN => n5881);
   U7443 : AOI221_X1 port map( B1 => n7028, B2 => n6804, C1 => n7025, C2 => 
                           n6828, A => n5889, ZN => n5886);
   U7444 : OAI22_X1 port map( A1 => n293, A2 => n7022, B1 => n261, B2 => n7019,
                           ZN => n5889);
   U7445 : AOI221_X1 port map( B1 => n7076, B2 => n6613, C1 => n7073, C2 => 
                           n6637, A => n5862, ZN => n5859);
   U7446 : OAI22_X1 port map( A1 => n804, A2 => n7070, B1 => n772, B2 => n7067,
                           ZN => n5862);
   U7447 : AOI221_X1 port map( B1 => n7028, B2 => n6805, C1 => n7025, C2 => 
                           n6829, A => n5870, ZN => n5867);
   U7448 : OAI22_X1 port map( A1 => n292, A2 => n7022, B1 => n260, B2 => n7019,
                           ZN => n5870);
   U7449 : AOI221_X1 port map( B1 => n7076, B2 => n6614, C1 => n7073, C2 => 
                           n6638, A => n5843, ZN => n5840);
   U7450 : OAI22_X1 port map( A1 => n803, A2 => n7070, B1 => n771, B2 => n7067,
                           ZN => n5843);
   U7451 : AOI221_X1 port map( B1 => n7028, B2 => n6806, C1 => n7025, C2 => 
                           n6830, A => n5851, ZN => n5848);
   U7452 : OAI22_X1 port map( A1 => n291, A2 => n7022, B1 => n259, B2 => n7019,
                           ZN => n5851);
   U7453 : AOI221_X1 port map( B1 => n7076, B2 => n6615, C1 => n7073, C2 => 
                           n6639, A => n5824, ZN => n5821);
   U7454 : OAI22_X1 port map( A1 => n802, A2 => n7070, B1 => n770, B2 => n7067,
                           ZN => n5824);
   U7455 : AOI221_X1 port map( B1 => n7028, B2 => n6807, C1 => n7025, C2 => 
                           n6831, A => n5832, ZN => n5829);
   U7456 : OAI22_X1 port map( A1 => n290, A2 => n7022, B1 => n258, B2 => n7019,
                           ZN => n5832);
   U7457 : AOI221_X1 port map( B1 => n7076, B2 => n6616, C1 => n7073, C2 => 
                           n6640, A => n5779, ZN => n5770);
   U7458 : OAI22_X1 port map( A1 => n801, A2 => n7070, B1 => n769, B2 => n7067,
                           ZN => n5779);
   U7459 : AOI221_X1 port map( B1 => n7028, B2 => n6808, C1 => n7025, C2 => 
                           n6832, A => n5803, ZN => n5794);
   U7460 : OAI22_X1 port map( A1 => n289, A2 => n7022, B1 => n257, B2 => n7019,
                           ZN => n5803);
   U7461 : AOI221_X1 port map( B1 => n7176, B2 => n6433, C1 => n7173, C2 => 
                           n6441, A => n5746, ZN => n5738);
   U7462 : OAI22_X1 port map( A1 => n832, A2 => n7170, B1 => n800, B2 => n7167,
                           ZN => n5746);
   U7463 : AOI221_X1 port map( B1 => n7128, B2 => n6497, C1 => n7125, C2 => 
                           n6505, A => n5760, ZN => n5756);
   U7464 : OAI22_X1 port map( A1 => n320, A2 => n7122, B1 => n288, B2 => n7119,
                           ZN => n5760);
   U7465 : AOI221_X1 port map( B1 => n7176, B2 => n6434, C1 => n7173, C2 => 
                           n6442, A => n5722, ZN => n5719);
   U7466 : OAI22_X1 port map( A1 => n831, A2 => n7170, B1 => n799, B2 => n7167,
                           ZN => n5722);
   U7467 : AOI221_X1 port map( B1 => n7128, B2 => n6498, C1 => n7125, C2 => 
                           n6506, A => n5730, ZN => n5727);
   U7468 : OAI22_X1 port map( A1 => n319, A2 => n7122, B1 => n287, B2 => n7119,
                           ZN => n5730);
   U7469 : AOI221_X1 port map( B1 => n7176, B2 => n6435, C1 => n7173, C2 => 
                           n6443, A => n5703, ZN => n5700);
   U7470 : OAI22_X1 port map( A1 => n830, A2 => n7170, B1 => n798, B2 => n7167,
                           ZN => n5703);
   U7471 : AOI221_X1 port map( B1 => n7128, B2 => n6499, C1 => n7125, C2 => 
                           n6507, A => n5711, ZN => n5708);
   U7472 : OAI22_X1 port map( A1 => n318, A2 => n7122, B1 => n286, B2 => n7119,
                           ZN => n5711);
   U7473 : AOI221_X1 port map( B1 => n7176, B2 => n6436, C1 => n7173, C2 => 
                           n6444, A => n5684, ZN => n5681);
   U7474 : OAI22_X1 port map( A1 => n829, A2 => n7170, B1 => n797, B2 => n7167,
                           ZN => n5684);
   U7475 : AOI221_X1 port map( B1 => n7128, B2 => n6500, C1 => n7125, C2 => 
                           n6508, A => n5692, ZN => n5689);
   U7476 : OAI22_X1 port map( A1 => n317, A2 => n7122, B1 => n285, B2 => n7119,
                           ZN => n5692);
   U7477 : AOI221_X1 port map( B1 => n7176, B2 => n6437, C1 => n7173, C2 => 
                           n6445, A => n5665, ZN => n5662);
   U7478 : OAI22_X1 port map( A1 => n828, A2 => n7170, B1 => n796, B2 => n7167,
                           ZN => n5665);
   U7479 : AOI221_X1 port map( B1 => n7128, B2 => n6501, C1 => n7125, C2 => 
                           n6509, A => n5673, ZN => n5670);
   U7480 : OAI22_X1 port map( A1 => n316, A2 => n7122, B1 => n284, B2 => n7119,
                           ZN => n5673);
   U7481 : AOI221_X1 port map( B1 => n7176, B2 => n6438, C1 => n7173, C2 => 
                           n6446, A => n5646, ZN => n5643);
   U7482 : OAI22_X1 port map( A1 => n827, A2 => n7170, B1 => n795, B2 => n7167,
                           ZN => n5646);
   U7483 : AOI221_X1 port map( B1 => n7128, B2 => n6502, C1 => n7125, C2 => 
                           n6510, A => n5654, ZN => n5651);
   U7484 : OAI22_X1 port map( A1 => n315, A2 => n7122, B1 => n283, B2 => n7119,
                           ZN => n5654);
   U7485 : AOI221_X1 port map( B1 => n7176, B2 => n6439, C1 => n7173, C2 => 
                           n6447, A => n5627, ZN => n5624);
   U7486 : OAI22_X1 port map( A1 => n826, A2 => n7170, B1 => n794, B2 => n7167,
                           ZN => n5627);
   U7487 : AOI221_X1 port map( B1 => n7128, B2 => n6503, C1 => n7125, C2 => 
                           n6511, A => n5635, ZN => n5632);
   U7488 : OAI22_X1 port map( A1 => n314, A2 => n7122, B1 => n282, B2 => n7119,
                           ZN => n5635);
   U7489 : AOI221_X1 port map( B1 => n7176, B2 => n6440, C1 => n7173, C2 => 
                           n6448, A => n5608, ZN => n5605);
   U7490 : OAI22_X1 port map( A1 => n825, A2 => n7170, B1 => n793, B2 => n7167,
                           ZN => n5608);
   U7491 : AOI221_X1 port map( B1 => n7128, B2 => n6504, C1 => n7125, C2 => 
                           n6512, A => n5616, ZN => n5613);
   U7492 : OAI22_X1 port map( A1 => n313, A2 => n7122, B1 => n281, B2 => n7119,
                           ZN => n5616);
   U7493 : AOI221_X1 port map( B1 => n7176, B2 => n6593, C1 => n7173, C2 => 
                           n6617, A => n5589, ZN => n5586);
   U7494 : OAI22_X1 port map( A1 => n824, A2 => n7170, B1 => n792, B2 => n7167,
                           ZN => n5589);
   U7495 : AOI221_X1 port map( B1 => n7128, B2 => n6785, C1 => n7125, C2 => 
                           n6809, A => n5597, ZN => n5594);
   U7496 : OAI22_X1 port map( A1 => n312, A2 => n7122, B1 => n280, B2 => n7119,
                           ZN => n5597);
   U7497 : AOI221_X1 port map( B1 => n7176, B2 => n6594, C1 => n7173, C2 => 
                           n6618, A => n5570, ZN => n5567);
   U7498 : OAI22_X1 port map( A1 => n823, A2 => n7170, B1 => n791, B2 => n7167,
                           ZN => n5570);
   U7499 : AOI221_X1 port map( B1 => n7128, B2 => n6786, C1 => n7125, C2 => 
                           n6810, A => n5578, ZN => n5575);
   U7500 : OAI22_X1 port map( A1 => n311, A2 => n7122, B1 => n279, B2 => n7119,
                           ZN => n5578);
   U7501 : AOI221_X1 port map( B1 => n7176, B2 => n6595, C1 => n7173, C2 => 
                           n6619, A => n5551, ZN => n5548);
   U7502 : OAI22_X1 port map( A1 => n822, A2 => n7170, B1 => n790, B2 => n7167,
                           ZN => n5551);
   U7503 : AOI221_X1 port map( B1 => n7128, B2 => n6787, C1 => n7125, C2 => 
                           n6811, A => n5559, ZN => n5556);
   U7504 : OAI22_X1 port map( A1 => n310, A2 => n7122, B1 => n278, B2 => n7119,
                           ZN => n5559);
   U7505 : AOI221_X1 port map( B1 => n7176, B2 => n6596, C1 => n7173, C2 => 
                           n6620, A => n5532, ZN => n5529);
   U7506 : OAI22_X1 port map( A1 => n821, A2 => n7170, B1 => n789, B2 => n7167,
                           ZN => n5532);
   U7507 : AOI221_X1 port map( B1 => n7128, B2 => n6788, C1 => n7125, C2 => 
                           n6812, A => n5540, ZN => n5537);
   U7508 : OAI22_X1 port map( A1 => n309, A2 => n7122, B1 => n277, B2 => n7119,
                           ZN => n5540);
   U7509 : AOI221_X1 port map( B1 => n7177, B2 => n6597, C1 => n7174, C2 => 
                           n6621, A => n5513, ZN => n5510);
   U7510 : OAI22_X1 port map( A1 => n820, A2 => n7171, B1 => n788, B2 => n7168,
                           ZN => n5513);
   U7511 : AOI221_X1 port map( B1 => n7129, B2 => n6789, C1 => n7126, C2 => 
                           n6813, A => n5521, ZN => n5518);
   U7512 : OAI22_X1 port map( A1 => n308, A2 => n7123, B1 => n276, B2 => n7120,
                           ZN => n5521);
   U7513 : AOI221_X1 port map( B1 => n7177, B2 => n6598, C1 => n7174, C2 => 
                           n6622, A => n5494, ZN => n5491);
   U7514 : OAI22_X1 port map( A1 => n819, A2 => n7171, B1 => n787, B2 => n7168,
                           ZN => n5494);
   U7515 : AOI221_X1 port map( B1 => n7129, B2 => n6790, C1 => n7126, C2 => 
                           n6814, A => n5502, ZN => n5499);
   U7516 : OAI22_X1 port map( A1 => n307, A2 => n7123, B1 => n275, B2 => n7120,
                           ZN => n5502);
   U7517 : AOI221_X1 port map( B1 => n7177, B2 => n6599, C1 => n7174, C2 => 
                           n6623, A => n5475, ZN => n5472);
   U7518 : OAI22_X1 port map( A1 => n818, A2 => n7171, B1 => n786, B2 => n7168,
                           ZN => n5475);
   U7519 : AOI221_X1 port map( B1 => n7129, B2 => n6791, C1 => n7126, C2 => 
                           n6815, A => n5483, ZN => n5480);
   U7520 : OAI22_X1 port map( A1 => n306, A2 => n7123, B1 => n274, B2 => n7120,
                           ZN => n5483);
   U7521 : AOI221_X1 port map( B1 => n7177, B2 => n6600, C1 => n7174, C2 => 
                           n6624, A => n5456, ZN => n5453);
   U7522 : OAI22_X1 port map( A1 => n817, A2 => n7171, B1 => n785, B2 => n7168,
                           ZN => n5456);
   U7523 : AOI221_X1 port map( B1 => n7129, B2 => n6792, C1 => n7126, C2 => 
                           n6816, A => n5464, ZN => n5461);
   U7524 : OAI22_X1 port map( A1 => n305, A2 => n7123, B1 => n273, B2 => n7120,
                           ZN => n5464);
   U7525 : AOI221_X1 port map( B1 => n7177, B2 => n6601, C1 => n7174, C2 => 
                           n6625, A => n5437, ZN => n5434);
   U7526 : OAI22_X1 port map( A1 => n816, A2 => n7171, B1 => n784, B2 => n7168,
                           ZN => n5437);
   U7527 : AOI221_X1 port map( B1 => n7129, B2 => n6793, C1 => n7126, C2 => 
                           n6817, A => n5445, ZN => n5442);
   U7528 : OAI22_X1 port map( A1 => n304, A2 => n7123, B1 => n272, B2 => n7120,
                           ZN => n5445);
   U7529 : AOI221_X1 port map( B1 => n7177, B2 => n6602, C1 => n7174, C2 => 
                           n6626, A => n5418, ZN => n5415);
   U7530 : OAI22_X1 port map( A1 => n815, A2 => n7171, B1 => n783, B2 => n7168,
                           ZN => n5418);
   U7531 : AOI221_X1 port map( B1 => n7129, B2 => n6794, C1 => n7126, C2 => 
                           n6818, A => n5426, ZN => n5423);
   U7532 : OAI22_X1 port map( A1 => n303, A2 => n7123, B1 => n271, B2 => n7120,
                           ZN => n5426);
   U7533 : AOI221_X1 port map( B1 => n7177, B2 => n6603, C1 => n7174, C2 => 
                           n6627, A => n5399, ZN => n5396);
   U7534 : OAI22_X1 port map( A1 => n814, A2 => n7171, B1 => n782, B2 => n7168,
                           ZN => n5399);
   U7535 : AOI221_X1 port map( B1 => n7129, B2 => n6795, C1 => n7126, C2 => 
                           n6819, A => n5407, ZN => n5404);
   U7536 : OAI22_X1 port map( A1 => n302, A2 => n7123, B1 => n270, B2 => n7120,
                           ZN => n5407);
   U7537 : AOI221_X1 port map( B1 => n7177, B2 => n6604, C1 => n7174, C2 => 
                           n6628, A => n5380, ZN => n5377);
   U7538 : OAI22_X1 port map( A1 => n813, A2 => n7171, B1 => n781, B2 => n7168,
                           ZN => n5380);
   U7539 : AOI221_X1 port map( B1 => n7129, B2 => n6796, C1 => n7126, C2 => 
                           n6820, A => n5388, ZN => n5385);
   U7540 : OAI22_X1 port map( A1 => n301, A2 => n7123, B1 => n269, B2 => n7120,
                           ZN => n5388);
   U7541 : AOI221_X1 port map( B1 => n7177, B2 => n6605, C1 => n7174, C2 => 
                           n6629, A => n5361, ZN => n5358);
   U7542 : OAI22_X1 port map( A1 => n812, A2 => n7171, B1 => n780, B2 => n7168,
                           ZN => n5361);
   U7543 : AOI221_X1 port map( B1 => n7129, B2 => n6797, C1 => n7126, C2 => 
                           n6821, A => n5369, ZN => n5366);
   U7544 : OAI22_X1 port map( A1 => n300, A2 => n7123, B1 => n268, B2 => n7120,
                           ZN => n5369);
   U7545 : AOI221_X1 port map( B1 => n7177, B2 => n6606, C1 => n7174, C2 => 
                           n6630, A => n5342, ZN => n5339);
   U7546 : OAI22_X1 port map( A1 => n811, A2 => n7171, B1 => n779, B2 => n7168,
                           ZN => n5342);
   U7547 : AOI221_X1 port map( B1 => n7129, B2 => n6798, C1 => n7126, C2 => 
                           n6822, A => n5350, ZN => n5347);
   U7548 : OAI22_X1 port map( A1 => n299, A2 => n7123, B1 => n267, B2 => n7120,
                           ZN => n5350);
   U7549 : AOI221_X1 port map( B1 => n7177, B2 => n6607, C1 => n7174, C2 => 
                           n6631, A => n5323, ZN => n5320);
   U7550 : OAI22_X1 port map( A1 => n810, A2 => n7171, B1 => n778, B2 => n7168,
                           ZN => n5323);
   U7551 : AOI221_X1 port map( B1 => n7129, B2 => n6799, C1 => n7126, C2 => 
                           n6823, A => n5331, ZN => n5328);
   U7552 : OAI22_X1 port map( A1 => n298, A2 => n7123, B1 => n266, B2 => n7120,
                           ZN => n5331);
   U7553 : AOI221_X1 port map( B1 => n7177, B2 => n6608, C1 => n7174, C2 => 
                           n6632, A => n5304, ZN => n5301);
   U7554 : OAI22_X1 port map( A1 => n809, A2 => n7171, B1 => n777, B2 => n7168,
                           ZN => n5304);
   U7555 : AOI221_X1 port map( B1 => n7129, B2 => n6800, C1 => n7126, C2 => 
                           n6824, A => n5312, ZN => n5309);
   U7556 : OAI22_X1 port map( A1 => n297, A2 => n7123, B1 => n265, B2 => n7120,
                           ZN => n5312);
   U7557 : AOI221_X1 port map( B1 => n7178, B2 => n6609, C1 => n7175, C2 => 
                           n6633, A => n5285, ZN => n5282);
   U7558 : OAI22_X1 port map( A1 => n808, A2 => n7172, B1 => n776, B2 => n7169,
                           ZN => n5285);
   U7559 : AOI221_X1 port map( B1 => n7130, B2 => n6801, C1 => n7127, C2 => 
                           n6825, A => n5293, ZN => n5290);
   U7560 : OAI22_X1 port map( A1 => n296, A2 => n7124, B1 => n264, B2 => n7121,
                           ZN => n5293);
   U7561 : AOI221_X1 port map( B1 => n7178, B2 => n6610, C1 => n7175, C2 => 
                           n6634, A => n5266, ZN => n5263);
   U7562 : OAI22_X1 port map( A1 => n807, A2 => n7172, B1 => n775, B2 => n7169,
                           ZN => n5266);
   U7563 : AOI221_X1 port map( B1 => n7130, B2 => n6802, C1 => n7127, C2 => 
                           n6826, A => n5274, ZN => n5271);
   U7564 : OAI22_X1 port map( A1 => n295, A2 => n7124, B1 => n263, B2 => n7121,
                           ZN => n5274);
   U7565 : AOI221_X1 port map( B1 => n7178, B2 => n6611, C1 => n7175, C2 => 
                           n6635, A => n5247, ZN => n5244);
   U7566 : OAI22_X1 port map( A1 => n806, A2 => n7172, B1 => n774, B2 => n7169,
                           ZN => n5247);
   U7567 : AOI221_X1 port map( B1 => n7130, B2 => n6803, C1 => n7127, C2 => 
                           n6827, A => n5255, ZN => n5252);
   U7568 : OAI22_X1 port map( A1 => n294, A2 => n7124, B1 => n262, B2 => n7121,
                           ZN => n5255);
   U7569 : AOI221_X1 port map( B1 => n7178, B2 => n6612, C1 => n7175, C2 => 
                           n6636, A => n5228, ZN => n5225);
   U7570 : OAI22_X1 port map( A1 => n805, A2 => n7172, B1 => n773, B2 => n7169,
                           ZN => n5228);
   U7571 : AOI221_X1 port map( B1 => n7130, B2 => n6804, C1 => n7127, C2 => 
                           n6828, A => n5236, ZN => n5233);
   U7572 : OAI22_X1 port map( A1 => n293, A2 => n7124, B1 => n261, B2 => n7121,
                           ZN => n5236);
   U7573 : AOI221_X1 port map( B1 => n7178, B2 => n6613, C1 => n7175, C2 => 
                           n6637, A => n5209, ZN => n5206);
   U7574 : OAI22_X1 port map( A1 => n804, A2 => n7172, B1 => n772, B2 => n7169,
                           ZN => n5209);
   U7575 : AOI221_X1 port map( B1 => n7130, B2 => n6805, C1 => n7127, C2 => 
                           n6829, A => n5217, ZN => n5214);
   U7576 : OAI22_X1 port map( A1 => n292, A2 => n7124, B1 => n260, B2 => n7121,
                           ZN => n5217);
   U7577 : AOI221_X1 port map( B1 => n7178, B2 => n6614, C1 => n7175, C2 => 
                           n6638, A => n5190, ZN => n5187);
   U7578 : OAI22_X1 port map( A1 => n803, A2 => n7172, B1 => n771, B2 => n7169,
                           ZN => n5190);
   U7579 : AOI221_X1 port map( B1 => n7130, B2 => n6806, C1 => n7127, C2 => 
                           n6830, A => n5198, ZN => n5195);
   U7580 : OAI22_X1 port map( A1 => n291, A2 => n7124, B1 => n259, B2 => n7121,
                           ZN => n5198);
   U7581 : AOI221_X1 port map( B1 => n7178, B2 => n6615, C1 => n7175, C2 => 
                           n6639, A => n5171, ZN => n5168);
   U7582 : OAI22_X1 port map( A1 => n802, A2 => n7172, B1 => n770, B2 => n7169,
                           ZN => n5171);
   U7583 : AOI221_X1 port map( B1 => n7130, B2 => n6807, C1 => n7127, C2 => 
                           n6831, A => n5179, ZN => n5176);
   U7584 : OAI22_X1 port map( A1 => n290, A2 => n7124, B1 => n258, B2 => n7121,
                           ZN => n5179);
   U7585 : AOI221_X1 port map( B1 => n7178, B2 => n6616, C1 => n7175, C2 => 
                           n6640, A => n5126, ZN => n5117);
   U7586 : OAI22_X1 port map( A1 => n801, A2 => n7172, B1 => n769, B2 => n7169,
                           ZN => n5126);
   U7587 : AOI221_X1 port map( B1 => n7130, B2 => n6808, C1 => n7127, C2 => 
                           n6832, A => n5150, ZN => n5141);
   U7588 : OAI22_X1 port map( A1 => n289, A2 => n7124, B1 => n257, B2 => n7121,
                           ZN => n5150);
   U7589 : AOI221_X1 port map( B1 => n7050, B2 => n6465, C1 => n7047, C2 => 
                           n6473, A => n6406, ZN => n6389);
   U7590 : OAI22_X1 port map( A1 => n576, A2 => n7044, B1 => n544, B2 => n7041,
                           ZN => n6406);
   U7591 : AOI221_X1 port map( B1 => n7002, B2 => n6529, C1 => n6999, C2 => 
                           n6537, A => n6416, ZN => n6407);
   U7592 : OAI22_X1 port map( A1 => n64, A2 => n6996, B1 => n32, B2 => n6993, 
                           ZN => n6416);
   U7593 : AOI221_X1 port map( B1 => n7050, B2 => n6466, C1 => n7047, C2 => 
                           n6474, A => n6377, ZN => n6370);
   U7594 : OAI22_X1 port map( A1 => n575, A2 => n7044, B1 => n543, B2 => n7041,
                           ZN => n6377);
   U7595 : AOI221_X1 port map( B1 => n7002, B2 => n6530, C1 => n6999, C2 => 
                           n6538, A => n6385, ZN => n6378);
   U7596 : OAI22_X1 port map( A1 => n63, A2 => n6996, B1 => n31, B2 => n6993, 
                           ZN => n6385);
   U7597 : AOI221_X1 port map( B1 => n7050, B2 => n6467, C1 => n7047, C2 => 
                           n6475, A => n6358, ZN => n6351);
   U7598 : OAI22_X1 port map( A1 => n574, A2 => n7044, B1 => n542, B2 => n7041,
                           ZN => n6358);
   U7599 : AOI221_X1 port map( B1 => n7002, B2 => n6531, C1 => n6999, C2 => 
                           n6539, A => n6366, ZN => n6359);
   U7600 : OAI22_X1 port map( A1 => n62, A2 => n6996, B1 => n30, B2 => n6993, 
                           ZN => n6366);
   U7601 : AOI221_X1 port map( B1 => n7050, B2 => n6468, C1 => n7047, C2 => 
                           n6476, A => n6339, ZN => n6332);
   U7602 : OAI22_X1 port map( A1 => n573, A2 => n7044, B1 => n541, B2 => n7041,
                           ZN => n6339);
   U7603 : AOI221_X1 port map( B1 => n7002, B2 => n6532, C1 => n6999, C2 => 
                           n6540, A => n6347, ZN => n6340);
   U7604 : OAI22_X1 port map( A1 => n61, A2 => n6996, B1 => n29, B2 => n6993, 
                           ZN => n6347);
   U7605 : AOI221_X1 port map( B1 => n7050, B2 => n6469, C1 => n7047, C2 => 
                           n6477, A => n6320, ZN => n6313);
   U7606 : OAI22_X1 port map( A1 => n572, A2 => n7044, B1 => n540, B2 => n7041,
                           ZN => n6320);
   U7607 : AOI221_X1 port map( B1 => n7002, B2 => n6533, C1 => n6999, C2 => 
                           n6541, A => n6328, ZN => n6321);
   U7608 : OAI22_X1 port map( A1 => n60, A2 => n6996, B1 => n28, B2 => n6993, 
                           ZN => n6328);
   U7609 : AOI221_X1 port map( B1 => n7050, B2 => n6470, C1 => n7047, C2 => 
                           n6478, A => n6301, ZN => n6294);
   U7610 : OAI22_X1 port map( A1 => n571, A2 => n7044, B1 => n539, B2 => n7041,
                           ZN => n6301);
   U7611 : AOI221_X1 port map( B1 => n7002, B2 => n6534, C1 => n6999, C2 => 
                           n6542, A => n6309, ZN => n6302);
   U7612 : OAI22_X1 port map( A1 => n59, A2 => n6996, B1 => n27, B2 => n6993, 
                           ZN => n6309);
   U7613 : AOI221_X1 port map( B1 => n7050, B2 => n6471, C1 => n7047, C2 => 
                           n6479, A => n6282, ZN => n6275);
   U7614 : OAI22_X1 port map( A1 => n570, A2 => n7044, B1 => n538, B2 => n7041,
                           ZN => n6282);
   U7615 : AOI221_X1 port map( B1 => n7002, B2 => n6535, C1 => n6999, C2 => 
                           n6543, A => n6290, ZN => n6283);
   U7616 : OAI22_X1 port map( A1 => n58, A2 => n6996, B1 => n26, B2 => n6993, 
                           ZN => n6290);
   U7617 : AOI221_X1 port map( B1 => n7050, B2 => n6472, C1 => n7047, C2 => 
                           n6480, A => n6263, ZN => n6256);
   U7618 : OAI22_X1 port map( A1 => n569, A2 => n7044, B1 => n537, B2 => n7041,
                           ZN => n6263);
   U7619 : AOI221_X1 port map( B1 => n7002, B2 => n6536, C1 => n6999, C2 => 
                           n6544, A => n6271, ZN => n6264);
   U7620 : OAI22_X1 port map( A1 => n57, A2 => n6996, B1 => n25, B2 => n6993, 
                           ZN => n6271);
   U7621 : AOI221_X1 port map( B1 => n7050, B2 => n6689, C1 => n7047, C2 => 
                           n6713, A => n6244, ZN => n6237);
   U7622 : OAI22_X1 port map( A1 => n568, A2 => n7044, B1 => n536, B2 => n7041,
                           ZN => n6244);
   U7623 : AOI221_X1 port map( B1 => n7002, B2 => n6881, C1 => n6999, C2 => 
                           n6905, A => n6252, ZN => n6245);
   U7624 : OAI22_X1 port map( A1 => n56, A2 => n6996, B1 => n24, B2 => n6993, 
                           ZN => n6252);
   U7625 : AOI221_X1 port map( B1 => n7050, B2 => n6690, C1 => n7047, C2 => 
                           n6714, A => n6225, ZN => n6218);
   U7626 : OAI22_X1 port map( A1 => n567, A2 => n7044, B1 => n535, B2 => n7041,
                           ZN => n6225);
   U7627 : AOI221_X1 port map( B1 => n7002, B2 => n6882, C1 => n6999, C2 => 
                           n6906, A => n6233, ZN => n6226);
   U7628 : OAI22_X1 port map( A1 => n55, A2 => n6996, B1 => n23, B2 => n6993, 
                           ZN => n6233);
   U7629 : AOI221_X1 port map( B1 => n7050, B2 => n6691, C1 => n7047, C2 => 
                           n6715, A => n6206, ZN => n6199);
   U7630 : OAI22_X1 port map( A1 => n566, A2 => n7044, B1 => n534, B2 => n7041,
                           ZN => n6206);
   U7631 : AOI221_X1 port map( B1 => n7002, B2 => n6883, C1 => n6999, C2 => 
                           n6907, A => n6214, ZN => n6207);
   U7632 : OAI22_X1 port map( A1 => n54, A2 => n6996, B1 => n22, B2 => n6993, 
                           ZN => n6214);
   U7633 : AOI221_X1 port map( B1 => n7050, B2 => n6692, C1 => n7047, C2 => 
                           n6716, A => n6187, ZN => n6180);
   U7634 : OAI22_X1 port map( A1 => n565, A2 => n7044, B1 => n533, B2 => n7041,
                           ZN => n6187);
   U7635 : AOI221_X1 port map( B1 => n7002, B2 => n6884, C1 => n6999, C2 => 
                           n6908, A => n6195, ZN => n6188);
   U7636 : OAI22_X1 port map( A1 => n53, A2 => n6996, B1 => n21, B2 => n6993, 
                           ZN => n6195);
   U7637 : AOI221_X1 port map( B1 => n7051, B2 => n6693, C1 => n7048, C2 => 
                           n6717, A => n6168, ZN => n6161);
   U7638 : OAI22_X1 port map( A1 => n564, A2 => n7045, B1 => n532, B2 => n7042,
                           ZN => n6168);
   U7639 : AOI221_X1 port map( B1 => n7003, B2 => n6885, C1 => n7000, C2 => 
                           n6909, A => n6176, ZN => n6169);
   U7640 : OAI22_X1 port map( A1 => n52, A2 => n6997, B1 => n20, B2 => n6994, 
                           ZN => n6176);
   U7641 : AOI221_X1 port map( B1 => n7051, B2 => n6694, C1 => n7048, C2 => 
                           n6718, A => n6149, ZN => n6142);
   U7642 : OAI22_X1 port map( A1 => n563, A2 => n7045, B1 => n531, B2 => n7042,
                           ZN => n6149);
   U7643 : AOI221_X1 port map( B1 => n7003, B2 => n6886, C1 => n7000, C2 => 
                           n6910, A => n6157, ZN => n6150);
   U7644 : OAI22_X1 port map( A1 => n51, A2 => n6997, B1 => n19, B2 => n6994, 
                           ZN => n6157);
   U7645 : AOI221_X1 port map( B1 => n7051, B2 => n6695, C1 => n7048, C2 => 
                           n6719, A => n6130, ZN => n6123);
   U7646 : OAI22_X1 port map( A1 => n562, A2 => n7045, B1 => n530, B2 => n7042,
                           ZN => n6130);
   U7647 : AOI221_X1 port map( B1 => n7003, B2 => n6887, C1 => n7000, C2 => 
                           n6911, A => n6138, ZN => n6131);
   U7648 : OAI22_X1 port map( A1 => n50, A2 => n6997, B1 => n18, B2 => n6994, 
                           ZN => n6138);
   U7649 : AOI221_X1 port map( B1 => n7051, B2 => n6696, C1 => n7048, C2 => 
                           n6720, A => n6111, ZN => n6104);
   U7650 : OAI22_X1 port map( A1 => n561, A2 => n7045, B1 => n529, B2 => n7042,
                           ZN => n6111);
   U7651 : AOI221_X1 port map( B1 => n7003, B2 => n6888, C1 => n7000, C2 => 
                           n6912, A => n6119, ZN => n6112);
   U7652 : OAI22_X1 port map( A1 => n49, A2 => n6997, B1 => n17, B2 => n6994, 
                           ZN => n6119);
   U7653 : AOI221_X1 port map( B1 => n7051, B2 => n6697, C1 => n7048, C2 => 
                           n6721, A => n6092, ZN => n6085);
   U7654 : OAI22_X1 port map( A1 => n560, A2 => n7045, B1 => n528, B2 => n7042,
                           ZN => n6092);
   U7655 : AOI221_X1 port map( B1 => n7003, B2 => n6889, C1 => n7000, C2 => 
                           n6913, A => n6100, ZN => n6093);
   U7656 : OAI22_X1 port map( A1 => n48, A2 => n6997, B1 => n16, B2 => n6994, 
                           ZN => n6100);
   U7657 : AOI221_X1 port map( B1 => n7051, B2 => n6698, C1 => n7048, C2 => 
                           n6722, A => n6073, ZN => n6066);
   U7658 : OAI22_X1 port map( A1 => n559, A2 => n7045, B1 => n527, B2 => n7042,
                           ZN => n6073);
   U7659 : AOI221_X1 port map( B1 => n7003, B2 => n6890, C1 => n7000, C2 => 
                           n6914, A => n6081, ZN => n6074);
   U7660 : OAI22_X1 port map( A1 => n47, A2 => n6997, B1 => n15, B2 => n6994, 
                           ZN => n6081);
   U7661 : AOI221_X1 port map( B1 => n7051, B2 => n6699, C1 => n7048, C2 => 
                           n6723, A => n6054, ZN => n6047);
   U7662 : OAI22_X1 port map( A1 => n558, A2 => n7045, B1 => n526, B2 => n7042,
                           ZN => n6054);
   U7663 : AOI221_X1 port map( B1 => n7003, B2 => n6891, C1 => n7000, C2 => 
                           n6915, A => n6062, ZN => n6055);
   U7664 : OAI22_X1 port map( A1 => n46, A2 => n6997, B1 => n14, B2 => n6994, 
                           ZN => n6062);
   U7665 : AOI221_X1 port map( B1 => n7051, B2 => n6700, C1 => n7048, C2 => 
                           n6724, A => n6035, ZN => n6028);
   U7666 : OAI22_X1 port map( A1 => n557, A2 => n7045, B1 => n525, B2 => n7042,
                           ZN => n6035);
   U7667 : AOI221_X1 port map( B1 => n7003, B2 => n6892, C1 => n7000, C2 => 
                           n6916, A => n6043, ZN => n6036);
   U7668 : OAI22_X1 port map( A1 => n45, A2 => n6997, B1 => n13, B2 => n6994, 
                           ZN => n6043);
   U7669 : AOI221_X1 port map( B1 => n7051, B2 => n6701, C1 => n7048, C2 => 
                           n6725, A => n6016, ZN => n6009);
   U7670 : OAI22_X1 port map( A1 => n556, A2 => n7045, B1 => n524, B2 => n7042,
                           ZN => n6016);
   U7671 : AOI221_X1 port map( B1 => n7003, B2 => n6893, C1 => n7000, C2 => 
                           n6917, A => n6024, ZN => n6017);
   U7672 : OAI22_X1 port map( A1 => n44, A2 => n6997, B1 => n12, B2 => n6994, 
                           ZN => n6024);
   U7673 : AOI221_X1 port map( B1 => n7051, B2 => n6702, C1 => n7048, C2 => 
                           n6726, A => n5997, ZN => n5990);
   U7674 : OAI22_X1 port map( A1 => n555, A2 => n7045, B1 => n523, B2 => n7042,
                           ZN => n5997);
   U7675 : AOI221_X1 port map( B1 => n7003, B2 => n6894, C1 => n7000, C2 => 
                           n6918, A => n6005, ZN => n5998);
   U7676 : OAI22_X1 port map( A1 => n43, A2 => n6997, B1 => n11, B2 => n6994, 
                           ZN => n6005);
   U7677 : AOI221_X1 port map( B1 => n7051, B2 => n6703, C1 => n7048, C2 => 
                           n6727, A => n5978, ZN => n5971);
   U7678 : OAI22_X1 port map( A1 => n554, A2 => n7045, B1 => n522, B2 => n7042,
                           ZN => n5978);
   U7679 : AOI221_X1 port map( B1 => n7003, B2 => n6895, C1 => n7000, C2 => 
                           n6919, A => n5986, ZN => n5979);
   U7680 : OAI22_X1 port map( A1 => n42, A2 => n6997, B1 => n10, B2 => n6994, 
                           ZN => n5986);
   U7681 : AOI221_X1 port map( B1 => n7051, B2 => n6704, C1 => n7048, C2 => 
                           n6728, A => n5959, ZN => n5952);
   U7682 : OAI22_X1 port map( A1 => n553, A2 => n7045, B1 => n521, B2 => n7042,
                           ZN => n5959);
   U7683 : AOI221_X1 port map( B1 => n7003, B2 => n6896, C1 => n7000, C2 => 
                           n6920, A => n5967, ZN => n5960);
   U7684 : OAI22_X1 port map( A1 => n41, A2 => n6997, B1 => n9, B2 => n6994, ZN
                           => n5967);
   U7685 : AOI221_X1 port map( B1 => n7052, B2 => n6705, C1 => n7049, C2 => 
                           n6729, A => n5940, ZN => n5933);
   U7686 : OAI22_X1 port map( A1 => n552, A2 => n7046, B1 => n520, B2 => n7043,
                           ZN => n5940);
   U7687 : AOI221_X1 port map( B1 => n7004, B2 => n6897, C1 => n7001, C2 => 
                           n6921, A => n5948, ZN => n5941);
   U7688 : OAI22_X1 port map( A1 => n40, A2 => n6998, B1 => n8, B2 => n6995, ZN
                           => n5948);
   U7689 : AOI221_X1 port map( B1 => n7052, B2 => n6706, C1 => n7049, C2 => 
                           n6730, A => n5921, ZN => n5914);
   U7690 : OAI22_X1 port map( A1 => n551, A2 => n7046, B1 => n519, B2 => n7043,
                           ZN => n5921);
   U7691 : AOI221_X1 port map( B1 => n7004, B2 => n6898, C1 => n7001, C2 => 
                           n6922, A => n5929, ZN => n5922);
   U7692 : OAI22_X1 port map( A1 => n39, A2 => n6998, B1 => n7, B2 => n6995, ZN
                           => n5929);
   U7693 : AOI221_X1 port map( B1 => n7052, B2 => n6707, C1 => n7049, C2 => 
                           n6731, A => n5902, ZN => n5895);
   U7694 : OAI22_X1 port map( A1 => n550, A2 => n7046, B1 => n518, B2 => n7043,
                           ZN => n5902);
   U7695 : AOI221_X1 port map( B1 => n7004, B2 => n6899, C1 => n7001, C2 => 
                           n6923, A => n5910, ZN => n5903);
   U7696 : OAI22_X1 port map( A1 => n38, A2 => n6998, B1 => n6, B2 => n6995, ZN
                           => n5910);
   U7697 : AOI221_X1 port map( B1 => n7052, B2 => n6708, C1 => n7049, C2 => 
                           n6732, A => n5883, ZN => n5876);
   U7698 : OAI22_X1 port map( A1 => n549, A2 => n7046, B1 => n517, B2 => n7043,
                           ZN => n5883);
   U7699 : AOI221_X1 port map( B1 => n7004, B2 => n6900, C1 => n7001, C2 => 
                           n6924, A => n5891, ZN => n5884);
   U7700 : OAI22_X1 port map( A1 => n37, A2 => n6998, B1 => n5, B2 => n6995, ZN
                           => n5891);
   U7701 : AOI221_X1 port map( B1 => n7052, B2 => n6709, C1 => n7049, C2 => 
                           n6733, A => n5864, ZN => n5857);
   U7702 : OAI22_X1 port map( A1 => n548, A2 => n7046, B1 => n516, B2 => n7043,
                           ZN => n5864);
   U7703 : AOI221_X1 port map( B1 => n7004, B2 => n6901, C1 => n7001, C2 => 
                           n6925, A => n5872, ZN => n5865);
   U7704 : OAI22_X1 port map( A1 => n36, A2 => n6998, B1 => n4, B2 => n6995, ZN
                           => n5872);
   U7705 : AOI221_X1 port map( B1 => n7052, B2 => n6710, C1 => n7049, C2 => 
                           n6734, A => n5845, ZN => n5838);
   U7706 : OAI22_X1 port map( A1 => n547, A2 => n7046, B1 => n515, B2 => n7043,
                           ZN => n5845);
   U7707 : AOI221_X1 port map( B1 => n7004, B2 => n6902, C1 => n7001, C2 => 
                           n6926, A => n5853, ZN => n5846);
   U7708 : OAI22_X1 port map( A1 => n35, A2 => n6998, B1 => n3, B2 => n6995, ZN
                           => n5853);
   U7709 : AOI221_X1 port map( B1 => n7052, B2 => n6711, C1 => n7049, C2 => 
                           n6735, A => n5826, ZN => n5819);
   U7710 : OAI22_X1 port map( A1 => n546, A2 => n7046, B1 => n514, B2 => n7043,
                           ZN => n5826);
   U7711 : AOI221_X1 port map( B1 => n7004, B2 => n6903, C1 => n7001, C2 => 
                           n6927, A => n5834, ZN => n5827);
   U7712 : OAI22_X1 port map( A1 => n34, A2 => n6998, B1 => n2, B2 => n6995, ZN
                           => n5834);
   U7713 : AOI221_X1 port map( B1 => n7052, B2 => n6712, C1 => n7049, C2 => 
                           n6736, A => n5789, ZN => n5768);
   U7714 : OAI22_X1 port map( A1 => n545, A2 => n7046, B1 => n513, B2 => n7043,
                           ZN => n5789);
   U7715 : AOI221_X1 port map( B1 => n7004, B2 => n6904, C1 => n7001, C2 => 
                           n6928, A => n5813, ZN => n5792);
   U7716 : OAI22_X1 port map( A1 => n33, A2 => n6998, B1 => n1, B2 => n6995, ZN
                           => n5813);
   U7717 : AOI221_X1 port map( B1 => n7152, B2 => n6465, C1 => n7149, C2 => 
                           n6473, A => n5753, ZN => n5736);
   U7718 : OAI22_X1 port map( A1 => n576, A2 => n7146, B1 => n544, B2 => n7143,
                           ZN => n5753);
   U7719 : AOI221_X1 port map( B1 => n7104, B2 => n6529, C1 => n7101, C2 => 
                           n6537, A => n5763, ZN => n5754);
   U7720 : OAI22_X1 port map( A1 => n64, A2 => n7098, B1 => n32, B2 => n7095, 
                           ZN => n5763);
   U7721 : AOI221_X1 port map( B1 => n7152, B2 => n6466, C1 => n7149, C2 => 
                           n6474, A => n5724, ZN => n5717);
   U7722 : OAI22_X1 port map( A1 => n575, A2 => n7146, B1 => n543, B2 => n7143,
                           ZN => n5724);
   U7723 : AOI221_X1 port map( B1 => n7104, B2 => n6530, C1 => n7101, C2 => 
                           n6538, A => n5732, ZN => n5725);
   U7724 : OAI22_X1 port map( A1 => n63, A2 => n7098, B1 => n31, B2 => n7095, 
                           ZN => n5732);
   U7725 : AOI221_X1 port map( B1 => n7152, B2 => n6467, C1 => n7149, C2 => 
                           n6475, A => n5705, ZN => n5698);
   U7726 : OAI22_X1 port map( A1 => n574, A2 => n7146, B1 => n542, B2 => n7143,
                           ZN => n5705);
   U7727 : AOI221_X1 port map( B1 => n7104, B2 => n6531, C1 => n7101, C2 => 
                           n6539, A => n5713, ZN => n5706);
   U7728 : OAI22_X1 port map( A1 => n62, A2 => n7098, B1 => n30, B2 => n7095, 
                           ZN => n5713);
   U7729 : AOI221_X1 port map( B1 => n7152, B2 => n6468, C1 => n7149, C2 => 
                           n6476, A => n5686, ZN => n5679);
   U7730 : OAI22_X1 port map( A1 => n573, A2 => n7146, B1 => n541, B2 => n7143,
                           ZN => n5686);
   U7731 : AOI221_X1 port map( B1 => n7104, B2 => n6532, C1 => n7101, C2 => 
                           n6540, A => n5694, ZN => n5687);
   U7732 : OAI22_X1 port map( A1 => n61, A2 => n7098, B1 => n29, B2 => n7095, 
                           ZN => n5694);
   U7733 : AOI221_X1 port map( B1 => n7152, B2 => n6469, C1 => n7149, C2 => 
                           n6477, A => n5667, ZN => n5660);
   U7734 : OAI22_X1 port map( A1 => n572, A2 => n7146, B1 => n540, B2 => n7143,
                           ZN => n5667);
   U7735 : AOI221_X1 port map( B1 => n7104, B2 => n6533, C1 => n7101, C2 => 
                           n6541, A => n5675, ZN => n5668);
   U7736 : OAI22_X1 port map( A1 => n60, A2 => n7098, B1 => n28, B2 => n7095, 
                           ZN => n5675);
   U7737 : AOI221_X1 port map( B1 => n7152, B2 => n6470, C1 => n7149, C2 => 
                           n6478, A => n5648, ZN => n5641);
   U7738 : OAI22_X1 port map( A1 => n571, A2 => n7146, B1 => n539, B2 => n7143,
                           ZN => n5648);
   U7739 : AOI221_X1 port map( B1 => n7104, B2 => n6534, C1 => n7101, C2 => 
                           n6542, A => n5656, ZN => n5649);
   U7740 : OAI22_X1 port map( A1 => n59, A2 => n7098, B1 => n27, B2 => n7095, 
                           ZN => n5656);
   U7741 : AOI221_X1 port map( B1 => n7152, B2 => n6471, C1 => n7149, C2 => 
                           n6479, A => n5629, ZN => n5622);
   U7742 : OAI22_X1 port map( A1 => n570, A2 => n7146, B1 => n538, B2 => n7143,
                           ZN => n5629);
   U7743 : AOI221_X1 port map( B1 => n7104, B2 => n6535, C1 => n7101, C2 => 
                           n6543, A => n5637, ZN => n5630);
   U7744 : OAI22_X1 port map( A1 => n58, A2 => n7098, B1 => n26, B2 => n7095, 
                           ZN => n5637);
   U7745 : AOI221_X1 port map( B1 => n7152, B2 => n6472, C1 => n7149, C2 => 
                           n6480, A => n5610, ZN => n5603);
   U7746 : OAI22_X1 port map( A1 => n569, A2 => n7146, B1 => n537, B2 => n7143,
                           ZN => n5610);
   U7747 : AOI221_X1 port map( B1 => n7104, B2 => n6536, C1 => n7101, C2 => 
                           n6544, A => n5618, ZN => n5611);
   U7748 : OAI22_X1 port map( A1 => n57, A2 => n7098, B1 => n25, B2 => n7095, 
                           ZN => n5618);
   U7749 : AOI221_X1 port map( B1 => n7152, B2 => n6689, C1 => n7149, C2 => 
                           n6713, A => n5591, ZN => n5584);
   U7750 : OAI22_X1 port map( A1 => n568, A2 => n7146, B1 => n536, B2 => n7143,
                           ZN => n5591);
   U7751 : AOI221_X1 port map( B1 => n7104, B2 => n6881, C1 => n7101, C2 => 
                           n6905, A => n5599, ZN => n5592);
   U7752 : OAI22_X1 port map( A1 => n56, A2 => n7098, B1 => n24, B2 => n7095, 
                           ZN => n5599);
   U7753 : AOI221_X1 port map( B1 => n7152, B2 => n6690, C1 => n7149, C2 => 
                           n6714, A => n5572, ZN => n5565);
   U7754 : OAI22_X1 port map( A1 => n567, A2 => n7146, B1 => n535, B2 => n7143,
                           ZN => n5572);
   U7755 : AOI221_X1 port map( B1 => n7104, B2 => n6882, C1 => n7101, C2 => 
                           n6906, A => n5580, ZN => n5573);
   U7756 : OAI22_X1 port map( A1 => n55, A2 => n7098, B1 => n23, B2 => n7095, 
                           ZN => n5580);
   U7757 : AOI221_X1 port map( B1 => n7152, B2 => n6691, C1 => n7149, C2 => 
                           n6715, A => n5553, ZN => n5546);
   U7758 : OAI22_X1 port map( A1 => n566, A2 => n7146, B1 => n534, B2 => n7143,
                           ZN => n5553);
   U7759 : AOI221_X1 port map( B1 => n7104, B2 => n6883, C1 => n7101, C2 => 
                           n6907, A => n5561, ZN => n5554);
   U7760 : OAI22_X1 port map( A1 => n54, A2 => n7098, B1 => n22, B2 => n7095, 
                           ZN => n5561);
   U7761 : AOI221_X1 port map( B1 => n7152, B2 => n6692, C1 => n7149, C2 => 
                           n6716, A => n5534, ZN => n5527);
   U7762 : OAI22_X1 port map( A1 => n565, A2 => n7146, B1 => n533, B2 => n7143,
                           ZN => n5534);
   U7763 : AOI221_X1 port map( B1 => n7104, B2 => n6884, C1 => n7101, C2 => 
                           n6908, A => n5542, ZN => n5535);
   U7764 : OAI22_X1 port map( A1 => n53, A2 => n7098, B1 => n21, B2 => n7095, 
                           ZN => n5542);
   U7765 : AOI221_X1 port map( B1 => n7153, B2 => n6693, C1 => n7150, C2 => 
                           n6717, A => n5515, ZN => n5508);
   U7766 : OAI22_X1 port map( A1 => n564, A2 => n7147, B1 => n532, B2 => n7144,
                           ZN => n5515);
   U7767 : AOI221_X1 port map( B1 => n7105, B2 => n6885, C1 => n7102, C2 => 
                           n6909, A => n5523, ZN => n5516);
   U7768 : OAI22_X1 port map( A1 => n52, A2 => n7099, B1 => n20, B2 => n7096, 
                           ZN => n5523);
   U7769 : AOI221_X1 port map( B1 => n7153, B2 => n6694, C1 => n7150, C2 => 
                           n6718, A => n5496, ZN => n5489);
   U7770 : OAI22_X1 port map( A1 => n563, A2 => n7147, B1 => n531, B2 => n7144,
                           ZN => n5496);
   U7771 : AOI221_X1 port map( B1 => n7105, B2 => n6886, C1 => n7102, C2 => 
                           n6910, A => n5504, ZN => n5497);
   U7772 : OAI22_X1 port map( A1 => n51, A2 => n7099, B1 => n19, B2 => n7096, 
                           ZN => n5504);
   U7773 : AOI221_X1 port map( B1 => n7153, B2 => n6695, C1 => n7150, C2 => 
                           n6719, A => n5477, ZN => n5470);
   U7774 : OAI22_X1 port map( A1 => n562, A2 => n7147, B1 => n530, B2 => n7144,
                           ZN => n5477);
   U7775 : AOI221_X1 port map( B1 => n7105, B2 => n6887, C1 => n7102, C2 => 
                           n6911, A => n5485, ZN => n5478);
   U7776 : OAI22_X1 port map( A1 => n50, A2 => n7099, B1 => n18, B2 => n7096, 
                           ZN => n5485);
   U7777 : AOI221_X1 port map( B1 => n7153, B2 => n6696, C1 => n7150, C2 => 
                           n6720, A => n5458, ZN => n5451);
   U7778 : OAI22_X1 port map( A1 => n561, A2 => n7147, B1 => n529, B2 => n7144,
                           ZN => n5458);
   U7779 : AOI221_X1 port map( B1 => n7105, B2 => n6888, C1 => n7102, C2 => 
                           n6912, A => n5466, ZN => n5459);
   U7780 : OAI22_X1 port map( A1 => n49, A2 => n7099, B1 => n17, B2 => n7096, 
                           ZN => n5466);
   U7781 : AOI221_X1 port map( B1 => n7153, B2 => n6697, C1 => n7150, C2 => 
                           n6721, A => n5439, ZN => n5432);
   U7782 : OAI22_X1 port map( A1 => n560, A2 => n7147, B1 => n528, B2 => n7144,
                           ZN => n5439);
   U7783 : AOI221_X1 port map( B1 => n7105, B2 => n6889, C1 => n7102, C2 => 
                           n6913, A => n5447, ZN => n5440);
   U7784 : OAI22_X1 port map( A1 => n48, A2 => n7099, B1 => n16, B2 => n7096, 
                           ZN => n5447);
   U7785 : AOI221_X1 port map( B1 => n7153, B2 => n6698, C1 => n7150, C2 => 
                           n6722, A => n5420, ZN => n5413);
   U7786 : OAI22_X1 port map( A1 => n559, A2 => n7147, B1 => n527, B2 => n7144,
                           ZN => n5420);
   U7787 : AOI221_X1 port map( B1 => n7105, B2 => n6890, C1 => n7102, C2 => 
                           n6914, A => n5428, ZN => n5421);
   U7788 : OAI22_X1 port map( A1 => n47, A2 => n7099, B1 => n15, B2 => n7096, 
                           ZN => n5428);
   U7789 : AOI221_X1 port map( B1 => n7153, B2 => n6699, C1 => n7150, C2 => 
                           n6723, A => n5401, ZN => n5394);
   U7790 : OAI22_X1 port map( A1 => n558, A2 => n7147, B1 => n526, B2 => n7144,
                           ZN => n5401);
   U7791 : AOI221_X1 port map( B1 => n7105, B2 => n6891, C1 => n7102, C2 => 
                           n6915, A => n5409, ZN => n5402);
   U7792 : OAI22_X1 port map( A1 => n46, A2 => n7099, B1 => n14, B2 => n7096, 
                           ZN => n5409);
   U7793 : AOI221_X1 port map( B1 => n7153, B2 => n6700, C1 => n7150, C2 => 
                           n6724, A => n5382, ZN => n5375);
   U7794 : OAI22_X1 port map( A1 => n557, A2 => n7147, B1 => n525, B2 => n7144,
                           ZN => n5382);
   U7795 : AOI221_X1 port map( B1 => n7105, B2 => n6892, C1 => n7102, C2 => 
                           n6916, A => n5390, ZN => n5383);
   U7796 : OAI22_X1 port map( A1 => n45, A2 => n7099, B1 => n13, B2 => n7096, 
                           ZN => n5390);
   U7797 : AOI221_X1 port map( B1 => n7153, B2 => n6701, C1 => n7150, C2 => 
                           n6725, A => n5363, ZN => n5356);
   U7798 : OAI22_X1 port map( A1 => n556, A2 => n7147, B1 => n524, B2 => n7144,
                           ZN => n5363);
   U7799 : AOI221_X1 port map( B1 => n7105, B2 => n6893, C1 => n7102, C2 => 
                           n6917, A => n5371, ZN => n5364);
   U7800 : OAI22_X1 port map( A1 => n44, A2 => n7099, B1 => n12, B2 => n7096, 
                           ZN => n5371);
   U7801 : AOI221_X1 port map( B1 => n7153, B2 => n6702, C1 => n7150, C2 => 
                           n6726, A => n5344, ZN => n5337);
   U7802 : OAI22_X1 port map( A1 => n555, A2 => n7147, B1 => n523, B2 => n7144,
                           ZN => n5344);
   U7803 : AOI221_X1 port map( B1 => n7105, B2 => n6894, C1 => n7102, C2 => 
                           n6918, A => n5352, ZN => n5345);
   U7804 : OAI22_X1 port map( A1 => n43, A2 => n7099, B1 => n11, B2 => n7096, 
                           ZN => n5352);
   U7805 : AOI221_X1 port map( B1 => n7153, B2 => n6703, C1 => n7150, C2 => 
                           n6727, A => n5325, ZN => n5318);
   U7806 : OAI22_X1 port map( A1 => n554, A2 => n7147, B1 => n522, B2 => n7144,
                           ZN => n5325);
   U7807 : AOI221_X1 port map( B1 => n7105, B2 => n6895, C1 => n7102, C2 => 
                           n6919, A => n5333, ZN => n5326);
   U7808 : OAI22_X1 port map( A1 => n42, A2 => n7099, B1 => n10, B2 => n7096, 
                           ZN => n5333);
   U7809 : AOI221_X1 port map( B1 => n7153, B2 => n6704, C1 => n7150, C2 => 
                           n6728, A => n5306, ZN => n5299);
   U7810 : OAI22_X1 port map( A1 => n553, A2 => n7147, B1 => n521, B2 => n7144,
                           ZN => n5306);
   U7811 : AOI221_X1 port map( B1 => n7105, B2 => n6896, C1 => n7102, C2 => 
                           n6920, A => n5314, ZN => n5307);
   U7812 : OAI22_X1 port map( A1 => n41, A2 => n7099, B1 => n9, B2 => n7096, ZN
                           => n5314);
   U7813 : AOI221_X1 port map( B1 => n7154, B2 => n6705, C1 => n7151, C2 => 
                           n6729, A => n5287, ZN => n5280);
   U7814 : OAI22_X1 port map( A1 => n552, A2 => n7148, B1 => n520, B2 => n7145,
                           ZN => n5287);
   U7815 : AOI221_X1 port map( B1 => n7106, B2 => n6897, C1 => n7103, C2 => 
                           n6921, A => n5295, ZN => n5288);
   U7816 : OAI22_X1 port map( A1 => n40, A2 => n7100, B1 => n8, B2 => n7097, ZN
                           => n5295);
   U7817 : AOI221_X1 port map( B1 => n7154, B2 => n6706, C1 => n7151, C2 => 
                           n6730, A => n5268, ZN => n5261);
   U7818 : OAI22_X1 port map( A1 => n551, A2 => n7148, B1 => n519, B2 => n7145,
                           ZN => n5268);
   U7819 : AOI221_X1 port map( B1 => n7106, B2 => n6898, C1 => n7103, C2 => 
                           n6922, A => n5276, ZN => n5269);
   U7820 : OAI22_X1 port map( A1 => n39, A2 => n7100, B1 => n7, B2 => n7097, ZN
                           => n5276);
   U7821 : AOI221_X1 port map( B1 => n7154, B2 => n6707, C1 => n7151, C2 => 
                           n6731, A => n5249, ZN => n5242);
   U7822 : OAI22_X1 port map( A1 => n550, A2 => n7148, B1 => n518, B2 => n7145,
                           ZN => n5249);
   U7823 : AOI221_X1 port map( B1 => n7106, B2 => n6899, C1 => n7103, C2 => 
                           n6923, A => n5257, ZN => n5250);
   U7824 : OAI22_X1 port map( A1 => n38, A2 => n7100, B1 => n6, B2 => n7097, ZN
                           => n5257);
   U7825 : AOI221_X1 port map( B1 => n7154, B2 => n6708, C1 => n7151, C2 => 
                           n6732, A => n5230, ZN => n5223);
   U7826 : OAI22_X1 port map( A1 => n549, A2 => n7148, B1 => n517, B2 => n7145,
                           ZN => n5230);
   U7827 : AOI221_X1 port map( B1 => n7106, B2 => n6900, C1 => n7103, C2 => 
                           n6924, A => n5238, ZN => n5231);
   U7828 : OAI22_X1 port map( A1 => n37, A2 => n7100, B1 => n5, B2 => n7097, ZN
                           => n5238);
   U7829 : AOI221_X1 port map( B1 => n7154, B2 => n6709, C1 => n7151, C2 => 
                           n6733, A => n5211, ZN => n5204);
   U7830 : OAI22_X1 port map( A1 => n548, A2 => n7148, B1 => n516, B2 => n7145,
                           ZN => n5211);
   U7831 : AOI221_X1 port map( B1 => n7106, B2 => n6901, C1 => n7103, C2 => 
                           n6925, A => n5219, ZN => n5212);
   U7832 : OAI22_X1 port map( A1 => n36, A2 => n7100, B1 => n4, B2 => n7097, ZN
                           => n5219);
   U7833 : AOI221_X1 port map( B1 => n7154, B2 => n6710, C1 => n7151, C2 => 
                           n6734, A => n5192, ZN => n5185);
   U7834 : OAI22_X1 port map( A1 => n547, A2 => n7148, B1 => n515, B2 => n7145,
                           ZN => n5192);
   U7835 : AOI221_X1 port map( B1 => n7106, B2 => n6902, C1 => n7103, C2 => 
                           n6926, A => n5200, ZN => n5193);
   U7836 : OAI22_X1 port map( A1 => n35, A2 => n7100, B1 => n3, B2 => n7097, ZN
                           => n5200);
   U7837 : AOI221_X1 port map( B1 => n7154, B2 => n6711, C1 => n7151, C2 => 
                           n6735, A => n5173, ZN => n5166);
   U7838 : OAI22_X1 port map( A1 => n546, A2 => n7148, B1 => n514, B2 => n7145,
                           ZN => n5173);
   U7839 : AOI221_X1 port map( B1 => n7106, B2 => n6903, C1 => n7103, C2 => 
                           n6927, A => n5181, ZN => n5174);
   U7840 : OAI22_X1 port map( A1 => n34, A2 => n7100, B1 => n2, B2 => n7097, ZN
                           => n5181);
   U7841 : AOI221_X1 port map( B1 => n7154, B2 => n6712, C1 => n7151, C2 => 
                           n6736, A => n5136, ZN => n5115);
   U7842 : OAI22_X1 port map( A1 => n545, A2 => n7148, B1 => n513, B2 => n7145,
                           ZN => n5136);
   U7843 : AOI221_X1 port map( B1 => n7106, B2 => n6904, C1 => n7103, C2 => 
                           n6928, A => n5160, ZN => n5139);
   U7844 : OAI22_X1 port map( A1 => n33, A2 => n7100, B1 => n1, B2 => n7097, ZN
                           => n5160);
   U7845 : OAI22_X1 port map( A1 => n7248, A2 => n7551, B1 => n5105, B2 => 
                           n4849, ZN => n2776);
   U7846 : OAI22_X1 port map( A1 => n7249, A2 => n7554, B1 => n5105, B2 => 
                           n4848, ZN => n2777);
   U7847 : OAI22_X1 port map( A1 => n7249, A2 => n7557, B1 => n5105, B2 => 
                           n4847, ZN => n2778);
   U7848 : OAI22_X1 port map( A1 => n7249, A2 => n7560, B1 => n5105, B2 => 
                           n4846, ZN => n2779);
   U7849 : OAI22_X1 port map( A1 => n7249, A2 => n7563, B1 => n5105, B2 => 
                           n4845, ZN => n2780);
   U7850 : OAI22_X1 port map( A1 => n7249, A2 => n7566, B1 => n5105, B2 => 
                           n4844, ZN => n2781);
   U7851 : OAI22_X1 port map( A1 => n7250, A2 => n7569, B1 => n5105, B2 => 
                           n4843, ZN => n2782);
   U7852 : OAI22_X1 port map( A1 => n7250, A2 => n7581, B1 => n5105, B2 => 
                           n4842, ZN => n2783);
   U7853 : OAI22_X1 port map( A1 => n7320, A2 => n7550, B1 => n5096, B2 => 
                           n4657, ZN => n3032);
   U7854 : OAI22_X1 port map( A1 => n7321, A2 => n7553, B1 => n5096, B2 => 
                           n4656, ZN => n3033);
   U7855 : OAI22_X1 port map( A1 => n7321, A2 => n7556, B1 => n5096, B2 => 
                           n4655, ZN => n3034);
   U7856 : OAI22_X1 port map( A1 => n7321, A2 => n7559, B1 => n5096, B2 => 
                           n4654, ZN => n3035);
   U7857 : OAI22_X1 port map( A1 => n7321, A2 => n7562, B1 => n5096, B2 => 
                           n4653, ZN => n3036);
   U7858 : OAI22_X1 port map( A1 => n7321, A2 => n7565, B1 => n5096, B2 => 
                           n4652, ZN => n3037);
   U7859 : OAI22_X1 port map( A1 => n7322, A2 => n7568, B1 => n5096, B2 => 
                           n4651, ZN => n3038);
   U7860 : OAI22_X1 port map( A1 => n7322, A2 => n7580, B1 => n5096, B2 => 
                           n4650, ZN => n3039);
   U7861 : OAI22_X1 port map( A1 => n7392, A2 => n7549, B1 => n5087, B2 => 
                           n4465, ZN => n3288);
   U7862 : OAI22_X1 port map( A1 => n7393, A2 => n7552, B1 => n5087, B2 => 
                           n4464, ZN => n3289);
   U7863 : OAI22_X1 port map( A1 => n7393, A2 => n7555, B1 => n5087, B2 => 
                           n4463, ZN => n3290);
   U7864 : OAI22_X1 port map( A1 => n7393, A2 => n7558, B1 => n5087, B2 => 
                           n4462, ZN => n3291);
   U7865 : OAI22_X1 port map( A1 => n7393, A2 => n7561, B1 => n5087, B2 => 
                           n4461, ZN => n3292);
   U7866 : OAI22_X1 port map( A1 => n7393, A2 => n7564, B1 => n5087, B2 => 
                           n4460, ZN => n3293);
   U7867 : OAI22_X1 port map( A1 => n7394, A2 => n7567, B1 => n5087, B2 => 
                           n4459, ZN => n3294);
   U7868 : OAI22_X1 port map( A1 => n7394, A2 => n7579, B1 => n5087, B2 => 
                           n4458, ZN => n3295);
   U7869 : OAI22_X1 port map( A1 => n7464, A2 => n7549, B1 => n5071, B2 => 
                           n4273, ZN => n3544);
   U7870 : OAI22_X1 port map( A1 => n7465, A2 => n7552, B1 => n5071, B2 => 
                           n4272, ZN => n3545);
   U7871 : OAI22_X1 port map( A1 => n7465, A2 => n7555, B1 => n5071, B2 => 
                           n4271, ZN => n3546);
   U7872 : OAI22_X1 port map( A1 => n7465, A2 => n7558, B1 => n5071, B2 => 
                           n4270, ZN => n3547);
   U7873 : OAI22_X1 port map( A1 => n7465, A2 => n7561, B1 => n5071, B2 => 
                           n4269, ZN => n3548);
   U7874 : OAI22_X1 port map( A1 => n7465, A2 => n7564, B1 => n5071, B2 => 
                           n4268, ZN => n3549);
   U7875 : OAI22_X1 port map( A1 => n7466, A2 => n7567, B1 => n5071, B2 => 
                           n4267, ZN => n3550);
   U7876 : OAI22_X1 port map( A1 => n7466, A2 => n7579, B1 => n5071, B2 => 
                           n4266, ZN => n3551);
   U7877 : OAI22_X1 port map( A1 => n7212, A2 => n7551, B1 => n968, B2 => n5109
                           , ZN => n2648);
   U7878 : OAI22_X1 port map( A1 => n7213, A2 => n7554, B1 => n967, B2 => n5109
                           , ZN => n2649);
   U7879 : OAI22_X1 port map( A1 => n7213, A2 => n7557, B1 => n966, B2 => n5109
                           , ZN => n2650);
   U7880 : OAI22_X1 port map( A1 => n7213, A2 => n7560, B1 => n965, B2 => n5109
                           , ZN => n2651);
   U7881 : OAI22_X1 port map( A1 => n7213, A2 => n7563, B1 => n964, B2 => n5109
                           , ZN => n2652);
   U7882 : OAI22_X1 port map( A1 => n7213, A2 => n7566, B1 => n963, B2 => n5109
                           , ZN => n2653);
   U7883 : OAI22_X1 port map( A1 => n7214, A2 => n7569, B1 => n962, B2 => n5109
                           , ZN => n2654);
   U7884 : OAI22_X1 port map( A1 => n7214, A2 => n7581, B1 => n961, B2 => n5109
                           , ZN => n2655);
   U7885 : OAI22_X1 port map( A1 => n7257, A2 => n7551, B1 => n808, B2 => n5104
                           , ZN => n2808);
   U7886 : OAI22_X1 port map( A1 => n7258, A2 => n7554, B1 => n807, B2 => n5104
                           , ZN => n2809);
   U7887 : OAI22_X1 port map( A1 => n7258, A2 => n7557, B1 => n806, B2 => n5104
                           , ZN => n2810);
   U7888 : OAI22_X1 port map( A1 => n7258, A2 => n7560, B1 => n805, B2 => n5104
                           , ZN => n2811);
   U7889 : OAI22_X1 port map( A1 => n7258, A2 => n7563, B1 => n804, B2 => n5104
                           , ZN => n2812);
   U7890 : OAI22_X1 port map( A1 => n7258, A2 => n7566, B1 => n803, B2 => n5104
                           , ZN => n2813);
   U7891 : OAI22_X1 port map( A1 => n7259, A2 => n7569, B1 => n802, B2 => n5104
                           , ZN => n2814);
   U7892 : OAI22_X1 port map( A1 => n7259, A2 => n7581, B1 => n801, B2 => n5104
                           , ZN => n2815);
   U7893 : OAI22_X1 port map( A1 => n7266, A2 => n7551, B1 => n776, B2 => n5102
                           , ZN => n2840);
   U7894 : OAI22_X1 port map( A1 => n7267, A2 => n7554, B1 => n775, B2 => n5102
                           , ZN => n2841);
   U7895 : OAI22_X1 port map( A1 => n7267, A2 => n7557, B1 => n774, B2 => n5102
                           , ZN => n2842);
   U7896 : OAI22_X1 port map( A1 => n7267, A2 => n7560, B1 => n773, B2 => n5102
                           , ZN => n2843);
   U7897 : OAI22_X1 port map( A1 => n7267, A2 => n7563, B1 => n772, B2 => n5102
                           , ZN => n2844);
   U7898 : OAI22_X1 port map( A1 => n7267, A2 => n7566, B1 => n771, B2 => n5102
                           , ZN => n2845);
   U7899 : OAI22_X1 port map( A1 => n7268, A2 => n7569, B1 => n770, B2 => n5102
                           , ZN => n2846);
   U7900 : OAI22_X1 port map( A1 => n7268, A2 => n7581, B1 => n769, B2 => n5102
                           , ZN => n2847);
   U7901 : OAI22_X1 port map( A1 => n7275, A2 => n7550, B1 => n744, B2 => n5101
                           , ZN => n2872);
   U7902 : OAI22_X1 port map( A1 => n7276, A2 => n7553, B1 => n743, B2 => n5101
                           , ZN => n2873);
   U7903 : OAI22_X1 port map( A1 => n7276, A2 => n7556, B1 => n742, B2 => n5101
                           , ZN => n2874);
   U7904 : OAI22_X1 port map( A1 => n7276, A2 => n7559, B1 => n741, B2 => n5101
                           , ZN => n2875);
   U7905 : OAI22_X1 port map( A1 => n7276, A2 => n7562, B1 => n740, B2 => n5101
                           , ZN => n2876);
   U7906 : OAI22_X1 port map( A1 => n7276, A2 => n7565, B1 => n739, B2 => n5101
                           , ZN => n2877);
   U7907 : OAI22_X1 port map( A1 => n7277, A2 => n7568, B1 => n738, B2 => n5101
                           , ZN => n2878);
   U7908 : OAI22_X1 port map( A1 => n7277, A2 => n7580, B1 => n737, B2 => n5101
                           , ZN => n2879);
   U7909 : OAI22_X1 port map( A1 => n7284, A2 => n7550, B1 => n712, B2 => n5100
                           , ZN => n2904);
   U7910 : OAI22_X1 port map( A1 => n7285, A2 => n7553, B1 => n711, B2 => n5100
                           , ZN => n2905);
   U7911 : OAI22_X1 port map( A1 => n7285, A2 => n7556, B1 => n710, B2 => n5100
                           , ZN => n2906);
   U7912 : OAI22_X1 port map( A1 => n7285, A2 => n7559, B1 => n709, B2 => n5100
                           , ZN => n2907);
   U7913 : OAI22_X1 port map( A1 => n7285, A2 => n7562, B1 => n708, B2 => n5100
                           , ZN => n2908);
   U7914 : OAI22_X1 port map( A1 => n7285, A2 => n7565, B1 => n707, B2 => n5100
                           , ZN => n2909);
   U7915 : OAI22_X1 port map( A1 => n7286, A2 => n7568, B1 => n706, B2 => n5100
                           , ZN => n2910);
   U7916 : OAI22_X1 port map( A1 => n7286, A2 => n7580, B1 => n705, B2 => n5100
                           , ZN => n2911);
   U7917 : OAI22_X1 port map( A1 => n7329, A2 => n7550, B1 => n552, B2 => n5095
                           , ZN => n3064);
   U7918 : OAI22_X1 port map( A1 => n7330, A2 => n7553, B1 => n551, B2 => n5095
                           , ZN => n3065);
   U7919 : OAI22_X1 port map( A1 => n7330, A2 => n7556, B1 => n550, B2 => n5095
                           , ZN => n3066);
   U7920 : OAI22_X1 port map( A1 => n7330, A2 => n7559, B1 => n549, B2 => n5095
                           , ZN => n3067);
   U7921 : OAI22_X1 port map( A1 => n7330, A2 => n7562, B1 => n548, B2 => n5095
                           , ZN => n3068);
   U7922 : OAI22_X1 port map( A1 => n7330, A2 => n7565, B1 => n547, B2 => n5095
                           , ZN => n3069);
   U7923 : OAI22_X1 port map( A1 => n7331, A2 => n7568, B1 => n546, B2 => n5095
                           , ZN => n3070);
   U7924 : OAI22_X1 port map( A1 => n7331, A2 => n7580, B1 => n545, B2 => n5095
                           , ZN => n3071);
   U7925 : OAI22_X1 port map( A1 => n7338, A2 => n7550, B1 => n520, B2 => n5093
                           , ZN => n3096);
   U7926 : OAI22_X1 port map( A1 => n7339, A2 => n7553, B1 => n519, B2 => n5093
                           , ZN => n3097);
   U7927 : OAI22_X1 port map( A1 => n7339, A2 => n7556, B1 => n518, B2 => n5093
                           , ZN => n3098);
   U7928 : OAI22_X1 port map( A1 => n7339, A2 => n7559, B1 => n517, B2 => n5093
                           , ZN => n3099);
   U7929 : OAI22_X1 port map( A1 => n7339, A2 => n7562, B1 => n516, B2 => n5093
                           , ZN => n3100);
   U7930 : OAI22_X1 port map( A1 => n7339, A2 => n7565, B1 => n515, B2 => n5093
                           , ZN => n3101);
   U7931 : OAI22_X1 port map( A1 => n7340, A2 => n7568, B1 => n514, B2 => n5093
                           , ZN => n3102);
   U7932 : OAI22_X1 port map( A1 => n7340, A2 => n7580, B1 => n513, B2 => n5093
                           , ZN => n3103);
   U7933 : OAI22_X1 port map( A1 => n7347, A2 => n7550, B1 => n488, B2 => n5092
                           , ZN => n3128);
   U7934 : OAI22_X1 port map( A1 => n7348, A2 => n7553, B1 => n487, B2 => n5092
                           , ZN => n3129);
   U7935 : OAI22_X1 port map( A1 => n7348, A2 => n7556, B1 => n486, B2 => n5092
                           , ZN => n3130);
   U7936 : OAI22_X1 port map( A1 => n7348, A2 => n7559, B1 => n485, B2 => n5092
                           , ZN => n3131);
   U7937 : OAI22_X1 port map( A1 => n7348, A2 => n7562, B1 => n484, B2 => n5092
                           , ZN => n3132);
   U7938 : OAI22_X1 port map( A1 => n7348, A2 => n7565, B1 => n483, B2 => n5092
                           , ZN => n3133);
   U7939 : OAI22_X1 port map( A1 => n7349, A2 => n7568, B1 => n482, B2 => n5092
                           , ZN => n3134);
   U7940 : OAI22_X1 port map( A1 => n7349, A2 => n7580, B1 => n481, B2 => n5092
                           , ZN => n3135);
   U7941 : OAI22_X1 port map( A1 => n7356, A2 => n7550, B1 => n456, B2 => n5091
                           , ZN => n3160);
   U7942 : OAI22_X1 port map( A1 => n7357, A2 => n7553, B1 => n455, B2 => n5091
                           , ZN => n3161);
   U7943 : OAI22_X1 port map( A1 => n7357, A2 => n7556, B1 => n454, B2 => n5091
                           , ZN => n3162);
   U7944 : OAI22_X1 port map( A1 => n7357, A2 => n7559, B1 => n453, B2 => n5091
                           , ZN => n3163);
   U7945 : OAI22_X1 port map( A1 => n7357, A2 => n7562, B1 => n452, B2 => n5091
                           , ZN => n3164);
   U7946 : OAI22_X1 port map( A1 => n7357, A2 => n7565, B1 => n451, B2 => n5091
                           , ZN => n3165);
   U7947 : OAI22_X1 port map( A1 => n7358, A2 => n7568, B1 => n450, B2 => n5091
                           , ZN => n3166);
   U7948 : OAI22_X1 port map( A1 => n7358, A2 => n7580, B1 => n449, B2 => n5091
                           , ZN => n3167);
   U7949 : OAI22_X1 port map( A1 => n7401, A2 => n7549, B1 => n296, B2 => n5086
                           , ZN => n3320);
   U7950 : OAI22_X1 port map( A1 => n7402, A2 => n7552, B1 => n295, B2 => n5086
                           , ZN => n3321);
   U7951 : OAI22_X1 port map( A1 => n7402, A2 => n7555, B1 => n294, B2 => n5086
                           , ZN => n3322);
   U7952 : OAI22_X1 port map( A1 => n7402, A2 => n7558, B1 => n293, B2 => n5086
                           , ZN => n3323);
   U7953 : OAI22_X1 port map( A1 => n7402, A2 => n7561, B1 => n292, B2 => n5086
                           , ZN => n3324);
   U7954 : OAI22_X1 port map( A1 => n7402, A2 => n7564, B1 => n291, B2 => n5086
                           , ZN => n3325);
   U7955 : OAI22_X1 port map( A1 => n7403, A2 => n7567, B1 => n290, B2 => n5086
                           , ZN => n3326);
   U7956 : OAI22_X1 port map( A1 => n7403, A2 => n7579, B1 => n289, B2 => n5086
                           , ZN => n3327);
   U7957 : OAI22_X1 port map( A1 => n7410, A2 => n7549, B1 => n264, B2 => n5084
                           , ZN => n3352);
   U7958 : OAI22_X1 port map( A1 => n7411, A2 => n7552, B1 => n263, B2 => n5084
                           , ZN => n3353);
   U7959 : OAI22_X1 port map( A1 => n7411, A2 => n7555, B1 => n262, B2 => n5084
                           , ZN => n3354);
   U7960 : OAI22_X1 port map( A1 => n7411, A2 => n7558, B1 => n261, B2 => n5084
                           , ZN => n3355);
   U7961 : OAI22_X1 port map( A1 => n7411, A2 => n7561, B1 => n260, B2 => n5084
                           , ZN => n3356);
   U7962 : OAI22_X1 port map( A1 => n7411, A2 => n7564, B1 => n259, B2 => n5084
                           , ZN => n3357);
   U7963 : OAI22_X1 port map( A1 => n7412, A2 => n7567, B1 => n258, B2 => n5084
                           , ZN => n3358);
   U7964 : OAI22_X1 port map( A1 => n7412, A2 => n7579, B1 => n257, B2 => n5084
                           , ZN => n3359);
   U7965 : OAI22_X1 port map( A1 => n7419, A2 => n7549, B1 => n232, B2 => n5081
                           , ZN => n3384);
   U7966 : OAI22_X1 port map( A1 => n7420, A2 => n7552, B1 => n231, B2 => n5081
                           , ZN => n3385);
   U7967 : OAI22_X1 port map( A1 => n7420, A2 => n7555, B1 => n230, B2 => n5081
                           , ZN => n3386);
   U7968 : OAI22_X1 port map( A1 => n7420, A2 => n7558, B1 => n229, B2 => n5081
                           , ZN => n3387);
   U7969 : OAI22_X1 port map( A1 => n7420, A2 => n7561, B1 => n228, B2 => n5081
                           , ZN => n3388);
   U7970 : OAI22_X1 port map( A1 => n7420, A2 => n7564, B1 => n227, B2 => n5081
                           , ZN => n3389);
   U7971 : OAI22_X1 port map( A1 => n7421, A2 => n7567, B1 => n226, B2 => n5081
                           , ZN => n3390);
   U7972 : OAI22_X1 port map( A1 => n7421, A2 => n7579, B1 => n225, B2 => n5081
                           , ZN => n3391);
   U7973 : OAI22_X1 port map( A1 => n7428, A2 => n7549, B1 => n200, B2 => n5079
                           , ZN => n3416);
   U7974 : OAI22_X1 port map( A1 => n7429, A2 => n7552, B1 => n199, B2 => n5079
                           , ZN => n3417);
   U7975 : OAI22_X1 port map( A1 => n7429, A2 => n7555, B1 => n198, B2 => n5079
                           , ZN => n3418);
   U7976 : OAI22_X1 port map( A1 => n7429, A2 => n7558, B1 => n197, B2 => n5079
                           , ZN => n3419);
   U7977 : OAI22_X1 port map( A1 => n7429, A2 => n7561, B1 => n196, B2 => n5079
                           , ZN => n3420);
   U7978 : OAI22_X1 port map( A1 => n7429, A2 => n7564, B1 => n195, B2 => n5079
                           , ZN => n3421);
   U7979 : OAI22_X1 port map( A1 => n7430, A2 => n7567, B1 => n194, B2 => n5079
                           , ZN => n3422);
   U7980 : OAI22_X1 port map( A1 => n7430, A2 => n7579, B1 => n193, B2 => n5079
                           , ZN => n3423);
   U7981 : OAI22_X1 port map( A1 => n7473, A2 => n7549, B1 => n40, B2 => n5069,
                           ZN => n3576);
   U7982 : OAI22_X1 port map( A1 => n7474, A2 => n7552, B1 => n39, B2 => n5069,
                           ZN => n3577);
   U7983 : OAI22_X1 port map( A1 => n7474, A2 => n7555, B1 => n38, B2 => n5069,
                           ZN => n3578);
   U7984 : OAI22_X1 port map( A1 => n7474, A2 => n7558, B1 => n37, B2 => n5069,
                           ZN => n3579);
   U7985 : OAI22_X1 port map( A1 => n7474, A2 => n7561, B1 => n36, B2 => n5069,
                           ZN => n3580);
   U7986 : OAI22_X1 port map( A1 => n7474, A2 => n7564, B1 => n35, B2 => n5069,
                           ZN => n3581);
   U7987 : OAI22_X1 port map( A1 => n7475, A2 => n7567, B1 => n34, B2 => n5069,
                           ZN => n3582);
   U7988 : OAI22_X1 port map( A1 => n7475, A2 => n7579, B1 => n33, B2 => n5069,
                           ZN => n3583);
   U7989 : OAI22_X1 port map( A1 => n7575, A2 => n7549, B1 => n8, B2 => n5035, 
                           ZN => n3608);
   U7990 : OAI22_X1 port map( A1 => n7576, A2 => n7552, B1 => n7, B2 => n5035, 
                           ZN => n3609);
   U7991 : OAI22_X1 port map( A1 => n7576, A2 => n7555, B1 => n6, B2 => n5035, 
                           ZN => n3610);
   U7992 : OAI22_X1 port map( A1 => n7576, A2 => n7558, B1 => n5, B2 => n5035, 
                           ZN => n3611);
   U7993 : OAI22_X1 port map( A1 => n7576, A2 => n7561, B1 => n4, B2 => n5035, 
                           ZN => n3612);
   U7994 : OAI22_X1 port map( A1 => n7576, A2 => n7564, B1 => n3, B2 => n5035, 
                           ZN => n3613);
   U7995 : OAI22_X1 port map( A1 => n7577, A2 => n7567, B1 => n2, B2 => n5035, 
                           ZN => n3614);
   U7996 : OAI22_X1 port map( A1 => n7577, A2 => n7579, B1 => n1, B2 => n5035, 
                           ZN => n3615);
   U7997 : OAI22_X1 port map( A1 => n7244, A2 => n7479, B1 => n7243, B2 => 
                           n4873, ZN => n2752);
   U7998 : OAI22_X1 port map( A1 => n7244, A2 => n7482, B1 => n7243, B2 => 
                           n4872, ZN => n2753);
   U7999 : OAI22_X1 port map( A1 => n7244, A2 => n7485, B1 => n7243, B2 => 
                           n4871, ZN => n2754);
   U8000 : OAI22_X1 port map( A1 => n7244, A2 => n7488, B1 => n7243, B2 => 
                           n4870, ZN => n2755);
   U8001 : OAI22_X1 port map( A1 => n7244, A2 => n7491, B1 => n7243, B2 => 
                           n4869, ZN => n2756);
   U8002 : OAI22_X1 port map( A1 => n7245, A2 => n7494, B1 => n7243, B2 => 
                           n4868, ZN => n2757);
   U8003 : OAI22_X1 port map( A1 => n7245, A2 => n7497, B1 => n7243, B2 => 
                           n4867, ZN => n2758);
   U8004 : OAI22_X1 port map( A1 => n7245, A2 => n7500, B1 => n7243, B2 => 
                           n4866, ZN => n2759);
   U8005 : OAI22_X1 port map( A1 => n7245, A2 => n7503, B1 => n7243, B2 => 
                           n4865, ZN => n2760);
   U8006 : OAI22_X1 port map( A1 => n7245, A2 => n7506, B1 => n7243, B2 => 
                           n4864, ZN => n2761);
   U8007 : OAI22_X1 port map( A1 => n7246, A2 => n7509, B1 => n7243, B2 => 
                           n4863, ZN => n2762);
   U8008 : OAI22_X1 port map( A1 => n7246, A2 => n7512, B1 => n7243, B2 => 
                           n4862, ZN => n2763);
   U8009 : OAI22_X1 port map( A1 => n7246, A2 => n7515, B1 => n5105, B2 => 
                           n4861, ZN => n2764);
   U8010 : OAI22_X1 port map( A1 => n7246, A2 => n7518, B1 => n5105, B2 => 
                           n4860, ZN => n2765);
   U8011 : OAI22_X1 port map( A1 => n7246, A2 => n7521, B1 => n5105, B2 => 
                           n4859, ZN => n2766);
   U8012 : OAI22_X1 port map( A1 => n7247, A2 => n7524, B1 => n7243, B2 => 
                           n4858, ZN => n2767);
   U8013 : OAI22_X1 port map( A1 => n7247, A2 => n7527, B1 => n7243, B2 => 
                           n4857, ZN => n2768);
   U8014 : OAI22_X1 port map( A1 => n7247, A2 => n7530, B1 => n7243, B2 => 
                           n4856, ZN => n2769);
   U8015 : OAI22_X1 port map( A1 => n7247, A2 => n7533, B1 => n7243, B2 => 
                           n4855, ZN => n2770);
   U8016 : OAI22_X1 port map( A1 => n7247, A2 => n7536, B1 => n7243, B2 => 
                           n4854, ZN => n2771);
   U8017 : OAI22_X1 port map( A1 => n7248, A2 => n7539, B1 => n7243, B2 => 
                           n4853, ZN => n2772);
   U8018 : OAI22_X1 port map( A1 => n7248, A2 => n7542, B1 => n7243, B2 => 
                           n4852, ZN => n2773);
   U8019 : OAI22_X1 port map( A1 => n7248, A2 => n7545, B1 => n7243, B2 => 
                           n4851, ZN => n2774);
   U8020 : OAI22_X1 port map( A1 => n7248, A2 => n7548, B1 => n7243, B2 => 
                           n4850, ZN => n2775);
   U8021 : OAI22_X1 port map( A1 => n7316, A2 => n7478, B1 => n7315, B2 => 
                           n4681, ZN => n3008);
   U8022 : OAI22_X1 port map( A1 => n7316, A2 => n7481, B1 => n7315, B2 => 
                           n4680, ZN => n3009);
   U8023 : OAI22_X1 port map( A1 => n7316, A2 => n7484, B1 => n7315, B2 => 
                           n4679, ZN => n3010);
   U8024 : OAI22_X1 port map( A1 => n7316, A2 => n7487, B1 => n7315, B2 => 
                           n4678, ZN => n3011);
   U8025 : OAI22_X1 port map( A1 => n7316, A2 => n7490, B1 => n7315, B2 => 
                           n4677, ZN => n3012);
   U8026 : OAI22_X1 port map( A1 => n7317, A2 => n7493, B1 => n7315, B2 => 
                           n4676, ZN => n3013);
   U8027 : OAI22_X1 port map( A1 => n7317, A2 => n7496, B1 => n7315, B2 => 
                           n4675, ZN => n3014);
   U8028 : OAI22_X1 port map( A1 => n7317, A2 => n7499, B1 => n7315, B2 => 
                           n4674, ZN => n3015);
   U8029 : OAI22_X1 port map( A1 => n7317, A2 => n7502, B1 => n7315, B2 => 
                           n4673, ZN => n3016);
   U8030 : OAI22_X1 port map( A1 => n7317, A2 => n7505, B1 => n7315, B2 => 
                           n4672, ZN => n3017);
   U8031 : OAI22_X1 port map( A1 => n7318, A2 => n7508, B1 => n7315, B2 => 
                           n4671, ZN => n3018);
   U8032 : OAI22_X1 port map( A1 => n7318, A2 => n7511, B1 => n7315, B2 => 
                           n4670, ZN => n3019);
   U8033 : OAI22_X1 port map( A1 => n7318, A2 => n7514, B1 => n5096, B2 => 
                           n4669, ZN => n3020);
   U8034 : OAI22_X1 port map( A1 => n7318, A2 => n7517, B1 => n5096, B2 => 
                           n4668, ZN => n3021);
   U8035 : OAI22_X1 port map( A1 => n7318, A2 => n7520, B1 => n5096, B2 => 
                           n4667, ZN => n3022);
   U8036 : OAI22_X1 port map( A1 => n7319, A2 => n7523, B1 => n7315, B2 => 
                           n4666, ZN => n3023);
   U8037 : OAI22_X1 port map( A1 => n7319, A2 => n7526, B1 => n7315, B2 => 
                           n4665, ZN => n3024);
   U8038 : OAI22_X1 port map( A1 => n7319, A2 => n7529, B1 => n7315, B2 => 
                           n4664, ZN => n3025);
   U8039 : OAI22_X1 port map( A1 => n7319, A2 => n7532, B1 => n7315, B2 => 
                           n4663, ZN => n3026);
   U8040 : OAI22_X1 port map( A1 => n7319, A2 => n7535, B1 => n7315, B2 => 
                           n4662, ZN => n3027);
   U8041 : OAI22_X1 port map( A1 => n7320, A2 => n7538, B1 => n7315, B2 => 
                           n4661, ZN => n3028);
   U8042 : OAI22_X1 port map( A1 => n7320, A2 => n7541, B1 => n7315, B2 => 
                           n4660, ZN => n3029);
   U8043 : OAI22_X1 port map( A1 => n7320, A2 => n7544, B1 => n7315, B2 => 
                           n4659, ZN => n3030);
   U8044 : OAI22_X1 port map( A1 => n7320, A2 => n7547, B1 => n7315, B2 => 
                           n4658, ZN => n3031);
   U8045 : OAI22_X1 port map( A1 => n7388, A2 => n7477, B1 => n7387, B2 => 
                           n4489, ZN => n3264);
   U8046 : OAI22_X1 port map( A1 => n7388, A2 => n7480, B1 => n7387, B2 => 
                           n4488, ZN => n3265);
   U8047 : OAI22_X1 port map( A1 => n7388, A2 => n7483, B1 => n7387, B2 => 
                           n4487, ZN => n3266);
   U8048 : OAI22_X1 port map( A1 => n7388, A2 => n7486, B1 => n7387, B2 => 
                           n4486, ZN => n3267);
   U8049 : OAI22_X1 port map( A1 => n7388, A2 => n7489, B1 => n7387, B2 => 
                           n4485, ZN => n3268);
   U8050 : OAI22_X1 port map( A1 => n7389, A2 => n7492, B1 => n7387, B2 => 
                           n4484, ZN => n3269);
   U8051 : OAI22_X1 port map( A1 => n7389, A2 => n7495, B1 => n7387, B2 => 
                           n4483, ZN => n3270);
   U8052 : OAI22_X1 port map( A1 => n7389, A2 => n7498, B1 => n7387, B2 => 
                           n4482, ZN => n3271);
   U8053 : OAI22_X1 port map( A1 => n7389, A2 => n7501, B1 => n7387, B2 => 
                           n4481, ZN => n3272);
   U8054 : OAI22_X1 port map( A1 => n7389, A2 => n7504, B1 => n7387, B2 => 
                           n4480, ZN => n3273);
   U8055 : OAI22_X1 port map( A1 => n7390, A2 => n7507, B1 => n7387, B2 => 
                           n4479, ZN => n3274);
   U8056 : OAI22_X1 port map( A1 => n7390, A2 => n7510, B1 => n7387, B2 => 
                           n4478, ZN => n3275);
   U8057 : OAI22_X1 port map( A1 => n7390, A2 => n7513, B1 => n5087, B2 => 
                           n4477, ZN => n3276);
   U8058 : OAI22_X1 port map( A1 => n7390, A2 => n7516, B1 => n5087, B2 => 
                           n4476, ZN => n3277);
   U8059 : OAI22_X1 port map( A1 => n7390, A2 => n7519, B1 => n5087, B2 => 
                           n4475, ZN => n3278);
   U8060 : OAI22_X1 port map( A1 => n7391, A2 => n7522, B1 => n7387, B2 => 
                           n4474, ZN => n3279);
   U8061 : OAI22_X1 port map( A1 => n7391, A2 => n7525, B1 => n7387, B2 => 
                           n4473, ZN => n3280);
   U8062 : OAI22_X1 port map( A1 => n7391, A2 => n7528, B1 => n7387, B2 => 
                           n4472, ZN => n3281);
   U8063 : OAI22_X1 port map( A1 => n7391, A2 => n7531, B1 => n7387, B2 => 
                           n4471, ZN => n3282);
   U8064 : OAI22_X1 port map( A1 => n7391, A2 => n7534, B1 => n7387, B2 => 
                           n4470, ZN => n3283);
   U8065 : OAI22_X1 port map( A1 => n7392, A2 => n7537, B1 => n7387, B2 => 
                           n4469, ZN => n3284);
   U8066 : OAI22_X1 port map( A1 => n7392, A2 => n7540, B1 => n7387, B2 => 
                           n4468, ZN => n3285);
   U8067 : OAI22_X1 port map( A1 => n7392, A2 => n7543, B1 => n7387, B2 => 
                           n4467, ZN => n3286);
   U8068 : OAI22_X1 port map( A1 => n7392, A2 => n7546, B1 => n7387, B2 => 
                           n4466, ZN => n3287);
   U8069 : OAI22_X1 port map( A1 => n7460, A2 => n7477, B1 => n7459, B2 => 
                           n4297, ZN => n3520);
   U8070 : OAI22_X1 port map( A1 => n7460, A2 => n7480, B1 => n7459, B2 => 
                           n4296, ZN => n3521);
   U8071 : OAI22_X1 port map( A1 => n7460, A2 => n7483, B1 => n7459, B2 => 
                           n4295, ZN => n3522);
   U8072 : OAI22_X1 port map( A1 => n7460, A2 => n7486, B1 => n7459, B2 => 
                           n4294, ZN => n3523);
   U8073 : OAI22_X1 port map( A1 => n7460, A2 => n7489, B1 => n7459, B2 => 
                           n4293, ZN => n3524);
   U8074 : OAI22_X1 port map( A1 => n7461, A2 => n7492, B1 => n7459, B2 => 
                           n4292, ZN => n3525);
   U8075 : OAI22_X1 port map( A1 => n7461, A2 => n7495, B1 => n7459, B2 => 
                           n4291, ZN => n3526);
   U8076 : OAI22_X1 port map( A1 => n7461, A2 => n7498, B1 => n7459, B2 => 
                           n4290, ZN => n3527);
   U8077 : OAI22_X1 port map( A1 => n7461, A2 => n7501, B1 => n7459, B2 => 
                           n4289, ZN => n3528);
   U8078 : OAI22_X1 port map( A1 => n7461, A2 => n7504, B1 => n7459, B2 => 
                           n4288, ZN => n3529);
   U8079 : OAI22_X1 port map( A1 => n7462, A2 => n7507, B1 => n7459, B2 => 
                           n4287, ZN => n3530);
   U8080 : OAI22_X1 port map( A1 => n7462, A2 => n7510, B1 => n7459, B2 => 
                           n4286, ZN => n3531);
   U8081 : OAI22_X1 port map( A1 => n7462, A2 => n7513, B1 => n5071, B2 => 
                           n4285, ZN => n3532);
   U8082 : OAI22_X1 port map( A1 => n7462, A2 => n7516, B1 => n5071, B2 => 
                           n4284, ZN => n3533);
   U8083 : OAI22_X1 port map( A1 => n7462, A2 => n7519, B1 => n5071, B2 => 
                           n4283, ZN => n3534);
   U8084 : OAI22_X1 port map( A1 => n7463, A2 => n7522, B1 => n7459, B2 => 
                           n4282, ZN => n3535);
   U8085 : OAI22_X1 port map( A1 => n7463, A2 => n7525, B1 => n7459, B2 => 
                           n4281, ZN => n3536);
   U8086 : OAI22_X1 port map( A1 => n7463, A2 => n7528, B1 => n7459, B2 => 
                           n4280, ZN => n3537);
   U8087 : OAI22_X1 port map( A1 => n7463, A2 => n7531, B1 => n7459, B2 => 
                           n4279, ZN => n3538);
   U8088 : OAI22_X1 port map( A1 => n7463, A2 => n7534, B1 => n7459, B2 => 
                           n4278, ZN => n3539);
   U8089 : OAI22_X1 port map( A1 => n7464, A2 => n7537, B1 => n7459, B2 => 
                           n4277, ZN => n3540);
   U8090 : OAI22_X1 port map( A1 => n7464, A2 => n7540, B1 => n7459, B2 => 
                           n4276, ZN => n3541);
   U8091 : OAI22_X1 port map( A1 => n7464, A2 => n7543, B1 => n7459, B2 => 
                           n4275, ZN => n3542);
   U8092 : OAI22_X1 port map( A1 => n7464, A2 => n7546, B1 => n7459, B2 => 
                           n4274, ZN => n3543);
   U8093 : OAI22_X1 port map( A1 => n1024, A2 => n5110, B1 => n7198, B2 => 
                           n7479, ZN => n2561);
   U8094 : OAI22_X1 port map( A1 => n1023, A2 => n7197, B1 => n7198, B2 => 
                           n7482, ZN => n2563);
   U8095 : OAI22_X1 port map( A1 => n1022, A2 => n7197, B1 => n7198, B2 => 
                           n7485, ZN => n2565);
   U8096 : OAI22_X1 port map( A1 => n1021, A2 => n7197, B1 => n7198, B2 => 
                           n7488, ZN => n2567);
   U8097 : OAI22_X1 port map( A1 => n1020, A2 => n7197, B1 => n7199, B2 => 
                           n7491, ZN => n2569);
   U8098 : OAI22_X1 port map( A1 => n1019, A2 => n7197, B1 => n7199, B2 => 
                           n7494, ZN => n2571);
   U8099 : OAI22_X1 port map( A1 => n1018, A2 => n7197, B1 => n7199, B2 => 
                           n7497, ZN => n2573);
   U8100 : OAI22_X1 port map( A1 => n1017, A2 => n7197, B1 => n7199, B2 => 
                           n7500, ZN => n2575);
   U8101 : OAI22_X1 port map( A1 => n1016, A2 => n7197, B1 => n7200, B2 => 
                           n7503, ZN => n2577);
   U8102 : OAI22_X1 port map( A1 => n1015, A2 => n7197, B1 => n7200, B2 => 
                           n7506, ZN => n2579);
   U8103 : OAI22_X1 port map( A1 => n1014, A2 => n7197, B1 => n7200, B2 => 
                           n7509, ZN => n2581);
   U8104 : OAI22_X1 port map( A1 => n1013, A2 => n7197, B1 => n7200, B2 => 
                           n7512, ZN => n2583);
   U8105 : OAI22_X1 port map( A1 => n1012, A2 => n5110, B1 => n7201, B2 => 
                           n7515, ZN => n2585);
   U8106 : OAI22_X1 port map( A1 => n1011, A2 => n7197, B1 => n7201, B2 => 
                           n7518, ZN => n2587);
   U8107 : OAI22_X1 port map( A1 => n1010, A2 => n5110, B1 => n7201, B2 => 
                           n7521, ZN => n2589);
   U8108 : OAI22_X1 port map( A1 => n1009, A2 => n7197, B1 => n7201, B2 => 
                           n7524, ZN => n2591);
   U8109 : OAI22_X1 port map( A1 => n1008, A2 => n5110, B1 => n7202, B2 => 
                           n7527, ZN => n2593);
   U8110 : OAI22_X1 port map( A1 => n1007, A2 => n7197, B1 => n7202, B2 => 
                           n7530, ZN => n2595);
   U8111 : OAI22_X1 port map( A1 => n1006, A2 => n5110, B1 => n7202, B2 => 
                           n7533, ZN => n2597);
   U8112 : OAI22_X1 port map( A1 => n1005, A2 => n7197, B1 => n7202, B2 => 
                           n7536, ZN => n2599);
   U8113 : OAI22_X1 port map( A1 => n1004, A2 => n5110, B1 => n7203, B2 => 
                           n7539, ZN => n2601);
   U8114 : OAI22_X1 port map( A1 => n1003, A2 => n7197, B1 => n7203, B2 => 
                           n7542, ZN => n2603);
   U8115 : OAI22_X1 port map( A1 => n1002, A2 => n5110, B1 => n7203, B2 => 
                           n7545, ZN => n2605);
   U8116 : OAI22_X1 port map( A1 => n1001, A2 => n7197, B1 => n7203, B2 => 
                           n7548, ZN => n2607);
   U8117 : OAI22_X1 port map( A1 => n1000, A2 => n5110, B1 => n7204, B2 => 
                           n7551, ZN => n2609);
   U8118 : OAI22_X1 port map( A1 => n999, A2 => n7197, B1 => n7204, B2 => n7554
                           , ZN => n2611);
   U8119 : OAI22_X1 port map( A1 => n998, A2 => n5110, B1 => n7204, B2 => n7557
                           , ZN => n2613);
   U8120 : OAI22_X1 port map( A1 => n997, A2 => n7197, B1 => n7204, B2 => n7560
                           , ZN => n2615);
   U8121 : OAI22_X1 port map( A1 => n996, A2 => n5110, B1 => n7205, B2 => n7563
                           , ZN => n2617);
   U8122 : OAI22_X1 port map( A1 => n995, A2 => n7197, B1 => n7205, B2 => n7566
                           , ZN => n2619);
   U8123 : OAI22_X1 port map( A1 => n994, A2 => n5110, B1 => n7205, B2 => n7569
                           , ZN => n2621);
   U8124 : OAI22_X1 port map( A1 => n993, A2 => n7197, B1 => n7205, B2 => n7581
                           , ZN => n2623);
   U8125 : OAI22_X1 port map( A1 => n7208, A2 => n7479, B1 => n992, B2 => n7207
                           , ZN => n2624);
   U8126 : OAI22_X1 port map( A1 => n7208, A2 => n7482, B1 => n991, B2 => n7207
                           , ZN => n2625);
   U8127 : OAI22_X1 port map( A1 => n7208, A2 => n7485, B1 => n990, B2 => n7207
                           , ZN => n2626);
   U8128 : OAI22_X1 port map( A1 => n7208, A2 => n7488, B1 => n989, B2 => n7207
                           , ZN => n2627);
   U8129 : OAI22_X1 port map( A1 => n7208, A2 => n7491, B1 => n988, B2 => n7207
                           , ZN => n2628);
   U8130 : OAI22_X1 port map( A1 => n7209, A2 => n7494, B1 => n987, B2 => n7207
                           , ZN => n2629);
   U8131 : OAI22_X1 port map( A1 => n7209, A2 => n7497, B1 => n986, B2 => n7207
                           , ZN => n2630);
   U8132 : OAI22_X1 port map( A1 => n7209, A2 => n7500, B1 => n985, B2 => n7207
                           , ZN => n2631);
   U8133 : OAI22_X1 port map( A1 => n7209, A2 => n7503, B1 => n984, B2 => n7207
                           , ZN => n2632);
   U8134 : OAI22_X1 port map( A1 => n7209, A2 => n7506, B1 => n983, B2 => n7207
                           , ZN => n2633);
   U8135 : OAI22_X1 port map( A1 => n7210, A2 => n7509, B1 => n982, B2 => n7207
                           , ZN => n2634);
   U8136 : OAI22_X1 port map( A1 => n7210, A2 => n7512, B1 => n981, B2 => n7207
                           , ZN => n2635);
   U8137 : OAI22_X1 port map( A1 => n7210, A2 => n7515, B1 => n980, B2 => n5109
                           , ZN => n2636);
   U8138 : OAI22_X1 port map( A1 => n7210, A2 => n7518, B1 => n979, B2 => n5109
                           , ZN => n2637);
   U8139 : OAI22_X1 port map( A1 => n7210, A2 => n7521, B1 => n978, B2 => n5109
                           , ZN => n2638);
   U8140 : OAI22_X1 port map( A1 => n7211, A2 => n7524, B1 => n977, B2 => n7207
                           , ZN => n2639);
   U8141 : OAI22_X1 port map( A1 => n7211, A2 => n7527, B1 => n976, B2 => n7207
                           , ZN => n2640);
   U8142 : OAI22_X1 port map( A1 => n7211, A2 => n7530, B1 => n975, B2 => n7207
                           , ZN => n2641);
   U8143 : OAI22_X1 port map( A1 => n7211, A2 => n7533, B1 => n974, B2 => n7207
                           , ZN => n2642);
   U8144 : OAI22_X1 port map( A1 => n7211, A2 => n7536, B1 => n973, B2 => n7207
                           , ZN => n2643);
   U8145 : OAI22_X1 port map( A1 => n7212, A2 => n7539, B1 => n972, B2 => n7207
                           , ZN => n2644);
   U8146 : OAI22_X1 port map( A1 => n7212, A2 => n7542, B1 => n971, B2 => n7207
                           , ZN => n2645);
   U8147 : OAI22_X1 port map( A1 => n7212, A2 => n7545, B1 => n970, B2 => n7207
                           , ZN => n2646);
   U8148 : OAI22_X1 port map( A1 => n7212, A2 => n7548, B1 => n969, B2 => n7207
                           , ZN => n2647);
   U8149 : OAI22_X1 port map( A1 => n7253, A2 => n7479, B1 => n832, B2 => n7252
                           , ZN => n2784);
   U8150 : OAI22_X1 port map( A1 => n7253, A2 => n7482, B1 => n831, B2 => n7252
                           , ZN => n2785);
   U8151 : OAI22_X1 port map( A1 => n7253, A2 => n7485, B1 => n830, B2 => n7252
                           , ZN => n2786);
   U8152 : OAI22_X1 port map( A1 => n7253, A2 => n7488, B1 => n829, B2 => n7252
                           , ZN => n2787);
   U8153 : OAI22_X1 port map( A1 => n7253, A2 => n7491, B1 => n828, B2 => n7252
                           , ZN => n2788);
   U8154 : OAI22_X1 port map( A1 => n7254, A2 => n7494, B1 => n827, B2 => n7252
                           , ZN => n2789);
   U8155 : OAI22_X1 port map( A1 => n7254, A2 => n7497, B1 => n826, B2 => n7252
                           , ZN => n2790);
   U8156 : OAI22_X1 port map( A1 => n7254, A2 => n7500, B1 => n825, B2 => n7252
                           , ZN => n2791);
   U8157 : OAI22_X1 port map( A1 => n7254, A2 => n7503, B1 => n824, B2 => n7252
                           , ZN => n2792);
   U8158 : OAI22_X1 port map( A1 => n7254, A2 => n7506, B1 => n823, B2 => n7252
                           , ZN => n2793);
   U8159 : OAI22_X1 port map( A1 => n7255, A2 => n7509, B1 => n822, B2 => n7252
                           , ZN => n2794);
   U8160 : OAI22_X1 port map( A1 => n7255, A2 => n7512, B1 => n821, B2 => n7252
                           , ZN => n2795);
   U8161 : OAI22_X1 port map( A1 => n7255, A2 => n7515, B1 => n820, B2 => n5104
                           , ZN => n2796);
   U8162 : OAI22_X1 port map( A1 => n7255, A2 => n7518, B1 => n819, B2 => n5104
                           , ZN => n2797);
   U8163 : OAI22_X1 port map( A1 => n7255, A2 => n7521, B1 => n818, B2 => n5104
                           , ZN => n2798);
   U8164 : OAI22_X1 port map( A1 => n7256, A2 => n7524, B1 => n817, B2 => n7252
                           , ZN => n2799);
   U8165 : OAI22_X1 port map( A1 => n7256, A2 => n7527, B1 => n816, B2 => n7252
                           , ZN => n2800);
   U8166 : OAI22_X1 port map( A1 => n7256, A2 => n7530, B1 => n815, B2 => n7252
                           , ZN => n2801);
   U8167 : OAI22_X1 port map( A1 => n7256, A2 => n7533, B1 => n814, B2 => n7252
                           , ZN => n2802);
   U8168 : OAI22_X1 port map( A1 => n7256, A2 => n7536, B1 => n813, B2 => n7252
                           , ZN => n2803);
   U8169 : OAI22_X1 port map( A1 => n7257, A2 => n7539, B1 => n812, B2 => n7252
                           , ZN => n2804);
   U8170 : OAI22_X1 port map( A1 => n7257, A2 => n7542, B1 => n811, B2 => n7252
                           , ZN => n2805);
   U8171 : OAI22_X1 port map( A1 => n7257, A2 => n7545, B1 => n810, B2 => n7252
                           , ZN => n2806);
   U8172 : OAI22_X1 port map( A1 => n7257, A2 => n7548, B1 => n809, B2 => n7252
                           , ZN => n2807);
   U8173 : OAI22_X1 port map( A1 => n7262, A2 => n7479, B1 => n800, B2 => n7261
                           , ZN => n2816);
   U8174 : OAI22_X1 port map( A1 => n7262, A2 => n7482, B1 => n799, B2 => n7261
                           , ZN => n2817);
   U8175 : OAI22_X1 port map( A1 => n7262, A2 => n7485, B1 => n798, B2 => n7261
                           , ZN => n2818);
   U8176 : OAI22_X1 port map( A1 => n7262, A2 => n7488, B1 => n797, B2 => n7261
                           , ZN => n2819);
   U8177 : OAI22_X1 port map( A1 => n7262, A2 => n7491, B1 => n796, B2 => n7261
                           , ZN => n2820);
   U8178 : OAI22_X1 port map( A1 => n7263, A2 => n7494, B1 => n795, B2 => n7261
                           , ZN => n2821);
   U8179 : OAI22_X1 port map( A1 => n7263, A2 => n7497, B1 => n794, B2 => n7261
                           , ZN => n2822);
   U8180 : OAI22_X1 port map( A1 => n7263, A2 => n7500, B1 => n793, B2 => n7261
                           , ZN => n2823);
   U8181 : OAI22_X1 port map( A1 => n7263, A2 => n7503, B1 => n792, B2 => n7261
                           , ZN => n2824);
   U8182 : OAI22_X1 port map( A1 => n7263, A2 => n7506, B1 => n791, B2 => n7261
                           , ZN => n2825);
   U8183 : OAI22_X1 port map( A1 => n7264, A2 => n7509, B1 => n790, B2 => n7261
                           , ZN => n2826);
   U8184 : OAI22_X1 port map( A1 => n7264, A2 => n7512, B1 => n789, B2 => n7261
                           , ZN => n2827);
   U8185 : OAI22_X1 port map( A1 => n7264, A2 => n7515, B1 => n788, B2 => n5102
                           , ZN => n2828);
   U8186 : OAI22_X1 port map( A1 => n7264, A2 => n7518, B1 => n787, B2 => n5102
                           , ZN => n2829);
   U8187 : OAI22_X1 port map( A1 => n7264, A2 => n7521, B1 => n786, B2 => n5102
                           , ZN => n2830);
   U8188 : OAI22_X1 port map( A1 => n7265, A2 => n7524, B1 => n785, B2 => n7261
                           , ZN => n2831);
   U8189 : OAI22_X1 port map( A1 => n7265, A2 => n7527, B1 => n784, B2 => n7261
                           , ZN => n2832);
   U8190 : OAI22_X1 port map( A1 => n7265, A2 => n7530, B1 => n783, B2 => n7261
                           , ZN => n2833);
   U8191 : OAI22_X1 port map( A1 => n7265, A2 => n7533, B1 => n782, B2 => n7261
                           , ZN => n2834);
   U8192 : OAI22_X1 port map( A1 => n7265, A2 => n7536, B1 => n781, B2 => n7261
                           , ZN => n2835);
   U8193 : OAI22_X1 port map( A1 => n7266, A2 => n7539, B1 => n780, B2 => n7261
                           , ZN => n2836);
   U8194 : OAI22_X1 port map( A1 => n7266, A2 => n7542, B1 => n779, B2 => n7261
                           , ZN => n2837);
   U8195 : OAI22_X1 port map( A1 => n7266, A2 => n7545, B1 => n778, B2 => n7261
                           , ZN => n2838);
   U8196 : OAI22_X1 port map( A1 => n7266, A2 => n7548, B1 => n777, B2 => n7261
                           , ZN => n2839);
   U8197 : OAI22_X1 port map( A1 => n7271, A2 => n7478, B1 => n768, B2 => n7270
                           , ZN => n2848);
   U8198 : OAI22_X1 port map( A1 => n7271, A2 => n7481, B1 => n767, B2 => n7270
                           , ZN => n2849);
   U8199 : OAI22_X1 port map( A1 => n7271, A2 => n7484, B1 => n766, B2 => n7270
                           , ZN => n2850);
   U8200 : OAI22_X1 port map( A1 => n7271, A2 => n7487, B1 => n765, B2 => n7270
                           , ZN => n2851);
   U8201 : OAI22_X1 port map( A1 => n7271, A2 => n7490, B1 => n764, B2 => n7270
                           , ZN => n2852);
   U8202 : OAI22_X1 port map( A1 => n7272, A2 => n7493, B1 => n763, B2 => n7270
                           , ZN => n2853);
   U8203 : OAI22_X1 port map( A1 => n7272, A2 => n7496, B1 => n762, B2 => n7270
                           , ZN => n2854);
   U8204 : OAI22_X1 port map( A1 => n7272, A2 => n7499, B1 => n761, B2 => n7270
                           , ZN => n2855);
   U8205 : OAI22_X1 port map( A1 => n7272, A2 => n7502, B1 => n760, B2 => n7270
                           , ZN => n2856);
   U8206 : OAI22_X1 port map( A1 => n7272, A2 => n7505, B1 => n759, B2 => n7270
                           , ZN => n2857);
   U8207 : OAI22_X1 port map( A1 => n7273, A2 => n7508, B1 => n758, B2 => n7270
                           , ZN => n2858);
   U8208 : OAI22_X1 port map( A1 => n7273, A2 => n7511, B1 => n757, B2 => n7270
                           , ZN => n2859);
   U8209 : OAI22_X1 port map( A1 => n7273, A2 => n7514, B1 => n756, B2 => n5101
                           , ZN => n2860);
   U8210 : OAI22_X1 port map( A1 => n7273, A2 => n7517, B1 => n755, B2 => n5101
                           , ZN => n2861);
   U8211 : OAI22_X1 port map( A1 => n7273, A2 => n7520, B1 => n754, B2 => n5101
                           , ZN => n2862);
   U8212 : OAI22_X1 port map( A1 => n7274, A2 => n7523, B1 => n753, B2 => n7270
                           , ZN => n2863);
   U8213 : OAI22_X1 port map( A1 => n7274, A2 => n7526, B1 => n752, B2 => n7270
                           , ZN => n2864);
   U8214 : OAI22_X1 port map( A1 => n7274, A2 => n7529, B1 => n751, B2 => n7270
                           , ZN => n2865);
   U8215 : OAI22_X1 port map( A1 => n7274, A2 => n7532, B1 => n750, B2 => n7270
                           , ZN => n2866);
   U8216 : OAI22_X1 port map( A1 => n7274, A2 => n7535, B1 => n749, B2 => n7270
                           , ZN => n2867);
   U8217 : OAI22_X1 port map( A1 => n7275, A2 => n7538, B1 => n748, B2 => n7270
                           , ZN => n2868);
   U8218 : OAI22_X1 port map( A1 => n7275, A2 => n7541, B1 => n747, B2 => n7270
                           , ZN => n2869);
   U8219 : OAI22_X1 port map( A1 => n7275, A2 => n7544, B1 => n746, B2 => n7270
                           , ZN => n2870);
   U8220 : OAI22_X1 port map( A1 => n7275, A2 => n7547, B1 => n745, B2 => n7270
                           , ZN => n2871);
   U8221 : OAI22_X1 port map( A1 => n7280, A2 => n7478, B1 => n736, B2 => n7279
                           , ZN => n2880);
   U8222 : OAI22_X1 port map( A1 => n7280, A2 => n7481, B1 => n735, B2 => n7279
                           , ZN => n2881);
   U8223 : OAI22_X1 port map( A1 => n7280, A2 => n7484, B1 => n734, B2 => n7279
                           , ZN => n2882);
   U8224 : OAI22_X1 port map( A1 => n7280, A2 => n7487, B1 => n733, B2 => n7279
                           , ZN => n2883);
   U8225 : OAI22_X1 port map( A1 => n7280, A2 => n7490, B1 => n732, B2 => n7279
                           , ZN => n2884);
   U8226 : OAI22_X1 port map( A1 => n7281, A2 => n7493, B1 => n731, B2 => n7279
                           , ZN => n2885);
   U8227 : OAI22_X1 port map( A1 => n7281, A2 => n7496, B1 => n730, B2 => n7279
                           , ZN => n2886);
   U8228 : OAI22_X1 port map( A1 => n7281, A2 => n7499, B1 => n729, B2 => n7279
                           , ZN => n2887);
   U8229 : OAI22_X1 port map( A1 => n7281, A2 => n7502, B1 => n728, B2 => n7279
                           , ZN => n2888);
   U8230 : OAI22_X1 port map( A1 => n7281, A2 => n7505, B1 => n727, B2 => n7279
                           , ZN => n2889);
   U8231 : OAI22_X1 port map( A1 => n7282, A2 => n7508, B1 => n726, B2 => n7279
                           , ZN => n2890);
   U8232 : OAI22_X1 port map( A1 => n7282, A2 => n7511, B1 => n725, B2 => n7279
                           , ZN => n2891);
   U8233 : OAI22_X1 port map( A1 => n7282, A2 => n7514, B1 => n724, B2 => n5100
                           , ZN => n2892);
   U8234 : OAI22_X1 port map( A1 => n7282, A2 => n7517, B1 => n723, B2 => n5100
                           , ZN => n2893);
   U8235 : OAI22_X1 port map( A1 => n7282, A2 => n7520, B1 => n722, B2 => n5100
                           , ZN => n2894);
   U8236 : OAI22_X1 port map( A1 => n7283, A2 => n7523, B1 => n721, B2 => n7279
                           , ZN => n2895);
   U8237 : OAI22_X1 port map( A1 => n7283, A2 => n7526, B1 => n720, B2 => n7279
                           , ZN => n2896);
   U8238 : OAI22_X1 port map( A1 => n7283, A2 => n7529, B1 => n719, B2 => n7279
                           , ZN => n2897);
   U8239 : OAI22_X1 port map( A1 => n7283, A2 => n7532, B1 => n718, B2 => n7279
                           , ZN => n2898);
   U8240 : OAI22_X1 port map( A1 => n7283, A2 => n7535, B1 => n717, B2 => n7279
                           , ZN => n2899);
   U8241 : OAI22_X1 port map( A1 => n7284, A2 => n7538, B1 => n716, B2 => n7279
                           , ZN => n2900);
   U8242 : OAI22_X1 port map( A1 => n7284, A2 => n7541, B1 => n715, B2 => n7279
                           , ZN => n2901);
   U8243 : OAI22_X1 port map( A1 => n7284, A2 => n7544, B1 => n714, B2 => n7279
                           , ZN => n2902);
   U8244 : OAI22_X1 port map( A1 => n7284, A2 => n7547, B1 => n713, B2 => n7279
                           , ZN => n2903);
   U8245 : OAI22_X1 port map( A1 => n7325, A2 => n7478, B1 => n576, B2 => n7324
                           , ZN => n3040);
   U8246 : OAI22_X1 port map( A1 => n7325, A2 => n7481, B1 => n575, B2 => n7324
                           , ZN => n3041);
   U8247 : OAI22_X1 port map( A1 => n7325, A2 => n7484, B1 => n574, B2 => n7324
                           , ZN => n3042);
   U8248 : OAI22_X1 port map( A1 => n7325, A2 => n7487, B1 => n573, B2 => n7324
                           , ZN => n3043);
   U8249 : OAI22_X1 port map( A1 => n7325, A2 => n7490, B1 => n572, B2 => n7324
                           , ZN => n3044);
   U8250 : OAI22_X1 port map( A1 => n7326, A2 => n7493, B1 => n571, B2 => n7324
                           , ZN => n3045);
   U8251 : OAI22_X1 port map( A1 => n7326, A2 => n7496, B1 => n570, B2 => n7324
                           , ZN => n3046);
   U8252 : OAI22_X1 port map( A1 => n7326, A2 => n7499, B1 => n569, B2 => n7324
                           , ZN => n3047);
   U8253 : OAI22_X1 port map( A1 => n7326, A2 => n7502, B1 => n568, B2 => n7324
                           , ZN => n3048);
   U8254 : OAI22_X1 port map( A1 => n7326, A2 => n7505, B1 => n567, B2 => n7324
                           , ZN => n3049);
   U8255 : OAI22_X1 port map( A1 => n7327, A2 => n7508, B1 => n566, B2 => n7324
                           , ZN => n3050);
   U8256 : OAI22_X1 port map( A1 => n7327, A2 => n7511, B1 => n565, B2 => n7324
                           , ZN => n3051);
   U8257 : OAI22_X1 port map( A1 => n7327, A2 => n7514, B1 => n564, B2 => n5095
                           , ZN => n3052);
   U8258 : OAI22_X1 port map( A1 => n7327, A2 => n7517, B1 => n563, B2 => n5095
                           , ZN => n3053);
   U8259 : OAI22_X1 port map( A1 => n7327, A2 => n7520, B1 => n562, B2 => n5095
                           , ZN => n3054);
   U8260 : OAI22_X1 port map( A1 => n7328, A2 => n7523, B1 => n561, B2 => n7324
                           , ZN => n3055);
   U8261 : OAI22_X1 port map( A1 => n7328, A2 => n7526, B1 => n560, B2 => n7324
                           , ZN => n3056);
   U8262 : OAI22_X1 port map( A1 => n7328, A2 => n7529, B1 => n559, B2 => n7324
                           , ZN => n3057);
   U8263 : OAI22_X1 port map( A1 => n7328, A2 => n7532, B1 => n558, B2 => n7324
                           , ZN => n3058);
   U8264 : OAI22_X1 port map( A1 => n7328, A2 => n7535, B1 => n557, B2 => n7324
                           , ZN => n3059);
   U8265 : OAI22_X1 port map( A1 => n7329, A2 => n7538, B1 => n556, B2 => n7324
                           , ZN => n3060);
   U8266 : OAI22_X1 port map( A1 => n7329, A2 => n7541, B1 => n555, B2 => n7324
                           , ZN => n3061);
   U8267 : OAI22_X1 port map( A1 => n7329, A2 => n7544, B1 => n554, B2 => n7324
                           , ZN => n3062);
   U8268 : OAI22_X1 port map( A1 => n7329, A2 => n7547, B1 => n553, B2 => n7324
                           , ZN => n3063);
   U8269 : OAI22_X1 port map( A1 => n7334, A2 => n7478, B1 => n544, B2 => n7333
                           , ZN => n3072);
   U8270 : OAI22_X1 port map( A1 => n7334, A2 => n7481, B1 => n543, B2 => n7333
                           , ZN => n3073);
   U8271 : OAI22_X1 port map( A1 => n7334, A2 => n7484, B1 => n542, B2 => n7333
                           , ZN => n3074);
   U8272 : OAI22_X1 port map( A1 => n7334, A2 => n7487, B1 => n541, B2 => n7333
                           , ZN => n3075);
   U8273 : OAI22_X1 port map( A1 => n7334, A2 => n7490, B1 => n540, B2 => n7333
                           , ZN => n3076);
   U8274 : OAI22_X1 port map( A1 => n7335, A2 => n7493, B1 => n539, B2 => n7333
                           , ZN => n3077);
   U8275 : OAI22_X1 port map( A1 => n7335, A2 => n7496, B1 => n538, B2 => n7333
                           , ZN => n3078);
   U8276 : OAI22_X1 port map( A1 => n7335, A2 => n7499, B1 => n537, B2 => n7333
                           , ZN => n3079);
   U8277 : OAI22_X1 port map( A1 => n7335, A2 => n7502, B1 => n536, B2 => n7333
                           , ZN => n3080);
   U8278 : OAI22_X1 port map( A1 => n7335, A2 => n7505, B1 => n535, B2 => n7333
                           , ZN => n3081);
   U8279 : OAI22_X1 port map( A1 => n7336, A2 => n7508, B1 => n534, B2 => n7333
                           , ZN => n3082);
   U8280 : OAI22_X1 port map( A1 => n7336, A2 => n7511, B1 => n533, B2 => n7333
                           , ZN => n3083);
   U8281 : OAI22_X1 port map( A1 => n7336, A2 => n7514, B1 => n532, B2 => n5093
                           , ZN => n3084);
   U8282 : OAI22_X1 port map( A1 => n7336, A2 => n7517, B1 => n531, B2 => n5093
                           , ZN => n3085);
   U8283 : OAI22_X1 port map( A1 => n7336, A2 => n7520, B1 => n530, B2 => n5093
                           , ZN => n3086);
   U8284 : OAI22_X1 port map( A1 => n7337, A2 => n7523, B1 => n529, B2 => n7333
                           , ZN => n3087);
   U8285 : OAI22_X1 port map( A1 => n7337, A2 => n7526, B1 => n528, B2 => n7333
                           , ZN => n3088);
   U8286 : OAI22_X1 port map( A1 => n7337, A2 => n7529, B1 => n527, B2 => n7333
                           , ZN => n3089);
   U8287 : OAI22_X1 port map( A1 => n7337, A2 => n7532, B1 => n526, B2 => n7333
                           , ZN => n3090);
   U8288 : OAI22_X1 port map( A1 => n7337, A2 => n7535, B1 => n525, B2 => n7333
                           , ZN => n3091);
   U8289 : OAI22_X1 port map( A1 => n7338, A2 => n7538, B1 => n524, B2 => n7333
                           , ZN => n3092);
   U8290 : OAI22_X1 port map( A1 => n7338, A2 => n7541, B1 => n523, B2 => n7333
                           , ZN => n3093);
   U8291 : OAI22_X1 port map( A1 => n7338, A2 => n7544, B1 => n522, B2 => n7333
                           , ZN => n3094);
   U8292 : OAI22_X1 port map( A1 => n7338, A2 => n7547, B1 => n521, B2 => n7333
                           , ZN => n3095);
   U8293 : OAI22_X1 port map( A1 => n7343, A2 => n7478, B1 => n512, B2 => n7342
                           , ZN => n3104);
   U8294 : OAI22_X1 port map( A1 => n7343, A2 => n7481, B1 => n511, B2 => n7342
                           , ZN => n3105);
   U8295 : OAI22_X1 port map( A1 => n7343, A2 => n7484, B1 => n510, B2 => n7342
                           , ZN => n3106);
   U8296 : OAI22_X1 port map( A1 => n7343, A2 => n7487, B1 => n509, B2 => n7342
                           , ZN => n3107);
   U8297 : OAI22_X1 port map( A1 => n7343, A2 => n7490, B1 => n508, B2 => n7342
                           , ZN => n3108);
   U8298 : OAI22_X1 port map( A1 => n7344, A2 => n7493, B1 => n507, B2 => n7342
                           , ZN => n3109);
   U8299 : OAI22_X1 port map( A1 => n7344, A2 => n7496, B1 => n506, B2 => n7342
                           , ZN => n3110);
   U8300 : OAI22_X1 port map( A1 => n7344, A2 => n7499, B1 => n505, B2 => n7342
                           , ZN => n3111);
   U8301 : OAI22_X1 port map( A1 => n7344, A2 => n7502, B1 => n504, B2 => n7342
                           , ZN => n3112);
   U8302 : OAI22_X1 port map( A1 => n7344, A2 => n7505, B1 => n503, B2 => n7342
                           , ZN => n3113);
   U8303 : OAI22_X1 port map( A1 => n7345, A2 => n7508, B1 => n502, B2 => n7342
                           , ZN => n3114);
   U8304 : OAI22_X1 port map( A1 => n7345, A2 => n7511, B1 => n501, B2 => n7342
                           , ZN => n3115);
   U8305 : OAI22_X1 port map( A1 => n7345, A2 => n7514, B1 => n500, B2 => n5092
                           , ZN => n3116);
   U8306 : OAI22_X1 port map( A1 => n7345, A2 => n7517, B1 => n499, B2 => n5092
                           , ZN => n3117);
   U8307 : OAI22_X1 port map( A1 => n7345, A2 => n7520, B1 => n498, B2 => n5092
                           , ZN => n3118);
   U8308 : OAI22_X1 port map( A1 => n7346, A2 => n7523, B1 => n497, B2 => n7342
                           , ZN => n3119);
   U8309 : OAI22_X1 port map( A1 => n7346, A2 => n7526, B1 => n496, B2 => n7342
                           , ZN => n3120);
   U8310 : OAI22_X1 port map( A1 => n7346, A2 => n7529, B1 => n495, B2 => n7342
                           , ZN => n3121);
   U8311 : OAI22_X1 port map( A1 => n7346, A2 => n7532, B1 => n494, B2 => n7342
                           , ZN => n3122);
   U8312 : OAI22_X1 port map( A1 => n7346, A2 => n7535, B1 => n493, B2 => n7342
                           , ZN => n3123);
   U8313 : OAI22_X1 port map( A1 => n7347, A2 => n7538, B1 => n492, B2 => n7342
                           , ZN => n3124);
   U8314 : OAI22_X1 port map( A1 => n7347, A2 => n7541, B1 => n491, B2 => n7342
                           , ZN => n3125);
   U8315 : OAI22_X1 port map( A1 => n7347, A2 => n7544, B1 => n490, B2 => n7342
                           , ZN => n3126);
   U8316 : OAI22_X1 port map( A1 => n7347, A2 => n7547, B1 => n489, B2 => n7342
                           , ZN => n3127);
   U8317 : OAI22_X1 port map( A1 => n7352, A2 => n7478, B1 => n480, B2 => n7351
                           , ZN => n3136);
   U8318 : OAI22_X1 port map( A1 => n7352, A2 => n7481, B1 => n479, B2 => n7351
                           , ZN => n3137);
   U8319 : OAI22_X1 port map( A1 => n7352, A2 => n7484, B1 => n478, B2 => n7351
                           , ZN => n3138);
   U8320 : OAI22_X1 port map( A1 => n7352, A2 => n7487, B1 => n477, B2 => n7351
                           , ZN => n3139);
   U8321 : OAI22_X1 port map( A1 => n7352, A2 => n7490, B1 => n476, B2 => n7351
                           , ZN => n3140);
   U8322 : OAI22_X1 port map( A1 => n7353, A2 => n7493, B1 => n475, B2 => n7351
                           , ZN => n3141);
   U8323 : OAI22_X1 port map( A1 => n7353, A2 => n7496, B1 => n474, B2 => n7351
                           , ZN => n3142);
   U8324 : OAI22_X1 port map( A1 => n7353, A2 => n7499, B1 => n473, B2 => n7351
                           , ZN => n3143);
   U8325 : OAI22_X1 port map( A1 => n7353, A2 => n7502, B1 => n472, B2 => n7351
                           , ZN => n3144);
   U8326 : OAI22_X1 port map( A1 => n7353, A2 => n7505, B1 => n471, B2 => n7351
                           , ZN => n3145);
   U8327 : OAI22_X1 port map( A1 => n7354, A2 => n7508, B1 => n470, B2 => n7351
                           , ZN => n3146);
   U8328 : OAI22_X1 port map( A1 => n7354, A2 => n7511, B1 => n469, B2 => n7351
                           , ZN => n3147);
   U8329 : OAI22_X1 port map( A1 => n7354, A2 => n7514, B1 => n468, B2 => n5091
                           , ZN => n3148);
   U8330 : OAI22_X1 port map( A1 => n7354, A2 => n7517, B1 => n467, B2 => n5091
                           , ZN => n3149);
   U8331 : OAI22_X1 port map( A1 => n7354, A2 => n7520, B1 => n466, B2 => n5091
                           , ZN => n3150);
   U8332 : OAI22_X1 port map( A1 => n7355, A2 => n7523, B1 => n465, B2 => n7351
                           , ZN => n3151);
   U8333 : OAI22_X1 port map( A1 => n7355, A2 => n7526, B1 => n464, B2 => n7351
                           , ZN => n3152);
   U8334 : OAI22_X1 port map( A1 => n7355, A2 => n7529, B1 => n463, B2 => n7351
                           , ZN => n3153);
   U8335 : OAI22_X1 port map( A1 => n7355, A2 => n7532, B1 => n462, B2 => n7351
                           , ZN => n3154);
   U8336 : OAI22_X1 port map( A1 => n7355, A2 => n7535, B1 => n461, B2 => n7351
                           , ZN => n3155);
   U8337 : OAI22_X1 port map( A1 => n7356, A2 => n7538, B1 => n460, B2 => n7351
                           , ZN => n3156);
   U8338 : OAI22_X1 port map( A1 => n7356, A2 => n7541, B1 => n459, B2 => n7351
                           , ZN => n3157);
   U8339 : OAI22_X1 port map( A1 => n7356, A2 => n7544, B1 => n458, B2 => n7351
                           , ZN => n3158);
   U8340 : OAI22_X1 port map( A1 => n7356, A2 => n7547, B1 => n457, B2 => n7351
                           , ZN => n3159);
   U8341 : OAI22_X1 port map( A1 => n7397, A2 => n7477, B1 => n320, B2 => n7396
                           , ZN => n3296);
   U8342 : OAI22_X1 port map( A1 => n7397, A2 => n7480, B1 => n319, B2 => n7396
                           , ZN => n3297);
   U8343 : OAI22_X1 port map( A1 => n7397, A2 => n7483, B1 => n318, B2 => n7396
                           , ZN => n3298);
   U8344 : OAI22_X1 port map( A1 => n7397, A2 => n7486, B1 => n317, B2 => n7396
                           , ZN => n3299);
   U8345 : OAI22_X1 port map( A1 => n7397, A2 => n7489, B1 => n316, B2 => n7396
                           , ZN => n3300);
   U8346 : OAI22_X1 port map( A1 => n7398, A2 => n7492, B1 => n315, B2 => n7396
                           , ZN => n3301);
   U8347 : OAI22_X1 port map( A1 => n7398, A2 => n7495, B1 => n314, B2 => n7396
                           , ZN => n3302);
   U8348 : OAI22_X1 port map( A1 => n7398, A2 => n7498, B1 => n313, B2 => n7396
                           , ZN => n3303);
   U8349 : OAI22_X1 port map( A1 => n7398, A2 => n7501, B1 => n312, B2 => n7396
                           , ZN => n3304);
   U8350 : OAI22_X1 port map( A1 => n7398, A2 => n7504, B1 => n311, B2 => n7396
                           , ZN => n3305);
   U8351 : OAI22_X1 port map( A1 => n7399, A2 => n7507, B1 => n310, B2 => n7396
                           , ZN => n3306);
   U8352 : OAI22_X1 port map( A1 => n7399, A2 => n7510, B1 => n309, B2 => n7396
                           , ZN => n3307);
   U8353 : OAI22_X1 port map( A1 => n7399, A2 => n7513, B1 => n308, B2 => n5086
                           , ZN => n3308);
   U8354 : OAI22_X1 port map( A1 => n7399, A2 => n7516, B1 => n307, B2 => n5086
                           , ZN => n3309);
   U8355 : OAI22_X1 port map( A1 => n7399, A2 => n7519, B1 => n306, B2 => n5086
                           , ZN => n3310);
   U8356 : OAI22_X1 port map( A1 => n7400, A2 => n7522, B1 => n305, B2 => n7396
                           , ZN => n3311);
   U8357 : OAI22_X1 port map( A1 => n7400, A2 => n7525, B1 => n304, B2 => n7396
                           , ZN => n3312);
   U8358 : OAI22_X1 port map( A1 => n7400, A2 => n7528, B1 => n303, B2 => n7396
                           , ZN => n3313);
   U8359 : OAI22_X1 port map( A1 => n7400, A2 => n7531, B1 => n302, B2 => n7396
                           , ZN => n3314);
   U8360 : OAI22_X1 port map( A1 => n7400, A2 => n7534, B1 => n301, B2 => n7396
                           , ZN => n3315);
   U8361 : OAI22_X1 port map( A1 => n7401, A2 => n7537, B1 => n300, B2 => n7396
                           , ZN => n3316);
   U8362 : OAI22_X1 port map( A1 => n7401, A2 => n7540, B1 => n299, B2 => n7396
                           , ZN => n3317);
   U8363 : OAI22_X1 port map( A1 => n7401, A2 => n7543, B1 => n298, B2 => n7396
                           , ZN => n3318);
   U8364 : OAI22_X1 port map( A1 => n7401, A2 => n7546, B1 => n297, B2 => n7396
                           , ZN => n3319);
   U8365 : OAI22_X1 port map( A1 => n7406, A2 => n7477, B1 => n288, B2 => n7405
                           , ZN => n3328);
   U8366 : OAI22_X1 port map( A1 => n7406, A2 => n7480, B1 => n287, B2 => n7405
                           , ZN => n3329);
   U8367 : OAI22_X1 port map( A1 => n7406, A2 => n7483, B1 => n286, B2 => n7405
                           , ZN => n3330);
   U8368 : OAI22_X1 port map( A1 => n7406, A2 => n7486, B1 => n285, B2 => n7405
                           , ZN => n3331);
   U8369 : OAI22_X1 port map( A1 => n7406, A2 => n7489, B1 => n284, B2 => n7405
                           , ZN => n3332);
   U8370 : OAI22_X1 port map( A1 => n7407, A2 => n7492, B1 => n283, B2 => n7405
                           , ZN => n3333);
   U8371 : OAI22_X1 port map( A1 => n7407, A2 => n7495, B1 => n282, B2 => n7405
                           , ZN => n3334);
   U8372 : OAI22_X1 port map( A1 => n7407, A2 => n7498, B1 => n281, B2 => n7405
                           , ZN => n3335);
   U8373 : OAI22_X1 port map( A1 => n7407, A2 => n7501, B1 => n280, B2 => n7405
                           , ZN => n3336);
   U8374 : OAI22_X1 port map( A1 => n7407, A2 => n7504, B1 => n279, B2 => n7405
                           , ZN => n3337);
   U8375 : OAI22_X1 port map( A1 => n7408, A2 => n7507, B1 => n278, B2 => n7405
                           , ZN => n3338);
   U8376 : OAI22_X1 port map( A1 => n7408, A2 => n7510, B1 => n277, B2 => n7405
                           , ZN => n3339);
   U8377 : OAI22_X1 port map( A1 => n7408, A2 => n7513, B1 => n276, B2 => n5084
                           , ZN => n3340);
   U8378 : OAI22_X1 port map( A1 => n7408, A2 => n7516, B1 => n275, B2 => n5084
                           , ZN => n3341);
   U8379 : OAI22_X1 port map( A1 => n7408, A2 => n7519, B1 => n274, B2 => n5084
                           , ZN => n3342);
   U8380 : OAI22_X1 port map( A1 => n7409, A2 => n7522, B1 => n273, B2 => n7405
                           , ZN => n3343);
   U8381 : OAI22_X1 port map( A1 => n7409, A2 => n7525, B1 => n272, B2 => n7405
                           , ZN => n3344);
   U8382 : OAI22_X1 port map( A1 => n7409, A2 => n7528, B1 => n271, B2 => n7405
                           , ZN => n3345);
   U8383 : OAI22_X1 port map( A1 => n7409, A2 => n7531, B1 => n270, B2 => n7405
                           , ZN => n3346);
   U8384 : OAI22_X1 port map( A1 => n7409, A2 => n7534, B1 => n269, B2 => n7405
                           , ZN => n3347);
   U8385 : OAI22_X1 port map( A1 => n7410, A2 => n7537, B1 => n268, B2 => n7405
                           , ZN => n3348);
   U8386 : OAI22_X1 port map( A1 => n7410, A2 => n7540, B1 => n267, B2 => n7405
                           , ZN => n3349);
   U8387 : OAI22_X1 port map( A1 => n7410, A2 => n7543, B1 => n266, B2 => n7405
                           , ZN => n3350);
   U8388 : OAI22_X1 port map( A1 => n7410, A2 => n7546, B1 => n265, B2 => n7405
                           , ZN => n3351);
   U8389 : OAI22_X1 port map( A1 => n7415, A2 => n7477, B1 => n256, B2 => n7414
                           , ZN => n3360);
   U8390 : OAI22_X1 port map( A1 => n7415, A2 => n7480, B1 => n255, B2 => n7414
                           , ZN => n3361);
   U8391 : OAI22_X1 port map( A1 => n7415, A2 => n7483, B1 => n254, B2 => n7414
                           , ZN => n3362);
   U8392 : OAI22_X1 port map( A1 => n7415, A2 => n7486, B1 => n253, B2 => n7414
                           , ZN => n3363);
   U8393 : OAI22_X1 port map( A1 => n7415, A2 => n7489, B1 => n252, B2 => n7414
                           , ZN => n3364);
   U8394 : OAI22_X1 port map( A1 => n7416, A2 => n7492, B1 => n251, B2 => n7414
                           , ZN => n3365);
   U8395 : OAI22_X1 port map( A1 => n7416, A2 => n7495, B1 => n250, B2 => n7414
                           , ZN => n3366);
   U8396 : OAI22_X1 port map( A1 => n7416, A2 => n7498, B1 => n249, B2 => n7414
                           , ZN => n3367);
   U8397 : OAI22_X1 port map( A1 => n7416, A2 => n7501, B1 => n248, B2 => n7414
                           , ZN => n3368);
   U8398 : OAI22_X1 port map( A1 => n7416, A2 => n7504, B1 => n247, B2 => n7414
                           , ZN => n3369);
   U8399 : OAI22_X1 port map( A1 => n7417, A2 => n7507, B1 => n246, B2 => n7414
                           , ZN => n3370);
   U8400 : OAI22_X1 port map( A1 => n7417, A2 => n7510, B1 => n245, B2 => n7414
                           , ZN => n3371);
   U8401 : OAI22_X1 port map( A1 => n7417, A2 => n7513, B1 => n244, B2 => n5081
                           , ZN => n3372);
   U8402 : OAI22_X1 port map( A1 => n7417, A2 => n7516, B1 => n243, B2 => n5081
                           , ZN => n3373);
   U8403 : OAI22_X1 port map( A1 => n7417, A2 => n7519, B1 => n242, B2 => n5081
                           , ZN => n3374);
   U8404 : OAI22_X1 port map( A1 => n7418, A2 => n7522, B1 => n241, B2 => n7414
                           , ZN => n3375);
   U8405 : OAI22_X1 port map( A1 => n7418, A2 => n7525, B1 => n240, B2 => n7414
                           , ZN => n3376);
   U8406 : OAI22_X1 port map( A1 => n7418, A2 => n7528, B1 => n239, B2 => n7414
                           , ZN => n3377);
   U8407 : OAI22_X1 port map( A1 => n7418, A2 => n7531, B1 => n238, B2 => n7414
                           , ZN => n3378);
   U8408 : OAI22_X1 port map( A1 => n7418, A2 => n7534, B1 => n237, B2 => n7414
                           , ZN => n3379);
   U8409 : OAI22_X1 port map( A1 => n7419, A2 => n7537, B1 => n236, B2 => n7414
                           , ZN => n3380);
   U8410 : OAI22_X1 port map( A1 => n7419, A2 => n7540, B1 => n235, B2 => n7414
                           , ZN => n3381);
   U8411 : OAI22_X1 port map( A1 => n7419, A2 => n7543, B1 => n234, B2 => n7414
                           , ZN => n3382);
   U8412 : OAI22_X1 port map( A1 => n7419, A2 => n7546, B1 => n233, B2 => n7414
                           , ZN => n3383);
   U8413 : OAI22_X1 port map( A1 => n7424, A2 => n7477, B1 => n224, B2 => n7423
                           , ZN => n3392);
   U8414 : OAI22_X1 port map( A1 => n7424, A2 => n7480, B1 => n223, B2 => n7423
                           , ZN => n3393);
   U8415 : OAI22_X1 port map( A1 => n7424, A2 => n7483, B1 => n222, B2 => n7423
                           , ZN => n3394);
   U8416 : OAI22_X1 port map( A1 => n7424, A2 => n7486, B1 => n221, B2 => n7423
                           , ZN => n3395);
   U8417 : OAI22_X1 port map( A1 => n7424, A2 => n7489, B1 => n220, B2 => n7423
                           , ZN => n3396);
   U8418 : OAI22_X1 port map( A1 => n7425, A2 => n7492, B1 => n219, B2 => n7423
                           , ZN => n3397);
   U8419 : OAI22_X1 port map( A1 => n7425, A2 => n7495, B1 => n218, B2 => n7423
                           , ZN => n3398);
   U8420 : OAI22_X1 port map( A1 => n7425, A2 => n7498, B1 => n217, B2 => n7423
                           , ZN => n3399);
   U8421 : OAI22_X1 port map( A1 => n7425, A2 => n7501, B1 => n216, B2 => n7423
                           , ZN => n3400);
   U8422 : OAI22_X1 port map( A1 => n7425, A2 => n7504, B1 => n215, B2 => n7423
                           , ZN => n3401);
   U8423 : OAI22_X1 port map( A1 => n7426, A2 => n7507, B1 => n214, B2 => n7423
                           , ZN => n3402);
   U8424 : OAI22_X1 port map( A1 => n7426, A2 => n7510, B1 => n213, B2 => n7423
                           , ZN => n3403);
   U8425 : OAI22_X1 port map( A1 => n7426, A2 => n7513, B1 => n212, B2 => n5079
                           , ZN => n3404);
   U8426 : OAI22_X1 port map( A1 => n7426, A2 => n7516, B1 => n211, B2 => n5079
                           , ZN => n3405);
   U8427 : OAI22_X1 port map( A1 => n7426, A2 => n7519, B1 => n210, B2 => n5079
                           , ZN => n3406);
   U8428 : OAI22_X1 port map( A1 => n7427, A2 => n7522, B1 => n209, B2 => n7423
                           , ZN => n3407);
   U8429 : OAI22_X1 port map( A1 => n7427, A2 => n7525, B1 => n208, B2 => n7423
                           , ZN => n3408);
   U8430 : OAI22_X1 port map( A1 => n7427, A2 => n7528, B1 => n207, B2 => n7423
                           , ZN => n3409);
   U8431 : OAI22_X1 port map( A1 => n7427, A2 => n7531, B1 => n206, B2 => n7423
                           , ZN => n3410);
   U8432 : OAI22_X1 port map( A1 => n7427, A2 => n7534, B1 => n205, B2 => n7423
                           , ZN => n3411);
   U8433 : OAI22_X1 port map( A1 => n7428, A2 => n7537, B1 => n204, B2 => n7423
                           , ZN => n3412);
   U8434 : OAI22_X1 port map( A1 => n7428, A2 => n7540, B1 => n203, B2 => n7423
                           , ZN => n3413);
   U8435 : OAI22_X1 port map( A1 => n7428, A2 => n7543, B1 => n202, B2 => n7423
                           , ZN => n3414);
   U8436 : OAI22_X1 port map( A1 => n7428, A2 => n7546, B1 => n201, B2 => n7423
                           , ZN => n3415);
   U8437 : OAI22_X1 port map( A1 => n7469, A2 => n7477, B1 => n64, B2 => n7468,
                           ZN => n3552);
   U8438 : OAI22_X1 port map( A1 => n7469, A2 => n7480, B1 => n63, B2 => n7468,
                           ZN => n3553);
   U8439 : OAI22_X1 port map( A1 => n7469, A2 => n7483, B1 => n62, B2 => n7468,
                           ZN => n3554);
   U8440 : OAI22_X1 port map( A1 => n7469, A2 => n7486, B1 => n61, B2 => n7468,
                           ZN => n3555);
   U8441 : OAI22_X1 port map( A1 => n7469, A2 => n7489, B1 => n60, B2 => n7468,
                           ZN => n3556);
   U8442 : OAI22_X1 port map( A1 => n7470, A2 => n7492, B1 => n59, B2 => n7468,
                           ZN => n3557);
   U8443 : OAI22_X1 port map( A1 => n7470, A2 => n7495, B1 => n58, B2 => n7468,
                           ZN => n3558);
   U8444 : OAI22_X1 port map( A1 => n7470, A2 => n7498, B1 => n57, B2 => n7468,
                           ZN => n3559);
   U8445 : OAI22_X1 port map( A1 => n7470, A2 => n7501, B1 => n56, B2 => n7468,
                           ZN => n3560);
   U8446 : OAI22_X1 port map( A1 => n7470, A2 => n7504, B1 => n55, B2 => n7468,
                           ZN => n3561);
   U8447 : OAI22_X1 port map( A1 => n7471, A2 => n7507, B1 => n54, B2 => n7468,
                           ZN => n3562);
   U8448 : OAI22_X1 port map( A1 => n7471, A2 => n7510, B1 => n53, B2 => n7468,
                           ZN => n3563);
   U8449 : OAI22_X1 port map( A1 => n7471, A2 => n7513, B1 => n52, B2 => n5069,
                           ZN => n3564);
   U8450 : OAI22_X1 port map( A1 => n7471, A2 => n7516, B1 => n51, B2 => n5069,
                           ZN => n3565);
   U8451 : OAI22_X1 port map( A1 => n7471, A2 => n7519, B1 => n50, B2 => n5069,
                           ZN => n3566);
   U8452 : OAI22_X1 port map( A1 => n7472, A2 => n7522, B1 => n49, B2 => n7468,
                           ZN => n3567);
   U8453 : OAI22_X1 port map( A1 => n7472, A2 => n7525, B1 => n48, B2 => n7468,
                           ZN => n3568);
   U8454 : OAI22_X1 port map( A1 => n7472, A2 => n7528, B1 => n47, B2 => n7468,
                           ZN => n3569);
   U8455 : OAI22_X1 port map( A1 => n7472, A2 => n7531, B1 => n46, B2 => n7468,
                           ZN => n3570);
   U8456 : OAI22_X1 port map( A1 => n7472, A2 => n7534, B1 => n45, B2 => n7468,
                           ZN => n3571);
   U8457 : OAI22_X1 port map( A1 => n7473, A2 => n7537, B1 => n44, B2 => n7468,
                           ZN => n3572);
   U8458 : OAI22_X1 port map( A1 => n7473, A2 => n7540, B1 => n43, B2 => n7468,
                           ZN => n3573);
   U8459 : OAI22_X1 port map( A1 => n7473, A2 => n7543, B1 => n42, B2 => n7468,
                           ZN => n3574);
   U8460 : OAI22_X1 port map( A1 => n7473, A2 => n7546, B1 => n41, B2 => n7468,
                           ZN => n3575);
   U8461 : OAI22_X1 port map( A1 => n7571, A2 => n7477, B1 => n32, B2 => n7570,
                           ZN => n3584);
   U8462 : OAI22_X1 port map( A1 => n7571, A2 => n7480, B1 => n31, B2 => n7570,
                           ZN => n3585);
   U8463 : OAI22_X1 port map( A1 => n7571, A2 => n7483, B1 => n30, B2 => n7570,
                           ZN => n3586);
   U8464 : OAI22_X1 port map( A1 => n7571, A2 => n7486, B1 => n29, B2 => n7570,
                           ZN => n3587);
   U8465 : OAI22_X1 port map( A1 => n7571, A2 => n7489, B1 => n28, B2 => n7570,
                           ZN => n3588);
   U8466 : OAI22_X1 port map( A1 => n7572, A2 => n7492, B1 => n27, B2 => n7570,
                           ZN => n3589);
   U8467 : OAI22_X1 port map( A1 => n7572, A2 => n7495, B1 => n26, B2 => n7570,
                           ZN => n3590);
   U8468 : OAI22_X1 port map( A1 => n7572, A2 => n7498, B1 => n25, B2 => n7570,
                           ZN => n3591);
   U8469 : OAI22_X1 port map( A1 => n7572, A2 => n7501, B1 => n24, B2 => n7570,
                           ZN => n3592);
   U8470 : OAI22_X1 port map( A1 => n7572, A2 => n7504, B1 => n23, B2 => n7570,
                           ZN => n3593);
   U8471 : OAI22_X1 port map( A1 => n7573, A2 => n7507, B1 => n22, B2 => n7570,
                           ZN => n3594);
   U8472 : OAI22_X1 port map( A1 => n7573, A2 => n7510, B1 => n21, B2 => n7570,
                           ZN => n3595);
   U8473 : OAI22_X1 port map( A1 => n7573, A2 => n7513, B1 => n20, B2 => n5035,
                           ZN => n3596);
   U8474 : OAI22_X1 port map( A1 => n7573, A2 => n7516, B1 => n19, B2 => n5035,
                           ZN => n3597);
   U8475 : OAI22_X1 port map( A1 => n7573, A2 => n7519, B1 => n18, B2 => n5035,
                           ZN => n3598);
   U8476 : OAI22_X1 port map( A1 => n7574, A2 => n7522, B1 => n17, B2 => n7570,
                           ZN => n3599);
   U8477 : OAI22_X1 port map( A1 => n7574, A2 => n7525, B1 => n16, B2 => n7570,
                           ZN => n3600);
   U8478 : OAI22_X1 port map( A1 => n7574, A2 => n7528, B1 => n15, B2 => n7570,
                           ZN => n3601);
   U8479 : OAI22_X1 port map( A1 => n7574, A2 => n7531, B1 => n14, B2 => n7570,
                           ZN => n3602);
   U8480 : OAI22_X1 port map( A1 => n7574, A2 => n7534, B1 => n13, B2 => n7570,
                           ZN => n3603);
   U8481 : OAI22_X1 port map( A1 => n7575, A2 => n7537, B1 => n12, B2 => n7570,
                           ZN => n3604);
   U8482 : OAI22_X1 port map( A1 => n7575, A2 => n7540, B1 => n11, B2 => n7570,
                           ZN => n3605);
   U8483 : OAI22_X1 port map( A1 => n7575, A2 => n7543, B1 => n10, B2 => n7570,
                           ZN => n3606);
   U8484 : OAI22_X1 port map( A1 => n7575, A2 => n7546, B1 => n9, B2 => n7570, 
                           ZN => n3607);
   U8485 : OAI21_X1 port map( B1 => n6937, B2 => n7090, A => n6253, ZN => n2535
                           );
   U8486 : OAI21_X1 port map( B1 => n6254, B2 => n6255, A => n7092, ZN => n6253
                           );
   U8487 : NAND4_X1 port map( A1 => n6264, A2 => n6265, A3 => n6266, A4 => 
                           n6267, ZN => n6254);
   U8488 : NAND4_X1 port map( A1 => n6256, A2 => n6257, A3 => n6258, A4 => 
                           n6259, ZN => n6255);
   U8489 : OAI21_X1 port map( B1 => n6970, B2 => n7090, A => n6215, ZN => n2537
                           );
   U8490 : OAI21_X1 port map( B1 => n6216, B2 => n6217, A => n7092, ZN => n6215
                           );
   U8491 : NAND4_X1 port map( A1 => n6226, A2 => n6227, A3 => n6228, A4 => 
                           n6229, ZN => n6216);
   U8492 : NAND4_X1 port map( A1 => n6218, A2 => n6219, A3 => n6220, A4 => 
                           n6221, ZN => n6217);
   U8493 : OAI21_X1 port map( B1 => n6971, B2 => n7090, A => n6196, ZN => n2538
                           );
   U8494 : OAI21_X1 port map( B1 => n6197, B2 => n6198, A => n7091, ZN => n6196
                           );
   U8495 : NAND4_X1 port map( A1 => n6207, A2 => n6208, A3 => n6209, A4 => 
                           n6210, ZN => n6197);
   U8496 : NAND4_X1 port map( A1 => n6199, A2 => n6200, A3 => n6201, A4 => 
                           n6202, ZN => n6198);
   U8497 : OAI21_X1 port map( B1 => n6972, B2 => n7090, A => n6177, ZN => n2539
                           );
   U8498 : OAI21_X1 port map( B1 => n6178, B2 => n6179, A => n7091, ZN => n6177
                           );
   U8499 : NAND4_X1 port map( A1 => n6188, A2 => n6189, A3 => n6190, A4 => 
                           n6191, ZN => n6178);
   U8500 : NAND4_X1 port map( A1 => n6180, A2 => n6181, A3 => n6182, A4 => 
                           n6183, ZN => n6179);
   U8501 : OAI21_X1 port map( B1 => n6973, B2 => n7090, A => n6158, ZN => n2540
                           );
   U8502 : OAI21_X1 port map( B1 => n6159, B2 => n6160, A => n7092, ZN => n6158
                           );
   U8503 : NAND4_X1 port map( A1 => n6169, A2 => n6170, A3 => n6171, A4 => 
                           n6172, ZN => n6159);
   U8504 : NAND4_X1 port map( A1 => n6161, A2 => n6162, A3 => n6163, A4 => 
                           n6164, ZN => n6160);
   U8505 : OAI21_X1 port map( B1 => n6974, B2 => n7090, A => n6139, ZN => n2541
                           );
   U8506 : OAI21_X1 port map( B1 => n6140, B2 => n6141, A => n7091, ZN => n6139
                           );
   U8507 : NAND4_X1 port map( A1 => n6150, A2 => n6151, A3 => n6152, A4 => 
                           n6153, ZN => n6140);
   U8508 : NAND4_X1 port map( A1 => n6142, A2 => n6143, A3 => n6144, A4 => 
                           n6145, ZN => n6141);
   U8509 : OAI21_X1 port map( B1 => n6975, B2 => n7090, A => n6120, ZN => n2542
                           );
   U8510 : OAI21_X1 port map( B1 => n6121, B2 => n6122, A => n7091, ZN => n6120
                           );
   U8511 : NAND4_X1 port map( A1 => n6131, A2 => n6132, A3 => n6133, A4 => 
                           n6134, ZN => n6121);
   U8512 : NAND4_X1 port map( A1 => n6123, A2 => n6124, A3 => n6125, A4 => 
                           n6126, ZN => n6122);
   U8513 : OAI21_X1 port map( B1 => n6976, B2 => n7090, A => n6101, ZN => n2543
                           );
   U8514 : OAI21_X1 port map( B1 => n6102, B2 => n6103, A => n7092, ZN => n6101
                           );
   U8515 : NAND4_X1 port map( A1 => n6112, A2 => n6113, A3 => n6114, A4 => 
                           n6115, ZN => n6102);
   U8516 : NAND4_X1 port map( A1 => n6104, A2 => n6105, A3 => n6106, A4 => 
                           n6107, ZN => n6103);
   U8517 : OAI21_X1 port map( B1 => n6977, B2 => n7090, A => n6082, ZN => n2544
                           );
   U8518 : OAI21_X1 port map( B1 => n6083, B2 => n6084, A => n7092, ZN => n6082
                           );
   U8519 : NAND4_X1 port map( A1 => n6093, A2 => n6094, A3 => n6095, A4 => 
                           n6096, ZN => n6083);
   U8520 : NAND4_X1 port map( A1 => n6085, A2 => n6086, A3 => n6087, A4 => 
                           n6088, ZN => n6084);
   U8521 : OAI21_X1 port map( B1 => n6978, B2 => n7090, A => n6063, ZN => n2545
                           );
   U8522 : OAI21_X1 port map( B1 => n6064, B2 => n6065, A => n7092, ZN => n6063
                           );
   U8523 : NAND4_X1 port map( A1 => n6074, A2 => n6075, A3 => n6076, A4 => 
                           n6077, ZN => n6064);
   U8524 : NAND4_X1 port map( A1 => n6066, A2 => n6067, A3 => n6068, A4 => 
                           n6069, ZN => n6065);
   U8525 : OAI21_X1 port map( B1 => n6979, B2 => n7090, A => n6044, ZN => n2546
                           );
   U8526 : OAI21_X1 port map( B1 => n6045, B2 => n6046, A => n7092, ZN => n6044
                           );
   U8527 : NAND4_X1 port map( A1 => n6055, A2 => n6056, A3 => n6057, A4 => 
                           n6058, ZN => n6045);
   U8528 : NAND4_X1 port map( A1 => n6047, A2 => n6048, A3 => n6049, A4 => 
                           n6050, ZN => n6046);
   U8529 : OAI21_X1 port map( B1 => n6929, B2 => n7090, A => n5765, ZN => n2559
                           );
   U8530 : OAI21_X1 port map( B1 => n5766, B2 => n5767, A => n7094, ZN => n5765
                           );
   U8531 : NAND4_X1 port map( A1 => n5792, A2 => n5793, A3 => n5794, A4 => 
                           n5795, ZN => n5766);
   U8532 : NAND4_X1 port map( A1 => n5768, A2 => n5769, A3 => n5770, A4 => 
                           n5771, ZN => n5767);
   U8533 : OAI21_X1 port map( B1 => n6945, B2 => n7192, A => n5600, ZN => n2574
                           );
   U8534 : OAI21_X1 port map( B1 => n5601, B2 => n5602, A => n7194, ZN => n5600
                           );
   U8535 : NAND4_X1 port map( A1 => n5611, A2 => n5612, A3 => n5613, A4 => 
                           n5614, ZN => n5601);
   U8536 : NAND4_X1 port map( A1 => n5603, A2 => n5604, A3 => n5605, A4 => 
                           n5606, ZN => n5602);
   U8537 : OAI21_X1 port map( B1 => n6947, B2 => n7192, A => n5562, ZN => n2578
                           );
   U8538 : OAI21_X1 port map( B1 => n5563, B2 => n5564, A => n7194, ZN => n5562
                           );
   U8539 : NAND4_X1 port map( A1 => n5573, A2 => n5574, A3 => n5575, A4 => 
                           n5576, ZN => n5563);
   U8540 : NAND4_X1 port map( A1 => n5565, A2 => n5566, A3 => n5567, A4 => 
                           n5568, ZN => n5564);
   U8541 : OAI21_X1 port map( B1 => n6948, B2 => n7192, A => n5543, ZN => n2580
                           );
   U8542 : OAI21_X1 port map( B1 => n5544, B2 => n5545, A => n7193, ZN => n5543
                           );
   U8543 : NAND4_X1 port map( A1 => n5554, A2 => n5555, A3 => n5556, A4 => 
                           n5557, ZN => n5544);
   U8544 : NAND4_X1 port map( A1 => n5546, A2 => n5547, A3 => n5548, A4 => 
                           n5549, ZN => n5545);
   U8545 : OAI21_X1 port map( B1 => n6949, B2 => n7192, A => n5524, ZN => n2582
                           );
   U8546 : OAI21_X1 port map( B1 => n5525, B2 => n5526, A => n7193, ZN => n5524
                           );
   U8547 : NAND4_X1 port map( A1 => n5535, A2 => n5536, A3 => n5537, A4 => 
                           n5538, ZN => n5525);
   U8548 : NAND4_X1 port map( A1 => n5527, A2 => n5528, A3 => n5529, A4 => 
                           n5530, ZN => n5526);
   U8549 : OAI21_X1 port map( B1 => n6950, B2 => n7192, A => n5505, ZN => n2584
                           );
   U8550 : OAI21_X1 port map( B1 => n5506, B2 => n5507, A => n7194, ZN => n5505
                           );
   U8551 : NAND4_X1 port map( A1 => n5516, A2 => n5517, A3 => n5518, A4 => 
                           n5519, ZN => n5506);
   U8552 : NAND4_X1 port map( A1 => n5508, A2 => n5509, A3 => n5510, A4 => 
                           n5511, ZN => n5507);
   U8553 : OAI21_X1 port map( B1 => n6951, B2 => n7192, A => n5486, ZN => n2586
                           );
   U8554 : OAI21_X1 port map( B1 => n5487, B2 => n5488, A => n7193, ZN => n5486
                           );
   U8555 : NAND4_X1 port map( A1 => n5497, A2 => n5498, A3 => n5499, A4 => 
                           n5500, ZN => n5487);
   U8556 : NAND4_X1 port map( A1 => n5489, A2 => n5490, A3 => n5491, A4 => 
                           n5492, ZN => n5488);
   U8557 : OAI21_X1 port map( B1 => n6952, B2 => n7192, A => n5467, ZN => n2588
                           );
   U8558 : OAI21_X1 port map( B1 => n5468, B2 => n5469, A => n7193, ZN => n5467
                           );
   U8559 : NAND4_X1 port map( A1 => n5478, A2 => n5479, A3 => n5480, A4 => 
                           n5481, ZN => n5468);
   U8560 : NAND4_X1 port map( A1 => n5470, A2 => n5471, A3 => n5472, A4 => 
                           n5473, ZN => n5469);
   U8561 : OAI21_X1 port map( B1 => n6953, B2 => n7192, A => n5448, ZN => n2590
                           );
   U8562 : OAI21_X1 port map( B1 => n5449, B2 => n5450, A => n7194, ZN => n5448
                           );
   U8563 : NAND4_X1 port map( A1 => n5459, A2 => n5460, A3 => n5461, A4 => 
                           n5462, ZN => n5449);
   U8564 : NAND4_X1 port map( A1 => n5451, A2 => n5452, A3 => n5453, A4 => 
                           n5454, ZN => n5450);
   U8565 : OAI21_X1 port map( B1 => n6954, B2 => n7192, A => n5429, ZN => n2592
                           );
   U8566 : OAI21_X1 port map( B1 => n5430, B2 => n5431, A => n7194, ZN => n5429
                           );
   U8567 : NAND4_X1 port map( A1 => n5440, A2 => n5441, A3 => n5442, A4 => 
                           n5443, ZN => n5430);
   U8568 : NAND4_X1 port map( A1 => n5432, A2 => n5433, A3 => n5434, A4 => 
                           n5435, ZN => n5431);
   U8569 : OAI21_X1 port map( B1 => n6955, B2 => n7192, A => n5410, ZN => n2594
                           );
   U8570 : OAI21_X1 port map( B1 => n5411, B2 => n5412, A => n7194, ZN => n5410
                           );
   U8571 : NAND4_X1 port map( A1 => n5421, A2 => n5422, A3 => n5423, A4 => 
                           n5424, ZN => n5411);
   U8572 : NAND4_X1 port map( A1 => n5413, A2 => n5414, A3 => n5415, A4 => 
                           n5416, ZN => n5412);
   U8573 : OAI21_X1 port map( B1 => n6956, B2 => n7192, A => n5391, ZN => n2596
                           );
   U8574 : OAI21_X1 port map( B1 => n5392, B2 => n5393, A => n7194, ZN => n5391
                           );
   U8575 : NAND4_X1 port map( A1 => n5402, A2 => n5403, A3 => n5404, A4 => 
                           n5405, ZN => n5392);
   U8576 : NAND4_X1 port map( A1 => n5394, A2 => n5395, A3 => n5396, A4 => 
                           n5397, ZN => n5393);
   U8577 : OAI21_X1 port map( B1 => n6992, B2 => n7192, A => n5112, ZN => n2622
                           );
   U8578 : OAI21_X1 port map( B1 => n5113, B2 => n5114, A => n7196, ZN => n5112
                           );
   U8579 : NAND4_X1 port map( A1 => n5139, A2 => n5140, A3 => n5141, A4 => 
                           n5142, ZN => n5113);
   U8580 : NAND4_X1 port map( A1 => n5115, A2 => n5116, A3 => n5117, A4 => 
                           n5118, ZN => n5114);
   U8581 : OAI21_X1 port map( B1 => n6930, B2 => n7091, A => n6386, ZN => n2528
                           );
   U8582 : OAI21_X1 port map( B1 => n6387, B2 => n6388, A => n7094, ZN => n6386
                           );
   U8583 : NAND4_X1 port map( A1 => n6407, A2 => n6408, A3 => n6409, A4 => 
                           n6410, ZN => n6387);
   U8584 : NAND4_X1 port map( A1 => n6389, A2 => n6390, A3 => n6391, A4 => 
                           n6392, ZN => n6388);
   U8585 : OAI21_X1 port map( B1 => n6931, B2 => n7091, A => n6367, ZN => n2529
                           );
   U8586 : OAI21_X1 port map( B1 => n6368, B2 => n6369, A => n7094, ZN => n6367
                           );
   U8587 : NAND4_X1 port map( A1 => n6378, A2 => n6379, A3 => n6380, A4 => 
                           n6381, ZN => n6368);
   U8588 : NAND4_X1 port map( A1 => n6370, A2 => n6371, A3 => n6372, A4 => 
                           n6373, ZN => n6369);
   U8589 : OAI21_X1 port map( B1 => n6932, B2 => n7091, A => n6348, ZN => n2530
                           );
   U8590 : OAI21_X1 port map( B1 => n6349, B2 => n6350, A => n7093, ZN => n6348
                           );
   U8591 : NAND4_X1 port map( A1 => n6359, A2 => n6360, A3 => n6361, A4 => 
                           n6362, ZN => n6349);
   U8592 : NAND4_X1 port map( A1 => n6351, A2 => n6352, A3 => n6353, A4 => 
                           n6354, ZN => n6350);
   U8593 : OAI21_X1 port map( B1 => n6933, B2 => n7091, A => n6329, ZN => n2531
                           );
   U8594 : OAI21_X1 port map( B1 => n6330, B2 => n6331, A => n7093, ZN => n6329
                           );
   U8595 : NAND4_X1 port map( A1 => n6340, A2 => n6341, A3 => n6342, A4 => 
                           n6343, ZN => n6330);
   U8596 : NAND4_X1 port map( A1 => n6332, A2 => n6333, A3 => n6334, A4 => 
                           n6335, ZN => n6331);
   U8597 : OAI21_X1 port map( B1 => n6934, B2 => n7091, A => n6310, ZN => n2532
                           );
   U8598 : OAI21_X1 port map( B1 => n6311, B2 => n6312, A => n7093, ZN => n6310
                           );
   U8599 : NAND4_X1 port map( A1 => n6321, A2 => n6322, A3 => n6323, A4 => 
                           n6324, ZN => n6311);
   U8600 : NAND4_X1 port map( A1 => n6313, A2 => n6314, A3 => n6315, A4 => 
                           n6316, ZN => n6312);
   U8601 : OAI21_X1 port map( B1 => n6935, B2 => n7091, A => n6291, ZN => n2533
                           );
   U8602 : OAI21_X1 port map( B1 => n6292, B2 => n6293, A => n7092, ZN => n6291
                           );
   U8603 : NAND4_X1 port map( A1 => n6302, A2 => n6303, A3 => n6304, A4 => 
                           n6305, ZN => n6292);
   U8604 : NAND4_X1 port map( A1 => n6294, A2 => n6295, A3 => n6296, A4 => 
                           n6297, ZN => n6293);
   U8605 : OAI21_X1 port map( B1 => n6936, B2 => n7091, A => n6272, ZN => n2534
                           );
   U8606 : OAI21_X1 port map( B1 => n6273, B2 => n6274, A => n7093, ZN => n6272
                           );
   U8607 : NAND4_X1 port map( A1 => n6283, A2 => n6284, A3 => n6285, A4 => 
                           n6286, ZN => n6273);
   U8608 : NAND4_X1 port map( A1 => n6275, A2 => n6276, A3 => n6277, A4 => 
                           n6278, ZN => n6274);
   U8609 : OAI21_X1 port map( B1 => n6969, B2 => n7091, A => n6234, ZN => n2536
                           );
   U8610 : OAI21_X1 port map( B1 => n6235, B2 => n6236, A => n7092, ZN => n6234
                           );
   U8611 : NAND4_X1 port map( A1 => n6245, A2 => n6246, A3 => n6247, A4 => 
                           n6248, ZN => n6235);
   U8612 : NAND4_X1 port map( A1 => n6237, A2 => n6238, A3 => n6239, A4 => 
                           n6240, ZN => n6236);
   U8613 : OAI21_X1 port map( B1 => n6938, B2 => n7193, A => n5733, ZN => n2560
                           );
   U8614 : OAI21_X1 port map( B1 => n5734, B2 => n5735, A => n7196, ZN => n5733
                           );
   U8615 : NAND4_X1 port map( A1 => n5754, A2 => n5755, A3 => n5756, A4 => 
                           n5757, ZN => n5734);
   U8616 : NAND4_X1 port map( A1 => n5736, A2 => n5737, A3 => n5738, A4 => 
                           n5739, ZN => n5735);
   U8617 : OAI21_X1 port map( B1 => n6939, B2 => n7193, A => n5714, ZN => n2562
                           );
   U8618 : OAI21_X1 port map( B1 => n5715, B2 => n5716, A => n7196, ZN => n5714
                           );
   U8619 : NAND4_X1 port map( A1 => n5725, A2 => n5726, A3 => n5727, A4 => 
                           n5728, ZN => n5715);
   U8620 : NAND4_X1 port map( A1 => n5717, A2 => n5718, A3 => n5719, A4 => 
                           n5720, ZN => n5716);
   U8621 : OAI21_X1 port map( B1 => n6940, B2 => n7193, A => n5695, ZN => n2564
                           );
   U8622 : OAI21_X1 port map( B1 => n5696, B2 => n5697, A => n7195, ZN => n5695
                           );
   U8623 : NAND4_X1 port map( A1 => n5706, A2 => n5707, A3 => n5708, A4 => 
                           n5709, ZN => n5696);
   U8624 : NAND4_X1 port map( A1 => n5698, A2 => n5699, A3 => n5700, A4 => 
                           n5701, ZN => n5697);
   U8625 : OAI21_X1 port map( B1 => n6941, B2 => n7193, A => n5676, ZN => n2566
                           );
   U8626 : OAI21_X1 port map( B1 => n5677, B2 => n5678, A => n7195, ZN => n5676
                           );
   U8627 : NAND4_X1 port map( A1 => n5687, A2 => n5688, A3 => n5689, A4 => 
                           n5690, ZN => n5677);
   U8628 : NAND4_X1 port map( A1 => n5679, A2 => n5680, A3 => n5681, A4 => 
                           n5682, ZN => n5678);
   U8629 : OAI21_X1 port map( B1 => n6942, B2 => n7193, A => n5657, ZN => n2568
                           );
   U8630 : OAI21_X1 port map( B1 => n5658, B2 => n5659, A => n7195, ZN => n5657
                           );
   U8631 : NAND4_X1 port map( A1 => n5668, A2 => n5669, A3 => n5670, A4 => 
                           n5671, ZN => n5658);
   U8632 : NAND4_X1 port map( A1 => n5660, A2 => n5661, A3 => n5662, A4 => 
                           n5663, ZN => n5659);
   U8633 : OAI21_X1 port map( B1 => n6943, B2 => n7193, A => n5638, ZN => n2570
                           );
   U8634 : OAI21_X1 port map( B1 => n5639, B2 => n5640, A => n7194, ZN => n5638
                           );
   U8635 : NAND4_X1 port map( A1 => n5649, A2 => n5650, A3 => n5651, A4 => 
                           n5652, ZN => n5639);
   U8636 : NAND4_X1 port map( A1 => n5641, A2 => n5642, A3 => n5643, A4 => 
                           n5644, ZN => n5640);
   U8637 : OAI21_X1 port map( B1 => n6944, B2 => n7193, A => n5619, ZN => n2572
                           );
   U8638 : OAI21_X1 port map( B1 => n5620, B2 => n5621, A => n7195, ZN => n5619
                           );
   U8639 : NAND4_X1 port map( A1 => n5630, A2 => n5631, A3 => n5632, A4 => 
                           n5633, ZN => n5620);
   U8640 : NAND4_X1 port map( A1 => n5622, A2 => n5623, A3 => n5624, A4 => 
                           n5625, ZN => n5621);
   U8641 : OAI21_X1 port map( B1 => n6946, B2 => n7193, A => n5581, ZN => n2576
                           );
   U8642 : OAI21_X1 port map( B1 => n5582, B2 => n5583, A => n7194, ZN => n5581
                           );
   U8643 : NAND4_X1 port map( A1 => n5592, A2 => n5593, A3 => n5594, A4 => 
                           n5595, ZN => n5582);
   U8644 : NAND4_X1 port map( A1 => n5584, A2 => n5585, A3 => n5586, A4 => 
                           n5587, ZN => n5583);
   U8645 : OAI21_X1 port map( B1 => n6980, B2 => n7089, A => n6025, ZN => n2547
                           );
   U8646 : OAI21_X1 port map( B1 => n6026, B2 => n6027, A => n7092, ZN => n6025
                           );
   U8647 : NAND4_X1 port map( A1 => n6036, A2 => n6037, A3 => n6038, A4 => 
                           n6039, ZN => n6026);
   U8648 : NAND4_X1 port map( A1 => n6028, A2 => n6029, A3 => n6030, A4 => 
                           n6031, ZN => n6027);
   U8649 : OAI21_X1 port map( B1 => n6981, B2 => n7089, A => n6006, ZN => n2548
                           );
   U8650 : OAI21_X1 port map( B1 => n6007, B2 => n6008, A => n7092, ZN => n6006
                           );
   U8651 : NAND4_X1 port map( A1 => n6017, A2 => n6018, A3 => n6019, A4 => 
                           n6020, ZN => n6007);
   U8652 : NAND4_X1 port map( A1 => n6009, A2 => n6010, A3 => n6011, A4 => 
                           n6012, ZN => n6008);
   U8653 : OAI21_X1 port map( B1 => n6982, B2 => n7089, A => n5987, ZN => n2549
                           );
   U8654 : OAI21_X1 port map( B1 => n5988, B2 => n5989, A => n7093, ZN => n5987
                           );
   U8655 : NAND4_X1 port map( A1 => n5998, A2 => n5999, A3 => n6000, A4 => 
                           n6001, ZN => n5988);
   U8656 : NAND4_X1 port map( A1 => n5990, A2 => n5991, A3 => n5992, A4 => 
                           n5993, ZN => n5989);
   U8657 : OAI21_X1 port map( B1 => n6983, B2 => n7089, A => n5968, ZN => n2550
                           );
   U8658 : OAI21_X1 port map( B1 => n5969, B2 => n5970, A => n7092, ZN => n5968
                           );
   U8659 : NAND4_X1 port map( A1 => n5979, A2 => n5980, A3 => n5981, A4 => 
                           n5982, ZN => n5969);
   U8660 : NAND4_X1 port map( A1 => n5971, A2 => n5972, A3 => n5973, A4 => 
                           n5974, ZN => n5970);
   U8661 : OAI21_X1 port map( B1 => n6984, B2 => n7089, A => n5949, ZN => n2551
                           );
   U8662 : OAI21_X1 port map( B1 => n5950, B2 => n5951, A => n7093, ZN => n5949
                           );
   U8663 : NAND4_X1 port map( A1 => n5960, A2 => n5961, A3 => n5962, A4 => 
                           n5963, ZN => n5950);
   U8664 : NAND4_X1 port map( A1 => n5952, A2 => n5953, A3 => n5954, A4 => 
                           n5955, ZN => n5951);
   U8665 : OAI21_X1 port map( B1 => n6985, B2 => n7089, A => n5930, ZN => n2552
                           );
   U8666 : OAI21_X1 port map( B1 => n5931, B2 => n5932, A => n7093, ZN => n5930
                           );
   U8667 : NAND4_X1 port map( A1 => n5941, A2 => n5942, A3 => n5943, A4 => 
                           n5944, ZN => n5931);
   U8668 : NAND4_X1 port map( A1 => n5933, A2 => n5934, A3 => n5935, A4 => 
                           n5936, ZN => n5932);
   U8669 : OAI21_X1 port map( B1 => n6986, B2 => n7089, A => n5911, ZN => n2553
                           );
   U8670 : OAI21_X1 port map( B1 => n5912, B2 => n5913, A => n7093, ZN => n5911
                           );
   U8671 : NAND4_X1 port map( A1 => n5922, A2 => n5923, A3 => n5924, A4 => 
                           n5925, ZN => n5912);
   U8672 : NAND4_X1 port map( A1 => n5914, A2 => n5915, A3 => n5916, A4 => 
                           n5917, ZN => n5913);
   U8673 : OAI21_X1 port map( B1 => n6987, B2 => n7089, A => n5892, ZN => n2554
                           );
   U8674 : OAI21_X1 port map( B1 => n5893, B2 => n5894, A => n7093, ZN => n5892
                           );
   U8675 : NAND4_X1 port map( A1 => n5903, A2 => n5904, A3 => n5905, A4 => 
                           n5906, ZN => n5893);
   U8676 : NAND4_X1 port map( A1 => n5895, A2 => n5896, A3 => n5897, A4 => 
                           n5898, ZN => n5894);
   U8677 : OAI21_X1 port map( B1 => n6988, B2 => n7089, A => n5873, ZN => n2555
                           );
   U8678 : OAI21_X1 port map( B1 => n5874, B2 => n5875, A => n7093, ZN => n5873
                           );
   U8679 : NAND4_X1 port map( A1 => n5884, A2 => n5885, A3 => n5886, A4 => 
                           n5887, ZN => n5874);
   U8680 : NAND4_X1 port map( A1 => n5876, A2 => n5877, A3 => n5878, A4 => 
                           n5879, ZN => n5875);
   U8681 : OAI21_X1 port map( B1 => n6989, B2 => n7089, A => n5854, ZN => n2556
                           );
   U8682 : OAI21_X1 port map( B1 => n5855, B2 => n5856, A => n7093, ZN => n5854
                           );
   U8683 : NAND4_X1 port map( A1 => n5865, A2 => n5866, A3 => n5867, A4 => 
                           n5868, ZN => n5855);
   U8684 : NAND4_X1 port map( A1 => n5857, A2 => n5858, A3 => n5859, A4 => 
                           n5860, ZN => n5856);
   U8685 : OAI21_X1 port map( B1 => n6990, B2 => n7089, A => n5835, ZN => n2557
                           );
   U8686 : OAI21_X1 port map( B1 => n5836, B2 => n5837, A => n7093, ZN => n5835
                           );
   U8687 : NAND4_X1 port map( A1 => n5846, A2 => n5847, A3 => n5848, A4 => 
                           n5849, ZN => n5836);
   U8688 : NAND4_X1 port map( A1 => n5838, A2 => n5839, A3 => n5840, A4 => 
                           n5841, ZN => n5837);
   U8689 : OAI21_X1 port map( B1 => n6991, B2 => n7089, A => n5816, ZN => n2558
                           );
   U8690 : OAI21_X1 port map( B1 => n5817, B2 => n5818, A => n7094, ZN => n5816
                           );
   U8691 : NAND4_X1 port map( A1 => n5827, A2 => n5828, A3 => n5829, A4 => 
                           n5830, ZN => n5817);
   U8692 : NAND4_X1 port map( A1 => n5819, A2 => n5820, A3 => n5821, A4 => 
                           n5822, ZN => n5818);
   U8693 : OAI21_X1 port map( B1 => n6957, B2 => n7191, A => n5372, ZN => n2598
                           );
   U8694 : OAI21_X1 port map( B1 => n5373, B2 => n5374, A => n7194, ZN => n5372
                           );
   U8695 : NAND4_X1 port map( A1 => n5383, A2 => n5384, A3 => n5385, A4 => 
                           n5386, ZN => n5373);
   U8696 : NAND4_X1 port map( A1 => n5375, A2 => n5376, A3 => n5377, A4 => 
                           n5378, ZN => n5374);
   U8697 : OAI21_X1 port map( B1 => n6958, B2 => n7191, A => n5353, ZN => n2600
                           );
   U8698 : OAI21_X1 port map( B1 => n5354, B2 => n5355, A => n7194, ZN => n5353
                           );
   U8699 : NAND4_X1 port map( A1 => n5364, A2 => n5365, A3 => n5366, A4 => 
                           n5367, ZN => n5354);
   U8700 : NAND4_X1 port map( A1 => n5356, A2 => n5357, A3 => n5358, A4 => 
                           n5359, ZN => n5355);
   U8701 : OAI21_X1 port map( B1 => n6959, B2 => n7191, A => n5334, ZN => n2602
                           );
   U8702 : OAI21_X1 port map( B1 => n5335, B2 => n5336, A => n7195, ZN => n5334
                           );
   U8703 : NAND4_X1 port map( A1 => n5345, A2 => n5346, A3 => n5347, A4 => 
                           n5348, ZN => n5335);
   U8704 : NAND4_X1 port map( A1 => n5337, A2 => n5338, A3 => n5339, A4 => 
                           n5340, ZN => n5336);
   U8705 : OAI21_X1 port map( B1 => n6960, B2 => n7191, A => n5315, ZN => n2604
                           );
   U8706 : OAI21_X1 port map( B1 => n5316, B2 => n5317, A => n7194, ZN => n5315
                           );
   U8707 : NAND4_X1 port map( A1 => n5326, A2 => n5327, A3 => n5328, A4 => 
                           n5329, ZN => n5316);
   U8708 : NAND4_X1 port map( A1 => n5318, A2 => n5319, A3 => n5320, A4 => 
                           n5321, ZN => n5317);
   U8709 : OAI21_X1 port map( B1 => n6961, B2 => n7191, A => n5296, ZN => n2606
                           );
   U8710 : OAI21_X1 port map( B1 => n5297, B2 => n5298, A => n7195, ZN => n5296
                           );
   U8711 : NAND4_X1 port map( A1 => n5307, A2 => n5308, A3 => n5309, A4 => 
                           n5310, ZN => n5297);
   U8712 : NAND4_X1 port map( A1 => n5299, A2 => n5300, A3 => n5301, A4 => 
                           n5302, ZN => n5298);
   U8713 : OAI21_X1 port map( B1 => n6962, B2 => n7191, A => n5277, ZN => n2608
                           );
   U8714 : OAI21_X1 port map( B1 => n5278, B2 => n5279, A => n7195, ZN => n5277
                           );
   U8715 : NAND4_X1 port map( A1 => n5288, A2 => n5289, A3 => n5290, A4 => 
                           n5291, ZN => n5278);
   U8716 : NAND4_X1 port map( A1 => n5280, A2 => n5281, A3 => n5282, A4 => 
                           n5283, ZN => n5279);
   U8717 : OAI21_X1 port map( B1 => n6963, B2 => n7191, A => n5258, ZN => n2610
                           );
   U8718 : OAI21_X1 port map( B1 => n5259, B2 => n5260, A => n7195, ZN => n5258
                           );
   U8719 : NAND4_X1 port map( A1 => n5269, A2 => n5270, A3 => n5271, A4 => 
                           n5272, ZN => n5259);
   U8720 : NAND4_X1 port map( A1 => n5261, A2 => n5262, A3 => n5263, A4 => 
                           n5264, ZN => n5260);
   U8721 : OAI21_X1 port map( B1 => n6964, B2 => n7191, A => n5239, ZN => n2612
                           );
   U8722 : OAI21_X1 port map( B1 => n5240, B2 => n5241, A => n7195, ZN => n5239
                           );
   U8723 : NAND4_X1 port map( A1 => n5250, A2 => n5251, A3 => n5252, A4 => 
                           n5253, ZN => n5240);
   U8724 : NAND4_X1 port map( A1 => n5242, A2 => n5243, A3 => n5244, A4 => 
                           n5245, ZN => n5241);
   U8725 : OAI21_X1 port map( B1 => n6965, B2 => n7191, A => n5220, ZN => n2614
                           );
   U8726 : OAI21_X1 port map( B1 => n5221, B2 => n5222, A => n7195, ZN => n5220
                           );
   U8727 : NAND4_X1 port map( A1 => n5231, A2 => n5232, A3 => n5233, A4 => 
                           n5234, ZN => n5221);
   U8728 : NAND4_X1 port map( A1 => n5223, A2 => n5224, A3 => n5225, A4 => 
                           n5226, ZN => n5222);
   U8729 : OAI21_X1 port map( B1 => n6966, B2 => n7191, A => n5201, ZN => n2616
                           );
   U8730 : OAI21_X1 port map( B1 => n5202, B2 => n5203, A => n7195, ZN => n5201
                           );
   U8731 : NAND4_X1 port map( A1 => n5212, A2 => n5213, A3 => n5214, A4 => 
                           n5215, ZN => n5202);
   U8732 : NAND4_X1 port map( A1 => n5204, A2 => n5205, A3 => n5206, A4 => 
                           n5207, ZN => n5203);
   U8733 : OAI21_X1 port map( B1 => n6967, B2 => n7191, A => n5182, ZN => n2618
                           );
   U8734 : OAI21_X1 port map( B1 => n5183, B2 => n5184, A => n7195, ZN => n5182
                           );
   U8735 : NAND4_X1 port map( A1 => n5193, A2 => n5194, A3 => n5195, A4 => 
                           n5196, ZN => n5183);
   U8736 : NAND4_X1 port map( A1 => n5185, A2 => n5186, A3 => n5187, A4 => 
                           n5188, ZN => n5184);
   U8737 : OAI21_X1 port map( B1 => n6968, B2 => n7191, A => n5163, ZN => n2620
                           );
   U8738 : OAI21_X1 port map( B1 => n5164, B2 => n5165, A => n7196, ZN => n5163
                           );
   U8739 : NAND4_X1 port map( A1 => n5174, A2 => n5175, A3 => n5176, A4 => 
                           n5177, ZN => n5164);
   U8740 : NAND4_X1 port map( A1 => n5166, A2 => n5167, A3 => n5168, A4 => 
                           n5169, ZN => n5165);
   U8741 : OAI22_X1 port map( A1 => n7235, A2 => n7479, B1 => n7234, B2 => 
                           n4905, ZN => n2720);
   U8742 : OAI22_X1 port map( A1 => n7235, A2 => n7482, B1 => n7234, B2 => 
                           n4904, ZN => n2721);
   U8743 : OAI22_X1 port map( A1 => n7235, A2 => n7485, B1 => n7234, B2 => 
                           n4903, ZN => n2722);
   U8744 : OAI22_X1 port map( A1 => n7235, A2 => n7488, B1 => n7234, B2 => 
                           n4902, ZN => n2723);
   U8745 : OAI22_X1 port map( A1 => n7235, A2 => n7491, B1 => n7234, B2 => 
                           n4901, ZN => n2724);
   U8746 : OAI22_X1 port map( A1 => n7236, A2 => n7494, B1 => n7234, B2 => 
                           n4900, ZN => n2725);
   U8747 : OAI22_X1 port map( A1 => n7236, A2 => n7497, B1 => n7234, B2 => 
                           n4899, ZN => n2726);
   U8748 : OAI22_X1 port map( A1 => n7236, A2 => n7500, B1 => n7234, B2 => 
                           n4898, ZN => n2727);
   U8749 : OAI22_X1 port map( A1 => n7236, A2 => n7503, B1 => n7234, B2 => 
                           n4897, ZN => n2728);
   U8750 : OAI22_X1 port map( A1 => n7236, A2 => n7506, B1 => n7234, B2 => 
                           n4896, ZN => n2729);
   U8751 : OAI22_X1 port map( A1 => n7237, A2 => n7509, B1 => n7234, B2 => 
                           n4895, ZN => n2730);
   U8752 : OAI22_X1 port map( A1 => n7237, A2 => n7512, B1 => n7234, B2 => 
                           n4894, ZN => n2731);
   U8753 : OAI22_X1 port map( A1 => n7237, A2 => n7515, B1 => n5106, B2 => 
                           n4893, ZN => n2732);
   U8754 : OAI22_X1 port map( A1 => n7237, A2 => n7518, B1 => n5106, B2 => 
                           n4892, ZN => n2733);
   U8755 : OAI22_X1 port map( A1 => n7237, A2 => n7521, B1 => n5106, B2 => 
                           n4891, ZN => n2734);
   U8756 : OAI22_X1 port map( A1 => n7238, A2 => n7524, B1 => n7234, B2 => 
                           n4890, ZN => n2735);
   U8757 : OAI22_X1 port map( A1 => n7238, A2 => n7527, B1 => n7234, B2 => 
                           n4889, ZN => n2736);
   U8758 : OAI22_X1 port map( A1 => n7238, A2 => n7530, B1 => n7234, B2 => 
                           n4888, ZN => n2737);
   U8759 : OAI22_X1 port map( A1 => n7238, A2 => n7533, B1 => n7234, B2 => 
                           n4887, ZN => n2738);
   U8760 : OAI22_X1 port map( A1 => n7238, A2 => n7536, B1 => n7234, B2 => 
                           n4886, ZN => n2739);
   U8761 : OAI22_X1 port map( A1 => n7239, A2 => n7539, B1 => n7234, B2 => 
                           n4885, ZN => n2740);
   U8762 : OAI22_X1 port map( A1 => n7239, A2 => n7542, B1 => n7234, B2 => 
                           n4884, ZN => n2741);
   U8763 : OAI22_X1 port map( A1 => n7239, A2 => n7545, B1 => n7234, B2 => 
                           n4883, ZN => n2742);
   U8764 : OAI22_X1 port map( A1 => n7239, A2 => n7548, B1 => n7234, B2 => 
                           n4882, ZN => n2743);
   U8765 : OAI22_X1 port map( A1 => n7239, A2 => n7551, B1 => n5106, B2 => 
                           n4881, ZN => n2744);
   U8766 : OAI22_X1 port map( A1 => n7240, A2 => n7554, B1 => n5106, B2 => 
                           n4880, ZN => n2745);
   U8767 : OAI22_X1 port map( A1 => n7240, A2 => n7557, B1 => n5106, B2 => 
                           n4879, ZN => n2746);
   U8768 : OAI22_X1 port map( A1 => n7240, A2 => n7560, B1 => n5106, B2 => 
                           n4878, ZN => n2747);
   U8769 : OAI22_X1 port map( A1 => n7240, A2 => n7563, B1 => n5106, B2 => 
                           n4877, ZN => n2748);
   U8770 : OAI22_X1 port map( A1 => n7240, A2 => n7566, B1 => n5106, B2 => 
                           n4876, ZN => n2749);
   U8771 : OAI22_X1 port map( A1 => n7241, A2 => n7569, B1 => n5106, B2 => 
                           n4875, ZN => n2750);
   U8772 : OAI22_X1 port map( A1 => n7241, A2 => n7581, B1 => n5106, B2 => 
                           n4874, ZN => n2751);
   U8773 : OAI22_X1 port map( A1 => n7307, A2 => n7478, B1 => n7306, B2 => 
                           n4713, ZN => n2976);
   U8774 : OAI22_X1 port map( A1 => n7307, A2 => n7481, B1 => n7306, B2 => 
                           n4712, ZN => n2977);
   U8775 : OAI22_X1 port map( A1 => n7307, A2 => n7484, B1 => n7306, B2 => 
                           n4711, ZN => n2978);
   U8776 : OAI22_X1 port map( A1 => n7307, A2 => n7487, B1 => n7306, B2 => 
                           n4710, ZN => n2979);
   U8777 : OAI22_X1 port map( A1 => n7307, A2 => n7490, B1 => n7306, B2 => 
                           n4709, ZN => n2980);
   U8778 : OAI22_X1 port map( A1 => n7308, A2 => n7493, B1 => n7306, B2 => 
                           n4708, ZN => n2981);
   U8779 : OAI22_X1 port map( A1 => n7308, A2 => n7496, B1 => n7306, B2 => 
                           n4707, ZN => n2982);
   U8780 : OAI22_X1 port map( A1 => n7308, A2 => n7499, B1 => n7306, B2 => 
                           n4706, ZN => n2983);
   U8781 : OAI22_X1 port map( A1 => n7308, A2 => n7502, B1 => n7306, B2 => 
                           n4705, ZN => n2984);
   U8782 : OAI22_X1 port map( A1 => n7308, A2 => n7505, B1 => n7306, B2 => 
                           n4704, ZN => n2985);
   U8783 : OAI22_X1 port map( A1 => n7309, A2 => n7508, B1 => n7306, B2 => 
                           n4703, ZN => n2986);
   U8784 : OAI22_X1 port map( A1 => n7309, A2 => n7511, B1 => n7306, B2 => 
                           n4702, ZN => n2987);
   U8785 : OAI22_X1 port map( A1 => n7309, A2 => n7514, B1 => n5097, B2 => 
                           n4701, ZN => n2988);
   U8786 : OAI22_X1 port map( A1 => n7309, A2 => n7517, B1 => n5097, B2 => 
                           n4700, ZN => n2989);
   U8787 : OAI22_X1 port map( A1 => n7309, A2 => n7520, B1 => n5097, B2 => 
                           n4699, ZN => n2990);
   U8788 : OAI22_X1 port map( A1 => n7310, A2 => n7523, B1 => n7306, B2 => 
                           n4698, ZN => n2991);
   U8789 : OAI22_X1 port map( A1 => n7310, A2 => n7526, B1 => n7306, B2 => 
                           n4697, ZN => n2992);
   U8790 : OAI22_X1 port map( A1 => n7310, A2 => n7529, B1 => n7306, B2 => 
                           n4696, ZN => n2993);
   U8791 : OAI22_X1 port map( A1 => n7310, A2 => n7532, B1 => n7306, B2 => 
                           n4695, ZN => n2994);
   U8792 : OAI22_X1 port map( A1 => n7310, A2 => n7535, B1 => n7306, B2 => 
                           n4694, ZN => n2995);
   U8793 : OAI22_X1 port map( A1 => n7311, A2 => n7538, B1 => n7306, B2 => 
                           n4693, ZN => n2996);
   U8794 : OAI22_X1 port map( A1 => n7311, A2 => n7541, B1 => n7306, B2 => 
                           n4692, ZN => n2997);
   U8795 : OAI22_X1 port map( A1 => n7311, A2 => n7544, B1 => n7306, B2 => 
                           n4691, ZN => n2998);
   U8796 : OAI22_X1 port map( A1 => n7311, A2 => n7547, B1 => n7306, B2 => 
                           n4690, ZN => n2999);
   U8797 : OAI22_X1 port map( A1 => n7311, A2 => n7550, B1 => n5097, B2 => 
                           n4689, ZN => n3000);
   U8798 : OAI22_X1 port map( A1 => n7312, A2 => n7553, B1 => n5097, B2 => 
                           n4688, ZN => n3001);
   U8799 : OAI22_X1 port map( A1 => n7312, A2 => n7556, B1 => n5097, B2 => 
                           n4687, ZN => n3002);
   U8800 : OAI22_X1 port map( A1 => n7312, A2 => n7559, B1 => n5097, B2 => 
                           n4686, ZN => n3003);
   U8801 : OAI22_X1 port map( A1 => n7312, A2 => n7562, B1 => n5097, B2 => 
                           n4685, ZN => n3004);
   U8802 : OAI22_X1 port map( A1 => n7312, A2 => n7565, B1 => n5097, B2 => 
                           n4684, ZN => n3005);
   U8803 : OAI22_X1 port map( A1 => n7313, A2 => n7568, B1 => n5097, B2 => 
                           n4683, ZN => n3006);
   U8804 : OAI22_X1 port map( A1 => n7313, A2 => n7580, B1 => n5097, B2 => 
                           n4682, ZN => n3007);
   U8805 : OAI22_X1 port map( A1 => n7379, A2 => n7477, B1 => n7378, B2 => 
                           n4521, ZN => n3232);
   U8806 : OAI22_X1 port map( A1 => n7379, A2 => n7480, B1 => n7378, B2 => 
                           n4520, ZN => n3233);
   U8807 : OAI22_X1 port map( A1 => n7379, A2 => n7483, B1 => n7378, B2 => 
                           n4519, ZN => n3234);
   U8808 : OAI22_X1 port map( A1 => n7379, A2 => n7486, B1 => n7378, B2 => 
                           n4518, ZN => n3235);
   U8809 : OAI22_X1 port map( A1 => n7379, A2 => n7489, B1 => n7378, B2 => 
                           n4517, ZN => n3236);
   U8810 : OAI22_X1 port map( A1 => n7380, A2 => n7492, B1 => n7378, B2 => 
                           n4516, ZN => n3237);
   U8811 : OAI22_X1 port map( A1 => n7380, A2 => n7495, B1 => n7378, B2 => 
                           n4515, ZN => n3238);
   U8812 : OAI22_X1 port map( A1 => n7380, A2 => n7498, B1 => n7378, B2 => 
                           n4514, ZN => n3239);
   U8813 : OAI22_X1 port map( A1 => n7380, A2 => n7501, B1 => n7378, B2 => 
                           n4513, ZN => n3240);
   U8814 : OAI22_X1 port map( A1 => n7380, A2 => n7504, B1 => n7378, B2 => 
                           n4512, ZN => n3241);
   U8815 : OAI22_X1 port map( A1 => n7381, A2 => n7507, B1 => n7378, B2 => 
                           n4511, ZN => n3242);
   U8816 : OAI22_X1 port map( A1 => n7381, A2 => n7510, B1 => n7378, B2 => 
                           n4510, ZN => n3243);
   U8817 : OAI22_X1 port map( A1 => n7381, A2 => n7513, B1 => n5088, B2 => 
                           n4509, ZN => n3244);
   U8818 : OAI22_X1 port map( A1 => n7381, A2 => n7516, B1 => n5088, B2 => 
                           n4508, ZN => n3245);
   U8819 : OAI22_X1 port map( A1 => n7381, A2 => n7519, B1 => n5088, B2 => 
                           n4507, ZN => n3246);
   U8820 : OAI22_X1 port map( A1 => n7382, A2 => n7522, B1 => n7378, B2 => 
                           n4506, ZN => n3247);
   U8821 : OAI22_X1 port map( A1 => n7382, A2 => n7525, B1 => n7378, B2 => 
                           n4505, ZN => n3248);
   U8822 : OAI22_X1 port map( A1 => n7382, A2 => n7528, B1 => n7378, B2 => 
                           n4504, ZN => n3249);
   U8823 : OAI22_X1 port map( A1 => n7382, A2 => n7531, B1 => n7378, B2 => 
                           n4503, ZN => n3250);
   U8824 : OAI22_X1 port map( A1 => n7382, A2 => n7534, B1 => n7378, B2 => 
                           n4502, ZN => n3251);
   U8825 : OAI22_X1 port map( A1 => n7383, A2 => n7537, B1 => n7378, B2 => 
                           n4501, ZN => n3252);
   U8826 : OAI22_X1 port map( A1 => n7383, A2 => n7540, B1 => n7378, B2 => 
                           n4500, ZN => n3253);
   U8827 : OAI22_X1 port map( A1 => n7383, A2 => n7543, B1 => n7378, B2 => 
                           n4499, ZN => n3254);
   U8828 : OAI22_X1 port map( A1 => n7383, A2 => n7546, B1 => n7378, B2 => 
                           n4498, ZN => n3255);
   U8829 : OAI22_X1 port map( A1 => n7383, A2 => n7549, B1 => n5088, B2 => 
                           n4497, ZN => n3256);
   U8830 : OAI22_X1 port map( A1 => n7384, A2 => n7552, B1 => n5088, B2 => 
                           n4496, ZN => n3257);
   U8831 : OAI22_X1 port map( A1 => n7384, A2 => n7555, B1 => n5088, B2 => 
                           n4495, ZN => n3258);
   U8832 : OAI22_X1 port map( A1 => n7384, A2 => n7558, B1 => n5088, B2 => 
                           n4494, ZN => n3259);
   U8833 : OAI22_X1 port map( A1 => n7384, A2 => n7561, B1 => n5088, B2 => 
                           n4493, ZN => n3260);
   U8834 : OAI22_X1 port map( A1 => n7384, A2 => n7564, B1 => n5088, B2 => 
                           n4492, ZN => n3261);
   U8835 : OAI22_X1 port map( A1 => n7385, A2 => n7567, B1 => n5088, B2 => 
                           n4491, ZN => n3262);
   U8836 : OAI22_X1 port map( A1 => n7385, A2 => n7579, B1 => n5088, B2 => 
                           n4490, ZN => n3263);
   U8837 : OAI22_X1 port map( A1 => n7451, A2 => n7477, B1 => n7450, B2 => 
                           n4329, ZN => n3488);
   U8838 : OAI22_X1 port map( A1 => n7451, A2 => n7480, B1 => n7450, B2 => 
                           n4328, ZN => n3489);
   U8839 : OAI22_X1 port map( A1 => n7451, A2 => n7483, B1 => n7450, B2 => 
                           n4327, ZN => n3490);
   U8840 : OAI22_X1 port map( A1 => n7451, A2 => n7486, B1 => n7450, B2 => 
                           n4326, ZN => n3491);
   U8841 : OAI22_X1 port map( A1 => n7451, A2 => n7489, B1 => n7450, B2 => 
                           n4325, ZN => n3492);
   U8842 : OAI22_X1 port map( A1 => n7452, A2 => n7492, B1 => n7450, B2 => 
                           n4324, ZN => n3493);
   U8843 : OAI22_X1 port map( A1 => n7452, A2 => n7495, B1 => n7450, B2 => 
                           n4323, ZN => n3494);
   U8844 : OAI22_X1 port map( A1 => n7452, A2 => n7498, B1 => n7450, B2 => 
                           n4322, ZN => n3495);
   U8845 : OAI22_X1 port map( A1 => n7452, A2 => n7501, B1 => n7450, B2 => 
                           n4321, ZN => n3496);
   U8846 : OAI22_X1 port map( A1 => n7452, A2 => n7504, B1 => n7450, B2 => 
                           n4320, ZN => n3497);
   U8847 : OAI22_X1 port map( A1 => n7453, A2 => n7507, B1 => n7450, B2 => 
                           n4319, ZN => n3498);
   U8848 : OAI22_X1 port map( A1 => n7453, A2 => n7510, B1 => n7450, B2 => 
                           n4318, ZN => n3499);
   U8849 : OAI22_X1 port map( A1 => n7453, A2 => n7513, B1 => n5073, B2 => 
                           n4317, ZN => n3500);
   U8850 : OAI22_X1 port map( A1 => n7453, A2 => n7516, B1 => n5073, B2 => 
                           n4316, ZN => n3501);
   U8851 : OAI22_X1 port map( A1 => n7453, A2 => n7519, B1 => n5073, B2 => 
                           n4315, ZN => n3502);
   U8852 : OAI22_X1 port map( A1 => n7454, A2 => n7522, B1 => n7450, B2 => 
                           n4314, ZN => n3503);
   U8853 : OAI22_X1 port map( A1 => n7454, A2 => n7525, B1 => n7450, B2 => 
                           n4313, ZN => n3504);
   U8854 : OAI22_X1 port map( A1 => n7454, A2 => n7528, B1 => n7450, B2 => 
                           n4312, ZN => n3505);
   U8855 : OAI22_X1 port map( A1 => n7454, A2 => n7531, B1 => n7450, B2 => 
                           n4311, ZN => n3506);
   U8856 : OAI22_X1 port map( A1 => n7454, A2 => n7534, B1 => n7450, B2 => 
                           n4310, ZN => n3507);
   U8857 : OAI22_X1 port map( A1 => n7455, A2 => n7537, B1 => n7450, B2 => 
                           n4309, ZN => n3508);
   U8858 : OAI22_X1 port map( A1 => n7455, A2 => n7540, B1 => n7450, B2 => 
                           n4308, ZN => n3509);
   U8859 : OAI22_X1 port map( A1 => n7455, A2 => n7543, B1 => n7450, B2 => 
                           n4307, ZN => n3510);
   U8860 : OAI22_X1 port map( A1 => n7455, A2 => n7546, B1 => n7450, B2 => 
                           n4306, ZN => n3511);
   U8861 : OAI22_X1 port map( A1 => n7455, A2 => n7549, B1 => n5073, B2 => 
                           n4305, ZN => n3512);
   U8862 : OAI22_X1 port map( A1 => n7456, A2 => n7552, B1 => n5073, B2 => 
                           n4304, ZN => n3513);
   U8863 : OAI22_X1 port map( A1 => n7456, A2 => n7555, B1 => n5073, B2 => 
                           n4303, ZN => n3514);
   U8864 : OAI22_X1 port map( A1 => n7456, A2 => n7558, B1 => n5073, B2 => 
                           n4302, ZN => n3515);
   U8865 : OAI22_X1 port map( A1 => n7456, A2 => n7561, B1 => n5073, B2 => 
                           n4301, ZN => n3516);
   U8866 : OAI22_X1 port map( A1 => n7456, A2 => n7564, B1 => n5073, B2 => 
                           n4300, ZN => n3517);
   U8867 : OAI22_X1 port map( A1 => n7457, A2 => n7567, B1 => n5073, B2 => 
                           n4299, ZN => n3518);
   U8868 : OAI22_X1 port map( A1 => n7457, A2 => n7579, B1 => n5073, B2 => 
                           n4298, ZN => n3519);
   U8869 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n6400);
   U8870 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n5747);
   U8871 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n4262, 
                           ZN => n6401);
   U8872 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n4265, 
                           ZN => n5748);
   U8873 : NOR2_X1 port map( A1 => n4260, A2 => ADD_RD1(4), ZN => n6412);
   U8874 : NOR2_X1 port map( A1 => n4263, A2 => ADD_RD2(4), ZN => n5759);
   U8875 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n6415);
   U8876 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n5762);
   U8877 : NOR3_X1 port map( A1 => n4262, A2 => ADD_RD1(2), A3 => n4261, ZN => 
                           n6403);
   U8878 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n4261, 
                           ZN => n6402);
   U8879 : NOR3_X1 port map( A1 => n4265, A2 => ADD_RD2(2), A3 => n4264, ZN => 
                           n5750);
   U8880 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n4264, 
                           ZN => n5749);
   U8881 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n6394);
   U8882 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n4260, ZN => n6405);
   U8883 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n5741);
   U8884 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n4263, ZN => n5752);
   U8885 : INV_X1 port map( A => RESET, ZN => n4254);
   U8886 : AND3_X1 port map( A1 => n4262, A2 => n4261, A3 => ADD_RD1(2), ZN => 
                           n6396);
   U8887 : AND3_X1 port map( A1 => n4265, A2 => n4264, A3 => ADD_RD2(2), ZN => 
                           n5743);
   U8888 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n4261, A3 => ADD_RD1(2), 
                           ZN => n6395);
   U8889 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n4264, A3 => ADD_RD2(2), 
                           ZN => n5742);
   U8890 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n5764);
   U8891 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n5111);
   U8892 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n7583, ZN => n5058);
   U8893 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n7583, ZN => n5057);
   U8894 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n7583, ZN => n5056);
   U8895 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n7583, ZN => n5055);
   U8896 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n7583, ZN => n5054);
   U8897 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n7583, ZN => n5053);
   U8898 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n7583, ZN => n5052);
   U8899 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n7583, ZN => n5051);
   U8900 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n7583, ZN => n5050);
   U8901 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n7583, ZN => n5049);
   U8902 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n7583, ZN => n5048);
   U8903 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n7583, ZN => n5047);
   U8904 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n7582, ZN => n5046);
   U8905 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n7582, ZN => n5045);
   U8906 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n7582, ZN => n5044);
   U8907 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n7582, ZN => n5043);
   U8908 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n7582, ZN => n5042);
   U8909 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n7582, ZN => n5041);
   U8910 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n7582, ZN => n5040);
   U8911 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n7582, ZN => n5039);
   U8912 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n7582, ZN => n5038);
   U8913 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n7582, ZN => n5037);
   U8914 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n7582, ZN => n5036);
   U8915 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n7582, ZN => n5034);
   U8916 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n7584, ZN => n5066);
   U8917 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n7584, ZN => n5065);
   U8918 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n7584, ZN => n5064);
   U8919 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n7584, ZN => n5063);
   U8920 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n7584, ZN => n5062);
   U8921 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n7584, ZN => n5061);
   U8922 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n7584, ZN => n5060);
   U8923 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n7584, ZN => n5059);
   U8924 : INV_X1 port map( A => ADD_RD1(1), ZN => n4261);
   U8925 : INV_X1 port map( A => ADD_RD2(1), ZN => n4264);
   U8926 : INV_X1 port map( A => ADD_RD1(0), ZN => n4262);
   U8927 : INV_X1 port map( A => ADD_RD2(0), ZN => n4265);
   U8928 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n4262, A3 => ADD_RD1(1), 
                           ZN => n6398);
   U8929 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n4265, A3 => ADD_RD2(1), 
                           ZN => n5745);
   U8930 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(1), ZN => n6397);
   U8931 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(1), ZN => n5744);
   U8932 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n5083);
   U8933 : INV_X1 port map( A => ADD_WR(2), ZN => n4257);
   U8934 : INV_X1 port map( A => ADD_WR(0), ZN => n4259);
   U8935 : INV_X1 port map( A => ADD_WR(1), ZN => n4258);
   U8936 : INV_X1 port map( A => ADD_RD1(3), ZN => n4260);
   U8937 : INV_X1 port map( A => ADD_RD2(3), ZN => n4263);
   U8938 : INV_X1 port map( A => ADD_WR(4), ZN => n4255);
   U8939 : INV_X1 port map( A => ADD_WR(3), ZN => n4256);
   U8940 : CLKBUF_X1 port map( A => n5764, Z => n7094);
   U8941 : CLKBUF_X1 port map( A => n5111, Z => n7196);
   U8942 : CLKBUF_X1 port map( A => n4254, Z => n7587);

end SYN_A;
