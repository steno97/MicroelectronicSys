
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windRF_M8_N8_F2_NBIT64 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windRF_M8_N8_F2_NBIT64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windRF_M8_N8_F2_NBIT64.all;

entity windRF_M8_N8_F2_NBIT64 is

   port( CLK, RESET, ENABLE, CALL, RETRN : in std_logic;  FILL, SPILL : out 
         std_logic;  BUSin : in std_logic_vector (63 downto 0);  BUSout : out 
         std_logic_vector (63 downto 0);  RD1, RD2, WR : in std_logic;  ADD_WR,
         ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end windRF_M8_N8_F2_NBIT64;

architecture SYN_bhv of windRF_M8_N8_F2_NBIT64 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal i_3_port, i_2_port, i_1_port, N659, N660, N661, N688, N689, N690, 
      N811, N812, N813, N929, N930, N931, N932, N6270, N6271, N6272, N6273, 
      N6395, N6396, N6397, N6398, U3_U193_Z_1, U3_U193_Z_2, U3_U193_Z_3, 
      U3_U193_Z_4, U3_U194_Z_1, U3_U194_Z_2, U3_U194_Z_3, U3_U194_Z_4, 
      U3_U195_Z_1, U3_U195_Z_2, U3_U195_Z_3, U3_U195_Z_4, n59, n60, n61, n62, 
      n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77
      , n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
      n92, n93, n94, n95, n96, n97, n98, n99, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811_port, n812_port, n813_port
      , n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
      n826, n2683, n2695, n2696, n2697, n2698, n2699, n2700, n2706, n2707, 
      n2709, n2710, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
      n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
      n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
      n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, 
      n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, 
      n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, 
      n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, 
      n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, 
      n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, 
      n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
      n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, 
      n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, 
      n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, 
      n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, 
      n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, 
      n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, 
      n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, 
      n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, 
      n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, 
      n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, 
      n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, 
      n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, 
      n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, 
      n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, 
      n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, 
      n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, 
      n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, 
      n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, 
      n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, 
      n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, 
      n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, 
      n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, 
      n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, 
      n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, 
      n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, 
      n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, 
      n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, 
      n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, 
      n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, 
      n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, 
      n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, 
      n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, 
      n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, 
      n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, 
      n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, 
      n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, 
      n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, 
      n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, 
      n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, 
      n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, 
      n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, 
      n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, 
      n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, 
      n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, 
      n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, 
      n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, 
      n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, 
      n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, 
      n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, 
      n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, 
      n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, 
      n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, 
      n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, 
      n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, 
      n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, 
      n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, 
      n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, 
      n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, 
      n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, 
      n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, 
      n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, 
      n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
      n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, 
      n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, 
      n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, 
      n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, 
      n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, 
      n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, 
      n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, 
      n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, 
      n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, 
      n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, 
      n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, 
      n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
      n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, 
      n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, 
      n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, 
      n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
      n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, 
      n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, 
      n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, 
      n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, 
      n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, 
      n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, 
      n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, 
      n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, 
      n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, 
      n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, 
      n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, 
      n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, 
      n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, 
      n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, 
      n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, 
      n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, 
      n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, 
      n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, 
      n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, 
      n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, 
      n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, 
      n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, 
      n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, 
      n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, 
      n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, 
      n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, 
      n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, 
      n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, 
      n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, 
      n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, 
      n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, 
      n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, 
      n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, 
      n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, 
      n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, 
      n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
      n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, 
      n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, 
      n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, 
      n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, 
      n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, 
      n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
      n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, 
      n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, 
      n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, 
      n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, 
      n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, 
      n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, 
      n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, 
      n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
      n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, 
      n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, 
      n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, 
      n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, 
      n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, 
      n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, 
      n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, 
      n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, 
      n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, 
      n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, 
      n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, 
      n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, 
      n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, 
      n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, 
      n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, 
      n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, 
      n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, 
      n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, 
      n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, 
      n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
      n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, 
      n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
      n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
      n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, 
      n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
      n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, 
      n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, 
      n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, 
      n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, 
      n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, 
      n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, 
      n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, 
      n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, 
      n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, 
      n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, 
      n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, 
      n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, 
      n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, 
      n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, 
      n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, 
      n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, 
      n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, 
      n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, 
      n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, 
      n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
      n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, 
      n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, 
      n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
      n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
      n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
      n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, 
      n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, 
      n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, 
      n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
      n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, 
      n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, 
      n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, 
      n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, 
      n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, 
      n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, 
      n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, 
      n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, 
      n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
      n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, 
      n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, 
      n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, 
      n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
      n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, 
      n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, 
      n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, 
      n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, 
      n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, 
      n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, 
      n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, 
      n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, 
      n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, 
      n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, 
      n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, 
      n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, 
      n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, 
      n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, 
      n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, 
      n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, 
      n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
      n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, 
      n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, 
      n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, 
      n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
      n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, 
      n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, 
      n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, 
      n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
      n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, 
      n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, 
      n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, 
      n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
      n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, 
      n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, 
      n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, 
      n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9895, n9896, 
      n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, 
      n9907, add_146_carry_2_port, add_146_carry_3_port, add_146_carry_4_port, 
      n12791, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, 
      n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, 
      n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, 
      n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, 
      n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, 
      n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, 
      n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, 
      n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, 
      n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, 
      n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, 
      n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, 
      n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, 
      n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, 
      n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, 
      n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, 
      n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, 
      n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, 
      n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, 
      n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, 
      n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, 
      n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, 
      n17066, n17067, n17068, n17069, n23853, n25394, r510_n3, 
      r510_carry_2_port, r510_carry_3_port, r510_carry_4_port, 
      r510_carry_5_port, r504_n3, r504_carry_2_port, r504_carry_3_port, 
      r504_carry_4_port, r504_carry_5_port, r498_n1, r498_carry_2_port, 
      r498_carry_3_port, r498_carry_4_port, r498_carry_5_port, 
      add_136_carry_2_port, add_136_carry_3_port, add_136_carry_4_port, n25395,
      n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, 
      n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, 
      n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, 
      n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, 
      n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, 
      n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, 
      n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, 
      n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, 
      n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, 
      n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, 
      n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, 
      n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, 
      n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n27870, 
      n27871, n27872, n27874, n27921, n27922, n27923, n27924, n27925, n27926, 
      n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, 
      n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, 
      n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, 
      n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, 
      n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, 
      n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, 
      n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, 
      n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, 
      n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, 
      n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, 
      n28849, n28850, n29043, n29044, n29045, n29046, n29047, n29048, n29049, 
      n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, 
      n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, 
      n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, 
      n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, 
      n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, 
      n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, 
      n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, 
      n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, 
      n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, 
      n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, 
      n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, 
      n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, 
      n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, 
      n29167, n29168, n29169, n29170, n29363, n29364, n29365, n29366, n29367, 
      n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, 
      n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, 
      n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, 
      n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, 
      n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, 
      n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, 
      n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, 
      n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, 
      n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, 
      n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, 
      n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, 
      n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, 
      n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, 
      n29485, n29486, n29487, n29488, n29489, n29490, n29683, n29684, n29685, 
      n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, 
      n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, 
      n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, 
      n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, 
      n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, 
      n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, 
      n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, 
      n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, 
      n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, 
      n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, 
      n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, 
      n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, 
      n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, 
      n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n30003, 
      n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, 
      n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, 
      n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, 
      n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, 
      n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, 
      n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, 
      n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, 
      n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, 
      n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, 
      n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, 
      n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, 
      n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, 
      n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, 
      n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, 
      n30130, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, 
      n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, 
      n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, 
      n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, 
      n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, 
      n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, 
      n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, 
      n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, 
      n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, 
      n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, 
      n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, 
      n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, 
      n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, 
      n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, 
      n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, 
      n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, 
      n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, 
      n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, 
      n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, 
      n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, 
      n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, 
      n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, 
      n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, 
      n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, 
      n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, 
      n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, 
      n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, 
      n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, 
      n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, 
      n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, 
      n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, 
      n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, 
      n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, 
      n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, 
      n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, 
      n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, 
      n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, 
      n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, 
      n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, 
      n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, 
      n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, 
      n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, 
      n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, 
      n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, 
      n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, 
      n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, 
      n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, 
      n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, 
      n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, 
      n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, 
      n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, 
      n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, 
      n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, 
      n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, 
      n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, 
      n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, 
      n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, 
      n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, 
      n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, 
      n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, 
      n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, 
      n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, 
      n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, 
      n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, 
      n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, 
      n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, 
      n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, 
      n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, 
      n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, 
      n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, 
      n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, 
      n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, 
      n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, 
      n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, 
      n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, 
      n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, 
      n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, 
      n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, 
      n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, 
      n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, 
      n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, 
      n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, 
      n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, 
      n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, 
      n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, 
      n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, 
      n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, 
      n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, 
      n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, 
      n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, 
      n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, 
      n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, 
      n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, 
      n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, 
      n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, 
      n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, 
      n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, 
      n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, 
      n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, 
      n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, 
      n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, 
      n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, 
      n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, 
      n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, 
      n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, 
      n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, 
      n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, 
      n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, 
      n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, 
      n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, 
      n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, 
      n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, 
      n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, 
      n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, 
      n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, 
      n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, 
      n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, 
      n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, 
      n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, 
      n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, 
      n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, 
      n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, 
      n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, 
      n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, 
      n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, 
      n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, 
      n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, 
      n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, 
      n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, 
      n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, 
      n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, 
      n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, 
      n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, 
      n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, 
      n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, 
      n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, 
      n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, 
      n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, 
      n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, 
      n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, 
      n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, 
      n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, 
      n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, 
      n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, 
      n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, 
      n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, 
      n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, 
      n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, 
      n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, 
      n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, 
      n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, 
      n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, 
      n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, 
      n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, 
      n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, 
      n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, 
      n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, 
      n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, 
      n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, 
      n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, 
      n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, 
      n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, 
      n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, 
      n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, 
      n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, 
      n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, 
      n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, 
      n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, 
      n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, 
      n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, 
      n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, 
      n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, 
      n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, 
      n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, 
      n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, 
      n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, 
      n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, 
      n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, 
      n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, 
      n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, 
      n32077, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, 
      n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, 
      n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, 
      n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, 
      n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, 
      n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, 
      n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, 
      n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, 
      n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, 
      n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, 
      n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, 
      n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, 
      n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, 
      n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, 
      n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, 
      n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, 
      n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, 
      n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, 
      n32240, n32241, n32242, n32243, n32244, n32246, n32247, n32248, n32249, 
      n32251, n32253, n32254, n32255, n32258, n32259, n32260, n32261, n32262, 
      n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, 
      n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, 
      n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, 
      n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, 
      n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, 
      n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, 
      n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32384, n32444, 
      n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, 
      n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, 
      n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, 
      n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, 
      n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, 
      n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, 
      n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, 
      n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, 
      n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, 
      n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, 
      n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, 
      n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, 
      n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, 
      n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, 
      n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, 
      n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, 
      n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, 
      n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, 
      n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, 
      n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, 
      n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, 
      n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, 
      n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, 
      n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, 
      n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, 
      n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, 
      n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, 
      n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, 
      n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, 
      n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, 
      n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, 
      n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, 
      n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, 
      n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, 
      n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, 
      n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, 
      n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, 
      n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, 
      n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, 
      n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, 
      n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, 
      n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, 
      n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, 
      n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, 
      n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, 
      n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, 
      n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, 
      n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, 
      n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, 
      n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, 
      n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, 
      n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, 
      n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, 
      n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, 
      n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, 
      n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, 
      n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, 
      n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, 
      n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, 
      n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, 
      n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, 
      n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, 
      n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, 
      n33037, n33038, n33087, n33088, n33089, n33090, n33091, n33092, n33093, 
      n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, 
      n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, 
      n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, 
      n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, 
      n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33139, 
      n33195, n33196, n33197, n33199, n33207, n33208, n33209, n33210, n33211, 
      n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, 
      n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, 
      n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, 
      n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, 
      n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, 
      n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, 
      n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, 
      n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, 
      n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, 
      n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, 
      n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, 
      n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, 
      n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, 
      n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, 
      n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, 
      n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, 
      n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, 
      n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, 
      n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, 
      n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, 
      n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, 
      n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, 
      n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, 
      n33419, n33420, n33422, n33423, n33424, n33425, n33426, n33427, n33428, 
      n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, 
      n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, 
      n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, 
      n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, 
      n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, 
      n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, 
      n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, 
      n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, 
      n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, 
      n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, 
      n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, 
      n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, 
      n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, 
      n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, 
      n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, 
      n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, 
      n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, 
      n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, 
      n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, 
      n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, 
      n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, 
      n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, 
      n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, 
      n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, 
      n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, 
      n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, 
      n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, 
      n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, 
      n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, 
      n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, 
      n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, 
      n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, 
      n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, 
      n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, 
      n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, 
      n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, 
      n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, 
      n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, 
      n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, 
      n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, 
      n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, 
      n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, 
      n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, 
      n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, 
      n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, 
      n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, 
      n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, 
      n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, 
      n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, 
      n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, 
      n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, 
      n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, 
      n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, 
      n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, 
      n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, 
      n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, 
      n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, 
      n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, 
      n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, 
      n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, 
      n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, 
      n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, 
      n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, 
      n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, 
      n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, 
      n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, 
      n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, 
      n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, 
      n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, 
      n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, 
      n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, 
      n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, 
      n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, 
      n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, 
      n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, 
      n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, 
      n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, 
      n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, 
      n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, 
      n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, 
      n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, 
      n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, 
      n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, 
      n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, 
      n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, 
      n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, 
      n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, 
      n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, 
      n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, 
      n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, 
      n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, 
      n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, 
      n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, 
      n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, 
      n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, 
      n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, 
      n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, 
      n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, 
      n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, 
      n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, 
      n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, 
      n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, 
      n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, 
      n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, 
      n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, 
      n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, 
      n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, 
      n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, 
      n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, 
      n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, 
      n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, 
      n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, 
      n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, 
      n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, 
      n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, 
      n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, 
      n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, 
      n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, 
      n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, 
      n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, 
      n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, 
      n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, 
      n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, 
      n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, 
      n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, 
      n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, 
      n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, 
      n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, 
      n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, 
      n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, 
      n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, 
      n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, 
      n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, 
      n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, 
      n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, 
      n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, 
      n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, 
      n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, 
      n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, 
      n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, 
      n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, 
      n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, 
      n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, 
      n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, 
      n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, 
      n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, 
      n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, 
      n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, 
      n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, 
      n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, 
      n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, 
      n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, 
      n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, 
      n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, 
      n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, 
      n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, 
      n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, 
      n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, 
      n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, 
      n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, 
      n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, 
      n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, 
      n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, 
      n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, 
      n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, 
      n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, 
      n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, 
      n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, 
      n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, 
      n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, 
      n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, 
      n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, 
      n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, 
      n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, 
      n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, 
      n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, 
      n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, 
      n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, 
      n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, 
      n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, 
      n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, 
      n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, 
      n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, 
      n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, 
      n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, 
      n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, 
      n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, 
      n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, 
      n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, 
      n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, 
      n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, 
      n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, 
      n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, 
      n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, 
      n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, 
      n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, 
      n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, 
      n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, 
      n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, 
      n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, 
      n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, 
      n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, 
      n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, 
      n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, 
      n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, 
      n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, 
      n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, 
      n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, 
      n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, 
      n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, 
      n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, 
      n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, 
      n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, 
      n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, 
      n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, 
      n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, 
      n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, 
      n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, 
      n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, 
      n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, 
      n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, 
      n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, 
      n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, 
      n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, 
      n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, 
      n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, 
      n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, 
      n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, 
      n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, 
      n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, 
      n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, 
      n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, 
      n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, 
      n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, 
      n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, 
      n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, 
      n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, 
      n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, 
      n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, 
      n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, 
      n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, 
      n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, 
      n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, 
      n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, 
      n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, 
      n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, 
      n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, 
      n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, 
      n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, 
      n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, 
      n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, 
      n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, 
      n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, 
      n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, 
      n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, 
      n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, 
      n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, 
      n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, 
      n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, 
      n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, 
      n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, 
      n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, 
      n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, 
      n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, 
      n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, 
      n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, 
      n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, 
      n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, 
      n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, 
      n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, 
      n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, 
      n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, 
      n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, 
      n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, 
      n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, 
      n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, 
      n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, 
      n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, 
      n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, 
      n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, 
      n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, 
      n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, 
      n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, 
      n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, 
      n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, 
      n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, 
      n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, 
      n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, 
      n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, 
      n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, 
      n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, 
      n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, 
      n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, 
      n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, 
      n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, 
      n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, 
      n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, 
      n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, 
      n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, 
      n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, 
      n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, 
      n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, 
      n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, 
      n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, 
      n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, 
      n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, 
      n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, 
      n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, 
      n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, 
      n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, 
      n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, 
      n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, 
      n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, 
      n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, 
      n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, 
      n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, 
      n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, 
      n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, 
      n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, 
      n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, 
      n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, 
      n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, 
      n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, 
      n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, 
      n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, 
      n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, 
      n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, 
      n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, 
      n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, 
      n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, 
      n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, 
      n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, 
      n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, 
      n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, 
      n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, 
      n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, 
      n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, 
      n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, 
      n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, 
      n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, 
      n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, 
      n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, 
      n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, 
      n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, 
      n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, 
      n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, 
      n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, 
      n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, 
      n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, 
      n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, 
      n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, 
      n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, 
      n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, 
      n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, 
      n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, 
      n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, 
      n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, 
      n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, 
      n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, 
      n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, 
      n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, 
      n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, 
      n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, 
      n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, 
      n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, 
      n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, 
      n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, 
      n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, 
      n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, 
      n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, 
      n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, 
      n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, 
      n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, 
      n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, 
      n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, 
      n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, 
      n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, 
      n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, 
      n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, 
      n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, 
      n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, 
      n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, 
      n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, 
      n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, 
      n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, 
      n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, 
      n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, 
      n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, 
      n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, 
      n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, 
      n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, 
      n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, 
      n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, 
      n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, 
      n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, 
      n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, 
      n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, 
      n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, 
      n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, 
      n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, 
      n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, 
      n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, 
      n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, 
      n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, 
      n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, 
      n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, 
      n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, 
      n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, 
      n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, 
      n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, 
      n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, 
      n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, 
      n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, 
      n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, 
      n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, 
      n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, 
      n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, 
      n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, 
      n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, 
      n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, 
      n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, 
      n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, 
      n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, 
      n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, 
      n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n38789, 
      n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, 
      n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, 
      n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, 
      n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, 
      n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, 
      n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, 
      n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, 
      n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, 
      n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, 
      n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, 
      n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, 
      n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, 
      n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, 
      n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, 
      n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, 
      n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, 
      n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, 
      n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, 
      n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, 
      n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, 
      n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, 
      n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, 
      n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, 
      n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, 
      n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, 
      n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, 
      n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, 
      n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, 
      n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, 
      n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, 
      n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, 
      n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, 
      n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, 
      n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, 
      n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, 
      n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, 
      n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, 
      n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, 
      n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, 
      n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, 
      n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, 
      n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, 
      n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, 
      n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, 
      n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, 
      n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, 
      n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, 
      n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, 
      n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, 
      n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, 
      n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, 
      n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, 
      n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, 
      n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, 
      n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, 
      n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, 
      n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, 
      n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, 
      n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, 
      n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, 
      n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, 
      n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, 
      n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, 
      n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, 
      n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, 
      n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, 
      n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, 
      n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, 
      n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, 
      n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, 
      n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, 
      n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, 
      n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, 
      n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, 
      n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, 
      n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, 
      n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, 
      n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, 
      n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, 
      n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, 
      n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, 
      n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, 
      n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, 
      n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, 
      n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, 
      n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, 
      n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, 
      n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, 
      n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, 
      n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, 
      n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, 
      n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, 
      n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, 
      n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, 
      n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, 
      n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, 
      n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, 
      n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, 
      n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, 
      n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, 
      n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, 
      n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, 
      n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, 
      n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, 
      n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, 
      n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, 
      n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, 
      n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, 
      n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, 
      n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, 
      n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, 
      n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, 
      n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, 
      n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, 
      n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, 
      n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833, 
      n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842, 
      n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851, 
      n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860, 
      n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869, 
      n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878, 
      n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887, 
      n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896, 
      n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905, 
      n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914, 
      n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923, 
      n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932, 
      n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941, 
      n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950, 
      n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959, 
      n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968, 
      n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977, 
      n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986, 
      n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, 
      n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, 
      n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013, 
      n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022, 
      n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031, 
      n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040, 
      n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049, 
      n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058, 
      n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067, 
      n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076, 
      n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085, 
      n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, 
      n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, 
      n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, 
      n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, 
      n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130, 
      n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139, 
      n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148, 
      n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, 
      n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, 
      n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175, 
      n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184, 
      n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193, 
      n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, 
      n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, 
      n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220, 
      n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229, 
      n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238, 
      n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247, 
      n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256, 
      n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265, 
      n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274, 
      n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283, 
      n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292, 
      n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301, 
      n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310, 
      n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319, 
      n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328, 
      n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337, 
      n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346, 
      n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355, 
      n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364, 
      n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373, 
      n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382, 
      n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391, 
      n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400, 
      n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409, 
      n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418, 
      n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, 
      n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, 
      n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445, 
      n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454, 
      n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463, 
      n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472, 
      n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, 
      n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, 
      n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, 
      n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, 
      n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, 
      n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, 
      n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, 
      n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, 
      n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, 
      n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, 
      n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, 
      n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, 
      n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, 
      n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, 
      n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, 
      n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, 
      n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, 
      n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, 
      n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, 
      n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, 
      n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, 
      n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, 
      n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, 
      n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, 
      n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, 
      n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, 
      n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, 
      n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, 
      n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, 
      n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, 
      n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, 
      n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, 
      n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769, 
      n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778, 
      n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787, 
      n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796, 
      n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805, 
      n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814, 
      n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823, 
      n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832, 
      n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, 
      n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850, 
      n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859, 
      n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868, 
      n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877, 
      n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886, 
      n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895, 
      n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904, 
      n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913, 
      n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922, 
      n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931, 
      n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940, 
      n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949, 
      n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958, 
      n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967, 
      n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976, 
      n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985, 
      n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994, 
      n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003, 
      n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012, 
      n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021, 
      n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030, 
      n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039, 
      n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, 
      n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057, 
      n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066, 
      n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075, 
      n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, 
      n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, 
      n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, 
      n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, 
      n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120, 
      n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129, 
      n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, 
      n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, 
      n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, 
      n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165, 
      n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174, 
      n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183, 
      n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192, 
      n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201, 
      n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210, 
      n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219, 
      n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228, 
      n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237, 
      n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246, 
      n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255, 
      n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264, 
      n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273, 
      n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282, 
      n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291, 
      n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300, 
      n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309, 
      n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318, 
      n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327, 
      n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336, 
      n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345, 
      n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354, 
      n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363, 
      n41364, n41365, n41366, n41367, n41368, n41369, n41370, n_1000, n_1001, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, 
      n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, 
      n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, 
      n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, 
      n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, 
      n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, 
      n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, 
      n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, 
      n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, 
      n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, 
      n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, 
      n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, 
      n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, 
      n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, 
      n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, 
      n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, 
      n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, 
      n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, 
      n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, 
      n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, 
      n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, 
      n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, 
      n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, 
      n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, 
      n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, 
      n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, 
      n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, 
      n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, 
      n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, 
      n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, 
      n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, 
      n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, 
      n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, 
      n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, 
      n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, 
      n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, 
      n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, 
      n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, 
      n_2532, n_2533, n_2534, n_2535 : std_logic;

begin
   
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => 
                           n_1000, QN => n30481);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => 
                           n_1001, QN => n30482);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => 
                           n_1002, QN => n30483);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => 
                           n_1003, QN => n30484);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => 
                           n_1004, QN => n30485);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => 
                           n_1005, QN => n30486);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => 
                           n_1006, QN => n30487);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => 
                           n_1007, QN => n30488);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => 
                           n_1008, QN => n30489);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => 
                           n_1009, QN => n30490);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => 
                           n_1010, QN => n30491);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => 
                           n_1011, QN => n30492);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => 
                           n_1012, QN => n30493);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => 
                           n_1013, QN => n30494);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => 
                           n_1014, QN => n30495);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => 
                           n_1015, QN => n30496);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => 
                           n_1016, QN => n30497);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => 
                           n_1017, QN => n30498);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => 
                           n_1018, QN => n30499);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => 
                           n_1019, QN => n30500);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => 
                           n_1020, QN => n30501);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => 
                           n_1021, QN => n30502);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => 
                           n_1022, QN => n30503);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => 
                           n_1023, QN => n30504);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => 
                           n_1024, QN => n30505);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => 
                           n_1025, QN => n30506);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => 
                           n_1026, QN => n30507);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => 
                           n_1027, QN => n30508);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7487, CK => CLK, Q => 
                           n_1028, QN => n30509);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7488, CK => CLK, Q => 
                           n_1029, QN => n30510);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7489, CK => CLK, Q => 
                           n_1030, QN => n30511);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7490, CK => CLK, Q => 
                           n_1031, QN => n30512);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7491, CK => CLK, Q => 
                           n_1032, QN => n30513);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7492, CK => CLK, Q => 
                           n_1033, QN => n30514);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7493, CK => CLK, Q => 
                           n_1034, QN => n30515);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7494, CK => CLK, Q => 
                           n_1035, QN => n30516);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7495, CK => CLK, Q => 
                           n_1036, QN => n30517);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7496, CK => CLK, Q => 
                           n_1037, QN => n30518);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7497, CK => CLK, Q => 
                           n_1038, QN => n30519);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7498, CK => CLK, Q => 
                           n_1039, QN => n30520);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7499, CK => CLK, Q => 
                           n_1040, QN => n30521);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7500, CK => CLK, Q => 
                           n_1041, QN => n30522);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7501, CK => CLK, Q => 
                           n_1042, QN => n30523);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7502, CK => CLK, Q => 
                           n_1043, QN => n30524);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7503, CK => CLK, Q => 
                           n_1044, QN => n30525);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7504, CK => CLK, Q => 
                           n_1045, QN => n30526);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7505, CK => CLK, Q => 
                           n_1046, QN => n30527);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7506, CK => CLK, Q => 
                           n_1047, QN => n30528);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7507, CK => CLK, Q => 
                           n_1048, QN => n30529);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7508, CK => CLK, Q => 
                           n_1049, QN => n30530);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7509, CK => CLK, Q => 
                           n_1050, QN => n30531);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7510, CK => CLK, Q => 
                           n_1051, QN => n30532);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7511, CK => CLK, Q => 
                           n_1052, QN => n30533);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7512, CK => CLK, Q => 
                           n_1053, QN => n30534);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7513, CK => CLK, Q => n_1054
                           , QN => n30535);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7514, CK => CLK, Q => n_1055
                           , QN => n30536);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7515, CK => CLK, Q => n_1056
                           , QN => n30537);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7516, CK => CLK, Q => n_1057
                           , QN => n30538);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7517, CK => CLK, Q => n_1058
                           , QN => n30539);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7518, CK => CLK, Q => n_1059
                           , QN => n30540);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7523, CK => CLK, Q => 
                           n_1060, QN => n30545);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7524, CK => CLK, Q => 
                           n_1061, QN => n30546);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7525, CK => CLK, Q => 
                           n_1062, QN => n30547);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7527, CK => CLK, Q => 
                           n_1063, QN => n30549);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7547, CK => CLK, Q => 
                           n_1064, QN => n30569);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7548, CK => CLK, Q => 
                           n_1065, QN => n30570);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7549, CK => CLK, Q => 
                           n_1066, QN => n30571);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7550, CK => CLK, Q => 
                           n_1067, QN => n30572);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7551, CK => CLK, Q => 
                           n_1068, QN => n30573);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7552, CK => CLK, Q => 
                           n_1069, QN => n30574);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7553, CK => CLK, Q => 
                           n_1070, QN => n30575);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7554, CK => CLK, Q => 
                           n_1071, QN => n30576);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7555, CK => CLK, Q => 
                           n_1072, QN => n30577);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7556, CK => CLK, Q => 
                           n_1073, QN => n30578);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7557, CK => CLK, Q => 
                           n_1074, QN => n30579);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7558, CK => CLK, Q => 
                           n_1075, QN => n30580);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7559, CK => CLK, Q => 
                           n_1076, QN => n30581);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7560, CK => CLK, Q => 
                           n_1077, QN => n30582);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7561, CK => CLK, Q => 
                           n_1078, QN => n30583);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7562, CK => CLK, Q => 
                           n_1079, QN => n30584);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7563, CK => CLK, Q => 
                           n_1080, QN => n30585);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7564, CK => CLK, Q => 
                           n_1081, QN => n30586);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7565, CK => CLK, Q => 
                           n_1082, QN => n30587);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7566, CK => CLK, Q => 
                           n_1083, QN => n30588);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7567, CK => CLK, Q => 
                           n_1084, QN => n30589);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7568, CK => CLK, Q => 
                           n_1085, QN => n30590);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7569, CK => CLK, Q => 
                           n_1086, QN => n30591);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7570, CK => CLK, Q => 
                           n_1087, QN => n30592);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7571, CK => CLK, Q => 
                           n_1088, QN => n30593);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7572, CK => CLK, Q => 
                           n_1089, QN => n30594);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7573, CK => CLK, Q => 
                           n_1090, QN => n30595);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7574, CK => CLK, Q => 
                           n_1091, QN => n30596);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7575, CK => CLK, Q => 
                           n_1092, QN => n30597);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7576, CK => CLK, Q => 
                           n_1093, QN => n30598);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7577, CK => CLK, Q => n_1094
                           , QN => n30599);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7578, CK => CLK, Q => n_1095
                           , QN => n30600);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7579, CK => CLK, Q => n_1096
                           , QN => n30601);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7580, CK => CLK, Q => n_1097
                           , QN => n30602);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7581, CK => CLK, Q => n_1098
                           , QN => n30603);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7582, CK => CLK, Q => n_1099
                           , QN => n30604);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7587, CK => CLK, Q => 
                           n_1100, QN => n30609);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7588, CK => CLK, Q => 
                           n_1101, QN => n30610);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7589, CK => CLK, Q => 
                           n_1102, QN => n30611);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7590, CK => CLK, Q => 
                           n_1103, QN => n30612);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7591, CK => CLK, Q => 
                           n_1104, QN => n30613);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7592, CK => CLK, Q => 
                           n_1105, QN => n30614);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7593, CK => CLK, Q => 
                           n_1106, QN => n30615);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7594, CK => CLK, Q => 
                           n_1107, QN => n30616);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7595, CK => CLK, Q => 
                           n_1108, QN => n30617);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7596, CK => CLK, Q => 
                           n_1109, QN => n30618);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7597, CK => CLK, Q => 
                           n_1110, QN => n30619);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7598, CK => CLK, Q => 
                           n_1111, QN => n30620);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7599, CK => CLK, Q => 
                           n_1112, QN => n30621);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7600, CK => CLK, Q => 
                           n_1113, QN => n30622);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7601, CK => CLK, Q => 
                           n_1114, QN => n30623);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7602, CK => CLK, Q => 
                           n_1115, QN => n30624);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7603, CK => CLK, Q => 
                           n_1116, QN => n30625);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7604, CK => CLK, Q => 
                           n_1117, QN => n30626);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7605, CK => CLK, Q => 
                           n_1118, QN => n30627);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7606, CK => CLK, Q => 
                           n_1119, QN => n30628);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7607, CK => CLK, Q => 
                           n_1120, QN => n30629);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7608, CK => CLK, Q => 
                           n_1121, QN => n30630);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7609, CK => CLK, Q => 
                           n_1122, QN => n30631);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7610, CK => CLK, Q => 
                           n_1123, QN => n30632);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7611, CK => CLK, Q => 
                           n_1124, QN => n30633);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7612, CK => CLK, Q => 
                           n_1125, QN => n30634);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7613, CK => CLK, Q => 
                           n_1126, QN => n30635);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7614, CK => CLK, Q => 
                           n_1127, QN => n30636);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7615, CK => CLK, Q => 
                           n_1128, QN => n30637);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7616, CK => CLK, Q => 
                           n_1129, QN => n30638);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7617, CK => CLK, Q => 
                           n_1130, QN => n30639);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7618, CK => CLK, Q => 
                           n_1131, QN => n30640);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7619, CK => CLK, Q => 
                           n_1132, QN => n30641);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7620, CK => CLK, Q => 
                           n_1133, QN => n30642);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7621, CK => CLK, Q => 
                           n_1134, QN => n30643);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7622, CK => CLK, Q => 
                           n_1135, QN => n30644);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7623, CK => CLK, Q => 
                           n_1136, QN => n30645);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7624, CK => CLK, Q => 
                           n_1137, QN => n30646);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7625, CK => CLK, Q => 
                           n_1138, QN => n30647);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7626, CK => CLK, Q => 
                           n_1139, QN => n30648);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7627, CK => CLK, Q => 
                           n_1140, QN => n30649);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7628, CK => CLK, Q => 
                           n_1141, QN => n30650);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7629, CK => CLK, Q => 
                           n_1142, QN => n30651);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7630, CK => CLK, Q => 
                           n_1143, QN => n30652);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7631, CK => CLK, Q => 
                           n_1144, QN => n30653);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7632, CK => CLK, Q => 
                           n_1145, QN => n30654);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7633, CK => CLK, Q => 
                           n_1146, QN => n30655);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7634, CK => CLK, Q => 
                           n_1147, QN => n30656);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7635, CK => CLK, Q => 
                           n_1148, QN => n30657);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7636, CK => CLK, Q => 
                           n_1149, QN => n30658);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7637, CK => CLK, Q => 
                           n_1150, QN => n30659);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7638, CK => CLK, Q => 
                           n_1151, QN => n30660);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7639, CK => CLK, Q => 
                           n_1152, QN => n30661);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7640, CK => CLK, Q => 
                           n_1153, QN => n30662);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7641, CK => CLK, Q => n_1154
                           , QN => n30663);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7642, CK => CLK, Q => n_1155
                           , QN => n30664);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7643, CK => CLK, Q => n_1156
                           , QN => n30665);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7644, CK => CLK, Q => n_1157
                           , QN => n30666);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7645, CK => CLK, Q => n_1158
                           , QN => n30667);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7646, CK => CLK, Q => n_1159
                           , QN => n30668);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7779, CK => CLK, Q => 
                           n_1160, QN => n30673);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7780, CK => CLK, Q => 
                           n_1161, QN => n30674);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7781, CK => CLK, Q => 
                           n_1162, QN => n30675);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7782, CK => CLK, Q => 
                           n_1163, QN => n30676);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7783, CK => CLK, Q => 
                           n_1164, QN => n30677);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7784, CK => CLK, Q => 
                           n_1165, QN => n30678);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7785, CK => CLK, Q => 
                           n_1166, QN => n30679);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7786, CK => CLK, Q => 
                           n_1167, QN => n30680);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7787, CK => CLK, Q => 
                           n_1168, QN => n30681);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7788, CK => CLK, Q => 
                           n_1169, QN => n30682);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7789, CK => CLK, Q => 
                           n_1170, QN => n30683);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7790, CK => CLK, Q => 
                           n_1171, QN => n30684);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7791, CK => CLK, Q => 
                           n_1172, QN => n30685);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7792, CK => CLK, Q => 
                           n_1173, QN => n30686);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7793, CK => CLK, Q => 
                           n_1174, QN => n30687);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7794, CK => CLK, Q => 
                           n_1175, QN => n30688);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7795, CK => CLK, Q => 
                           n_1176, QN => n30689);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7796, CK => CLK, Q => 
                           n_1177, QN => n30690);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7797, CK => CLK, Q => 
                           n_1178, QN => n30691);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7798, CK => CLK, Q => 
                           n_1179, QN => n30692);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7799, CK => CLK, Q => 
                           n_1180, QN => n30693);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7800, CK => CLK, Q => 
                           n_1181, QN => n30694);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7801, CK => CLK, Q => 
                           n_1182, QN => n30695);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7802, CK => CLK, Q => 
                           n_1183, QN => n30696);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7803, CK => CLK, Q => 
                           n_1184, QN => n30697);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7804, CK => CLK, Q => 
                           n_1185, QN => n30698);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7805, CK => CLK, Q => 
                           n_1186, QN => n30699);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7806, CK => CLK, Q => 
                           n_1187, QN => n30700);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7807, CK => CLK, Q => 
                           n_1188, QN => n30701);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7808, CK => CLK, Q => 
                           n_1189, QN => n30702);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7809, CK => CLK, Q => 
                           n_1190, QN => n30703);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7810, CK => CLK, Q => 
                           n_1191, QN => n30704);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7811, CK => CLK, Q => 
                           n_1192, QN => n30705);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7812, CK => CLK, Q => 
                           n_1193, QN => n30706);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7813, CK => CLK, Q => 
                           n_1194, QN => n30707);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7814, CK => CLK, Q => 
                           n_1195, QN => n30708);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7815, CK => CLK, Q => 
                           n_1196, QN => n30709);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7816, CK => CLK, Q => 
                           n_1197, QN => n30710);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7817, CK => CLK, Q => 
                           n_1198, QN => n30711);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n7818, CK => CLK, Q => 
                           n_1199, QN => n30712);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n7819, CK => CLK, Q => 
                           n_1200, QN => n30713);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n7820, CK => CLK, Q => 
                           n_1201, QN => n30714);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n7821, CK => CLK, Q => 
                           n_1202, QN => n30715);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n7822, CK => CLK, Q => 
                           n_1203, QN => n30716);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n7823, CK => CLK, Q => 
                           n_1204, QN => n30717);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n7824, CK => CLK, Q => 
                           n_1205, QN => n30718);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n7825, CK => CLK, Q => 
                           n_1206, QN => n30719);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n7826, CK => CLK, Q => 
                           n_1207, QN => n30720);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n7827, CK => CLK, Q => 
                           n_1208, QN => n30721);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n7828, CK => CLK, Q => 
                           n_1209, QN => n30722);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n7829, CK => CLK, Q => 
                           n_1210, QN => n30723);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n7830, CK => CLK, Q => 
                           n_1211, QN => n30724);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n7831, CK => CLK, Q => 
                           n_1212, QN => n30725);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n7832, CK => CLK, Q => 
                           n_1213, QN => n30726);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n7833, CK => CLK, Q => n_1214
                           , QN => n30727);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n7834, CK => CLK, Q => n_1215
                           , QN => n30728);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n7835, CK => CLK, Q => n_1216
                           , QN => n30729);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n7836, CK => CLK, Q => n_1217
                           , QN => n30730);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n7837, CK => CLK, Q => n_1218
                           , QN => n30731);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n7838, CK => CLK, Q => n_1219
                           , QN => n30732);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n7843, CK => CLK, Q => 
                           n_1220, QN => n30737);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n7844, CK => CLK, Q => 
                           n_1221, QN => n30738);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n7845, CK => CLK, Q => 
                           n_1222, QN => n30739);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n7846, CK => CLK, Q => 
                           n_1223, QN => n30740);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n7847, CK => CLK, Q => 
                           n_1224, QN => n30741);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n7848, CK => CLK, Q => 
                           n_1225, QN => n30742);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n7849, CK => CLK, Q => 
                           n_1226, QN => n30743);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n7850, CK => CLK, Q => 
                           n_1227, QN => n30744);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n7851, CK => CLK, Q => 
                           n_1228, QN => n30745);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n7852, CK => CLK, Q => 
                           n_1229, QN => n30746);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n7853, CK => CLK, Q => 
                           n_1230, QN => n30747);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => 
                           n_1231, QN => n30748);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n7855, CK => CLK, Q => 
                           n_1232, QN => n30749);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n7856, CK => CLK, Q => 
                           n_1233, QN => n30750);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n7857, CK => CLK, Q => 
                           n_1234, QN => n30751);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n7858, CK => CLK, Q => 
                           n_1235, QN => n30752);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n7859, CK => CLK, Q => 
                           n_1236, QN => n30753);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n7860, CK => CLK, Q => 
                           n_1237, QN => n30754);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n7861, CK => CLK, Q => 
                           n_1238, QN => n30755);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n7862, CK => CLK, Q => 
                           n_1239, QN => n30756);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n7863, CK => CLK, Q => 
                           n_1240, QN => n30757);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n7864, CK => CLK, Q => 
                           n_1241, QN => n30758);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n7865, CK => CLK, Q => 
                           n_1242, QN => n30759);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n7866, CK => CLK, Q => 
                           n_1243, QN => n30760);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n7867, CK => CLK, Q => 
                           n_1244, QN => n30761);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n7868, CK => CLK, Q => 
                           n_1245, QN => n30762);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n7869, CK => CLK, Q => 
                           n_1246, QN => n30763);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n7870, CK => CLK, Q => 
                           n_1247, QN => n30764);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n7871, CK => CLK, Q => 
                           n_1248, QN => n30765);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n7872, CK => CLK, Q => 
                           n_1249, QN => n30766);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n7873, CK => CLK, Q => 
                           n_1250, QN => n30767);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n7874, CK => CLK, Q => 
                           n_1251, QN => n30768);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n7875, CK => CLK, Q => 
                           n_1252, QN => n30769);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n7876, CK => CLK, Q => 
                           n_1253, QN => n30770);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n7877, CK => CLK, Q => 
                           n_1254, QN => n30771);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n7878, CK => CLK, Q => 
                           n_1255, QN => n30772);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n7879, CK => CLK, Q => 
                           n_1256, QN => n30773);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n7880, CK => CLK, Q => 
                           n_1257, QN => n30774);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n7881, CK => CLK, Q => 
                           n_1258, QN => n30775);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n7882, CK => CLK, Q => 
                           n_1259, QN => n30776);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n7883, CK => CLK, Q => 
                           n_1260, QN => n30777);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n7884, CK => CLK, Q => 
                           n_1261, QN => n30778);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n7885, CK => CLK, Q => 
                           n_1262, QN => n30779);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n7886, CK => CLK, Q => 
                           n_1263, QN => n30780);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n7887, CK => CLK, Q => 
                           n_1264, QN => n30781);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n7888, CK => CLK, Q => 
                           n_1265, QN => n30782);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n7889, CK => CLK, Q => 
                           n_1266, QN => n30783);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n7890, CK => CLK, Q => 
                           n_1267, QN => n30784);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n7891, CK => CLK, Q => 
                           n_1268, QN => n30785);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n7892, CK => CLK, Q => 
                           n_1269, QN => n30786);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n7893, CK => CLK, Q => 
                           n_1270, QN => n30787);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n7894, CK => CLK, Q => 
                           n_1271, QN => n30788);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n7895, CK => CLK, Q => 
                           n_1272, QN => n30789);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n7896, CK => CLK, Q => 
                           n_1273, QN => n30790);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n7897, CK => CLK, Q => n_1274
                           , QN => n30791);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n7898, CK => CLK, Q => n_1275
                           , QN => n30792);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n7899, CK => CLK, Q => n_1276
                           , QN => n30793);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n7900, CK => CLK, Q => n_1277
                           , QN => n30794);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n7901, CK => CLK, Q => n_1278
                           , QN => n30795);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n7902, CK => CLK, Q => n_1279
                           , QN => n30796);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n7907, CK => CLK, Q => 
                           n_1280, QN => n30801);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n7908, CK => CLK, Q => 
                           n_1281, QN => n30802);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n7909, CK => CLK, Q => 
                           n_1282, QN => n30803);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n7910, CK => CLK, Q => 
                           n_1283, QN => n30804);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n7911, CK => CLK, Q => 
                           n_1284, QN => n30805);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n7912, CK => CLK, Q => 
                           n_1285, QN => n30806);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n7913, CK => CLK, Q => 
                           n_1286, QN => n30807);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n7914, CK => CLK, Q => 
                           n_1287, QN => n30808);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n7915, CK => CLK, Q => 
                           n_1288, QN => n30809);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n7916, CK => CLK, Q => 
                           n_1289, QN => n30810);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n7917, CK => CLK, Q => 
                           n_1290, QN => n30811);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n7918, CK => CLK, Q => 
                           n_1291, QN => n30812);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n7919, CK => CLK, Q => 
                           n_1292, QN => n30813);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n7920, CK => CLK, Q => 
                           n_1293, QN => n30814);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n7921, CK => CLK, Q => 
                           n_1294, QN => n30815);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n7922, CK => CLK, Q => 
                           n_1295, QN => n30816);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n7923, CK => CLK, Q => 
                           n_1296, QN => n30817);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n7924, CK => CLK, Q => 
                           n_1297, QN => n30818);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n7925, CK => CLK, Q => 
                           n_1298, QN => n30819);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n7926, CK => CLK, Q => 
                           n_1299, QN => n30820);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n7927, CK => CLK, Q => 
                           n_1300, QN => n30821);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n7928, CK => CLK, Q => 
                           n_1301, QN => n30822);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n7929, CK => CLK, Q => 
                           n_1302, QN => n30823);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n7930, CK => CLK, Q => 
                           n_1303, QN => n30824);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n7931, CK => CLK, Q => 
                           n_1304, QN => n30825);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n7932, CK => CLK, Q => 
                           n_1305, QN => n30826);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n7933, CK => CLK, Q => 
                           n_1306, QN => n30827);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n7934, CK => CLK, Q => 
                           n_1307, QN => n30828);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n7935, CK => CLK, Q => 
                           n_1308, QN => n30829);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n7936, CK => CLK, Q => 
                           n_1309, QN => n30830);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n7937, CK => CLK, Q => 
                           n_1310, QN => n30831);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n7938, CK => CLK, Q => 
                           n_1311, QN => n30832);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n7939, CK => CLK, Q => 
                           n_1312, QN => n30833);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n7940, CK => CLK, Q => 
                           n_1313, QN => n30834);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n7941, CK => CLK, Q => 
                           n_1314, QN => n30835);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n7942, CK => CLK, Q => 
                           n_1315, QN => n30836);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n7943, CK => CLK, Q => 
                           n_1316, QN => n30837);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n7944, CK => CLK, Q => 
                           n_1317, QN => n30838);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n7945, CK => CLK, Q => 
                           n_1318, QN => n30839);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n7946, CK => CLK, Q => 
                           n_1319, QN => n30840);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n7947, CK => CLK, Q => 
                           n_1320, QN => n30841);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n7948, CK => CLK, Q => 
                           n_1321, QN => n30842);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n7949, CK => CLK, Q => 
                           n_1322, QN => n30843);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n7950, CK => CLK, Q => 
                           n_1323, QN => n30844);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n7951, CK => CLK, Q => 
                           n_1324, QN => n30845);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n7952, CK => CLK, Q => 
                           n_1325, QN => n30846);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n7953, CK => CLK, Q => 
                           n_1326, QN => n30847);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n7954, CK => CLK, Q => 
                           n_1327, QN => n30848);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n7955, CK => CLK, Q => 
                           n_1328, QN => n30849);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n7956, CK => CLK, Q => 
                           n_1329, QN => n30850);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n7957, CK => CLK, Q => 
                           n_1330, QN => n30851);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n7958, CK => CLK, Q => 
                           n_1331, QN => n30852);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n7959, CK => CLK, Q => 
                           n_1332, QN => n30853);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n7960, CK => CLK, Q => 
                           n_1333, QN => n30854);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n7961, CK => CLK, Q => n_1334
                           , QN => n30855);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n7962, CK => CLK, Q => n_1335
                           , QN => n30856);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n7963, CK => CLK, Q => n_1336
                           , QN => n30857);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n7964, CK => CLK, Q => n_1337
                           , QN => n30858);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n7965, CK => CLK, Q => n_1338
                           , QN => n30859);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n7966, CK => CLK, Q => n_1339
                           , QN => n30860);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n8099, CK => CLK, Q => 
                           n_1340, QN => n30865);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n8100, CK => CLK, Q => 
                           n_1341, QN => n30866);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n8101, CK => CLK, Q => 
                           n_1342, QN => n30867);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n8102, CK => CLK, Q => 
                           n_1343, QN => n30868);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n8103, CK => CLK, Q => 
                           n_1344, QN => n30869);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n8104, CK => CLK, Q => 
                           n_1345, QN => n30870);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n8105, CK => CLK, Q => 
                           n_1346, QN => n30871);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n8106, CK => CLK, Q => 
                           n_1347, QN => n30872);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n8107, CK => CLK, Q => 
                           n_1348, QN => n30873);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n8108, CK => CLK, Q => 
                           n_1349, QN => n30874);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n8109, CK => CLK, Q => 
                           n_1350, QN => n30875);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n8110, CK => CLK, Q => 
                           n_1351, QN => n30876);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n8111, CK => CLK, Q => 
                           n_1352, QN => n30877);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n8112, CK => CLK, Q => 
                           n_1353, QN => n30878);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n8113, CK => CLK, Q => 
                           n_1354, QN => n30879);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n8114, CK => CLK, Q => 
                           n_1355, QN => n30880);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n8115, CK => CLK, Q => 
                           n_1356, QN => n30881);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n8116, CK => CLK, Q => 
                           n_1357, QN => n30882);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n8117, CK => CLK, Q => 
                           n_1358, QN => n30883);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n8118, CK => CLK, Q => 
                           n_1359, QN => n30884);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n8119, CK => CLK, Q => 
                           n_1360, QN => n30885);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n8120, CK => CLK, Q => 
                           n_1361, QN => n30886);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n8121, CK => CLK, Q => 
                           n_1362, QN => n30887);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n8122, CK => CLK, Q => 
                           n_1363, QN => n30888);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n8123, CK => CLK, Q => 
                           n_1364, QN => n30889);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n8124, CK => CLK, Q => 
                           n_1365, QN => n30890);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n8125, CK => CLK, Q => 
                           n_1366, QN => n30891);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n8126, CK => CLK, Q => 
                           n_1367, QN => n30892);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n8127, CK => CLK, Q => 
                           n_1368, QN => n30893);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n8128, CK => CLK, Q => 
                           n_1369, QN => n30894);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n8129, CK => CLK, Q => 
                           n_1370, QN => n30895);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n8130, CK => CLK, Q => 
                           n_1371, QN => n30896);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n8131, CK => CLK, Q => 
                           n_1372, QN => n30897);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n8132, CK => CLK, Q => 
                           n_1373, QN => n30898);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n8133, CK => CLK, Q => 
                           n_1374, QN => n30899);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n8134, CK => CLK, Q => 
                           n_1375, QN => n30900);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n8135, CK => CLK, Q => 
                           n_1376, QN => n30901);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n8136, CK => CLK, Q => 
                           n_1377, QN => n30902);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n8137, CK => CLK, Q => 
                           n_1378, QN => n30903);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n8138, CK => CLK, Q => 
                           n_1379, QN => n30904);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n8139, CK => CLK, Q => 
                           n_1380, QN => n30905);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n8140, CK => CLK, Q => 
                           n_1381, QN => n30906);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n8141, CK => CLK, Q => 
                           n_1382, QN => n30907);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n8142, CK => CLK, Q => 
                           n_1383, QN => n30908);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n8143, CK => CLK, Q => 
                           n_1384, QN => n30909);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n8144, CK => CLK, Q => 
                           n_1385, QN => n30910);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n8145, CK => CLK, Q => 
                           n_1386, QN => n30911);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n8146, CK => CLK, Q => 
                           n_1387, QN => n30912);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n8147, CK => CLK, Q => 
                           n_1388, QN => n30913);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n8148, CK => CLK, Q => 
                           n_1389, QN => n30914);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n8149, CK => CLK, Q => 
                           n_1390, QN => n30915);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n8150, CK => CLK, Q => 
                           n_1391, QN => n30916);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n8151, CK => CLK, Q => 
                           n_1392, QN => n30917);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n8152, CK => CLK, Q => 
                           n_1393, QN => n30918);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n8153, CK => CLK, Q => 
                           n_1394, QN => n30919);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n8154, CK => CLK, Q => 
                           n_1395, QN => n30920);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n8155, CK => CLK, Q => 
                           n_1396, QN => n30921);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n8156, CK => CLK, Q => 
                           n_1397, QN => n30922);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n8157, CK => CLK, Q => 
                           n_1398, QN => n30923);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n8158, CK => CLK, Q => 
                           n_1399, QN => n30924);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n8159, CK => CLK, Q => 
                           n_1400, QN => n30925);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n8160, CK => CLK, Q => 
                           n_1401, QN => n30926);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n8161, CK => CLK, Q => 
                           n_1402, QN => n30927);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n8162, CK => CLK, Q => 
                           n_1403, QN => n30928);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n8163, CK => CLK, Q => 
                           n_1404, QN => n30929);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n8164, CK => CLK, Q => 
                           n_1405, QN => n30930);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n8165, CK => CLK, Q => 
                           n_1406, QN => n30931);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n8166, CK => CLK, Q => 
                           n_1407, QN => n30932);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n8167, CK => CLK, Q => 
                           n_1408, QN => n30933);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n8168, CK => CLK, Q => 
                           n_1409, QN => n30934);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n8169, CK => CLK, Q => 
                           n_1410, QN => n30935);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n8170, CK => CLK, Q => 
                           n_1411, QN => n30936);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n8171, CK => CLK, Q => 
                           n_1412, QN => n30937);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n8172, CK => CLK, Q => 
                           n_1413, QN => n30938);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n8173, CK => CLK, Q => 
                           n_1414, QN => n30939);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n8174, CK => CLK, Q => 
                           n_1415, QN => n30940);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n8175, CK => CLK, Q => 
                           n_1416, QN => n30941);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n8176, CK => CLK, Q => 
                           n_1417, QN => n30942);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n8177, CK => CLK, Q => 
                           n_1418, QN => n30943);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n8178, CK => CLK, Q => 
                           n_1419, QN => n30944);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n8179, CK => CLK, Q => 
                           n_1420, QN => n30945);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n8180, CK => CLK, Q => 
                           n_1421, QN => n30946);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n8181, CK => CLK, Q => 
                           n_1422, QN => n30947);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n8182, CK => CLK, Q => 
                           n_1423, QN => n30948);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n8183, CK => CLK, Q => 
                           n_1424, QN => n30949);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n8184, CK => CLK, Q => 
                           n_1425, QN => n30950);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n8185, CK => CLK, Q => 
                           n_1426, QN => n30951);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n8186, CK => CLK, Q => 
                           n_1427, QN => n30952);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n8187, CK => CLK, Q => 
                           n_1428, QN => n30953);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n8188, CK => CLK, Q => 
                           n_1429, QN => n30954);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n8189, CK => CLK, Q => 
                           n_1430, QN => n30955);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n8190, CK => CLK, Q => 
                           n_1431, QN => n30956);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n8191, CK => CLK, Q => 
                           n_1432, QN => n30957);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n8192, CK => CLK, Q => 
                           n_1433, QN => n30958);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n8193, CK => CLK, Q => 
                           n_1434, QN => n30959);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n8194, CK => CLK, Q => 
                           n_1435, QN => n30960);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n8195, CK => CLK, Q => 
                           n_1436, QN => n30961);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n8196, CK => CLK, Q => 
                           n_1437, QN => n30962);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n8197, CK => CLK, Q => 
                           n_1438, QN => n30963);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n8198, CK => CLK, Q => 
                           n_1439, QN => n30964);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n8199, CK => CLK, Q => 
                           n_1440, QN => n30965);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n8200, CK => CLK, Q => 
                           n_1441, QN => n30966);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n8201, CK => CLK, Q => 
                           n_1442, QN => n30967);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n8202, CK => CLK, Q => 
                           n_1443, QN => n30968);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n8203, CK => CLK, Q => 
                           n_1444, QN => n30969);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n8204, CK => CLK, Q => 
                           n_1445, QN => n30970);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n8205, CK => CLK, Q => 
                           n_1446, QN => n30971);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n8206, CK => CLK, Q => 
                           n_1447, QN => n30972);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n8207, CK => CLK, Q => 
                           n_1448, QN => n30973);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n8208, CK => CLK, Q => 
                           n_1449, QN => n30974);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n8209, CK => CLK, Q => 
                           n_1450, QN => n30975);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n8210, CK => CLK, Q => 
                           n_1451, QN => n30976);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n8211, CK => CLK, Q => 
                           n_1452, QN => n30977);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n8212, CK => CLK, Q => 
                           n_1453, QN => n30978);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n8213, CK => CLK, Q => 
                           n_1454, QN => n30979);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n8214, CK => CLK, Q => 
                           n_1455, QN => n30980);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n8215, CK => CLK, Q => 
                           n_1456, QN => n30981);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n8216, CK => CLK, Q => 
                           n_1457, QN => n30982);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n8217, CK => CLK, Q => 
                           n_1458, QN => n30983);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n8218, CK => CLK, Q => 
                           n_1459, QN => n30984);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n8219, CK => CLK, Q => 
                           n_1460, QN => n30985);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n8220, CK => CLK, Q => 
                           n_1461, QN => n30986);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n8221, CK => CLK, Q => 
                           n_1462, QN => n30987);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n8222, CK => CLK, Q => 
                           n_1463, QN => n30988);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n8223, CK => CLK, Q => 
                           n_1464, QN => n30989);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n8224, CK => CLK, Q => 
                           n_1465, QN => n30990);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n8225, CK => CLK, Q => 
                           n_1466, QN => n30991);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n8226, CK => CLK, Q => 
                           n_1467, QN => n30992);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n8227, CK => CLK, Q => 
                           n_1468, QN => n30993);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n8228, CK => CLK, Q => 
                           n_1469, QN => n30994);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n8229, CK => CLK, Q => 
                           n_1470, QN => n30995);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n8230, CK => CLK, Q => 
                           n_1471, QN => n30996);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n8231, CK => CLK, Q => 
                           n_1472, QN => n30997);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n8232, CK => CLK, Q => 
                           n_1473, QN => n30998);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n8233, CK => CLK, Q => 
                           n_1474, QN => n30999);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n8234, CK => CLK, Q => 
                           n_1475, QN => n31000);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n8235, CK => CLK, Q => 
                           n_1476, QN => n31001);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n8236, CK => CLK, Q => 
                           n_1477, QN => n31002);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n8237, CK => CLK, Q => 
                           n_1478, QN => n31003);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n8238, CK => CLK, Q => 
                           n_1479, QN => n31004);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n8239, CK => CLK, Q => 
                           n_1480, QN => n31005);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n8240, CK => CLK, Q => 
                           n_1481, QN => n31006);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n8241, CK => CLK, Q => 
                           n_1482, QN => n31007);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n8242, CK => CLK, Q => 
                           n_1483, QN => n31008);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n8243, CK => CLK, Q => 
                           n_1484, QN => n31009);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n8244, CK => CLK, Q => 
                           n_1485, QN => n31010);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n8245, CK => CLK, Q => 
                           n_1486, QN => n31011);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n8246, CK => CLK, Q => 
                           n_1487, QN => n31012);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n8247, CK => CLK, Q => 
                           n_1488, QN => n31013);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n8248, CK => CLK, Q => 
                           n_1489, QN => n31014);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n8249, CK => CLK, Q => 
                           n_1490, QN => n31015);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n8250, CK => CLK, Q => 
                           n_1491, QN => n31016);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n8251, CK => CLK, Q => 
                           n_1492, QN => n31017);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n8252, CK => CLK, Q => 
                           n_1493, QN => n31018);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n8253, CK => CLK, Q => 
                           n_1494, QN => n31019);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n8254, CK => CLK, Q => 
                           n_1495, QN => n31020);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n8255, CK => CLK, Q => 
                           n_1496, QN => n31021);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n8256, CK => CLK, Q => 
                           n_1497, QN => n31022);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n8257, CK => CLK, Q => 
                           n_1498, QN => n31023);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n8258, CK => CLK, Q => 
                           n_1499, QN => n31024);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n8259, CK => CLK, Q => 
                           n_1500, QN => n31025);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n8260, CK => CLK, Q => 
                           n_1501, QN => n31026);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n8261, CK => CLK, Q => 
                           n_1502, QN => n31027);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n8262, CK => CLK, Q => 
                           n_1503, QN => n31028);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n8263, CK => CLK, Q => 
                           n_1504, QN => n31029);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n8264, CK => CLK, Q => 
                           n_1505, QN => n31030);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n8265, CK => CLK, Q => 
                           n_1506, QN => n31031);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n8266, CK => CLK, Q => 
                           n_1507, QN => n31032);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n8267, CK => CLK, Q => 
                           n_1508, QN => n31033);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n8268, CK => CLK, Q => 
                           n_1509, QN => n31034);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n8269, CK => CLK, Q => 
                           n_1510, QN => n31035);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n8270, CK => CLK, Q => 
                           n_1511, QN => n31036);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n8271, CK => CLK, Q => 
                           n_1512, QN => n31037);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n8272, CK => CLK, Q => 
                           n_1513, QN => n31038);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n8273, CK => CLK, Q => 
                           n_1514, QN => n31039);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n8274, CK => CLK, Q => 
                           n_1515, QN => n31040);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n8275, CK => CLK, Q => 
                           n_1516, QN => n31041);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n8276, CK => CLK, Q => 
                           n_1517, QN => n31042);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n8277, CK => CLK, Q => 
                           n_1518, QN => n31043);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n8278, CK => CLK, Q => 
                           n_1519, QN => n31044);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n8279, CK => CLK, Q => 
                           n_1520, QN => n31045);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n8280, CK => CLK, Q => 
                           n_1521, QN => n31046);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n8281, CK => CLK, Q => 
                           n_1522, QN => n31047);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n8282, CK => CLK, Q => 
                           n_1523, QN => n31048);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n8283, CK => CLK, Q => 
                           n_1524, QN => n31049);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n8284, CK => CLK, Q => 
                           n_1525, QN => n31050);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n8285, CK => CLK, Q => 
                           n_1526, QN => n31051);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n8286, CK => CLK, Q => 
                           n_1527, QN => n31052);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n8287, CK => CLK, Q => 
                           n_1528, QN => n31053);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n8288, CK => CLK, Q => 
                           n_1529, QN => n31054);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n8289, CK => CLK, Q => 
                           n_1530, QN => n31055);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n8290, CK => CLK, Q => 
                           n_1531, QN => n31056);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n8419, CK => CLK, Q => 
                           n_1532, QN => n31175);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n8420, CK => CLK, Q => 
                           n_1533, QN => n31176);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n8421, CK => CLK, Q => 
                           n_1534, QN => n31177);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n8422, CK => CLK, Q => 
                           n_1535, QN => n31178);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n8423, CK => CLK, Q => 
                           n_1536, QN => n31179);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n8424, CK => CLK, Q => 
                           n_1537, QN => n31180);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n8425, CK => CLK, Q => 
                           n_1538, QN => n31181);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n8426, CK => CLK, Q => 
                           n_1539, QN => n31182);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n8427, CK => CLK, Q => 
                           n_1540, QN => n31183);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n8428, CK => CLK, Q => 
                           n_1541, QN => n31184);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n8429, CK => CLK, Q => 
                           n_1542, QN => n31185);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n8430, CK => CLK, Q => 
                           n_1543, QN => n31186);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n8431, CK => CLK, Q => 
                           n_1544, QN => n31187);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n8432, CK => CLK, Q => 
                           n_1545, QN => n31188);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n8433, CK => CLK, Q => 
                           n_1546, QN => n31189);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n8434, CK => CLK, Q => 
                           n_1547, QN => n31190);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n8435, CK => CLK, Q => 
                           n_1548, QN => n31191);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n8436, CK => CLK, Q => 
                           n_1549, QN => n31192);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n8437, CK => CLK, Q => 
                           n_1550, QN => n31193);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n8438, CK => CLK, Q => 
                           n_1551, QN => n31194);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n8439, CK => CLK, Q => 
                           n_1552, QN => n31195);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n8440, CK => CLK, Q => 
                           n_1553, QN => n31196);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n8441, CK => CLK, Q => 
                           n_1554, QN => n31197);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n8442, CK => CLK, Q => 
                           n_1555, QN => n31198);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n8443, CK => CLK, Q => 
                           n_1556, QN => n31199);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n8444, CK => CLK, Q => 
                           n_1557, QN => n31200);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n8445, CK => CLK, Q => 
                           n_1558, QN => n31201);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n8446, CK => CLK, Q => 
                           n_1559, QN => n31202);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n8447, CK => CLK, Q => 
                           n_1560, QN => n31203);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n8448, CK => CLK, Q => 
                           n_1561, QN => n31204);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n8449, CK => CLK, Q => 
                           n_1562, QN => n31205);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n8450, CK => CLK, Q => 
                           n_1563, QN => n31206);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n8451, CK => CLK, Q => 
                           n_1564, QN => n31207);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n8452, CK => CLK, Q => 
                           n_1565, QN => n31208);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n8453, CK => CLK, Q => 
                           n_1566, QN => n31209);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n8454, CK => CLK, Q => 
                           n_1567, QN => n31210);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n8455, CK => CLK, Q => 
                           n_1568, QN => n31211);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n8456, CK => CLK, Q => 
                           n_1569, QN => n31212);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n8457, CK => CLK, Q => 
                           n_1570, QN => n31213);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n8458, CK => CLK, Q => 
                           n_1571, QN => n31214);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n8459, CK => CLK, Q => 
                           n_1572, QN => n31215);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n8460, CK => CLK, Q => 
                           n_1573, QN => n31216);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n8461, CK => CLK, Q => 
                           n_1574, QN => n31217);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n8462, CK => CLK, Q => 
                           n_1575, QN => n31218);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n8463, CK => CLK, Q => 
                           n_1576, QN => n31219);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n8464, CK => CLK, Q => 
                           n_1577, QN => n31220);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n8465, CK => CLK, Q => 
                           n_1578, QN => n31221);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n8466, CK => CLK, Q => 
                           n_1579, QN => n31222);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n8467, CK => CLK, Q => 
                           n_1580, QN => n31223);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n8468, CK => CLK, Q => 
                           n_1581, QN => n31224);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n8469, CK => CLK, Q => 
                           n_1582, QN => n31225);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n8470, CK => CLK, Q => 
                           n_1583, QN => n31226);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n8471, CK => CLK, Q => 
                           n_1584, QN => n31227);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n8472, CK => CLK, Q => 
                           n_1585, QN => n31228);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n8473, CK => CLK, Q => 
                           n_1586, QN => n31229);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n8474, CK => CLK, Q => 
                           n_1587, QN => n31230);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n8475, CK => CLK, Q => 
                           n_1588, QN => n31231);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n8476, CK => CLK, Q => 
                           n_1589, QN => n31232);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n8477, CK => CLK, Q => 
                           n_1590, QN => n31233);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n8478, CK => CLK, Q => 
                           n_1591, QN => n31234);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n8483, CK => CLK, Q => 
                           n_1592, QN => n31239);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n8484, CK => CLK, Q => 
                           n_1593, QN => n31240);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n8485, CK => CLK, Q => 
                           n_1594, QN => n31241);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n8486, CK => CLK, Q => 
                           n_1595, QN => n31242);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n8487, CK => CLK, Q => 
                           n_1596, QN => n31243);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n8488, CK => CLK, Q => 
                           n_1597, QN => n31244);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n8489, CK => CLK, Q => 
                           n_1598, QN => n31245);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n8490, CK => CLK, Q => 
                           n_1599, QN => n31246);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n8491, CK => CLK, Q => 
                           n_1600, QN => n31247);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n8492, CK => CLK, Q => 
                           n_1601, QN => n31248);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n8493, CK => CLK, Q => 
                           n_1602, QN => n31249);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n8494, CK => CLK, Q => 
                           n_1603, QN => n31250);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n8495, CK => CLK, Q => 
                           n_1604, QN => n31251);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n8496, CK => CLK, Q => 
                           n_1605, QN => n31252);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n8497, CK => CLK, Q => 
                           n_1606, QN => n31253);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n8498, CK => CLK, Q => 
                           n_1607, QN => n31254);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n8499, CK => CLK, Q => 
                           n_1608, QN => n31255);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n8500, CK => CLK, Q => 
                           n_1609, QN => n31256);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n8501, CK => CLK, Q => 
                           n_1610, QN => n31257);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n8502, CK => CLK, Q => 
                           n_1611, QN => n31258);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n8503, CK => CLK, Q => 
                           n_1612, QN => n31259);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n8504, CK => CLK, Q => 
                           n_1613, QN => n31260);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n8505, CK => CLK, Q => 
                           n_1614, QN => n31261);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n8506, CK => CLK, Q => 
                           n_1615, QN => n31262);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n8507, CK => CLK, Q => 
                           n_1616, QN => n31263);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n8508, CK => CLK, Q => 
                           n_1617, QN => n31264);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n8509, CK => CLK, Q => 
                           n_1618, QN => n31265);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n8510, CK => CLK, Q => 
                           n_1619, QN => n31266);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n8511, CK => CLK, Q => 
                           n_1620, QN => n31267);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n8512, CK => CLK, Q => 
                           n_1621, QN => n31268);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n8513, CK => CLK, Q => 
                           n_1622, QN => n31269);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n8514, CK => CLK, Q => 
                           n_1623, QN => n31270);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n8515, CK => CLK, Q => 
                           n_1624, QN => n31271);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n8516, CK => CLK, Q => 
                           n_1625, QN => n31272);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n8517, CK => CLK, Q => 
                           n_1626, QN => n31273);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n8518, CK => CLK, Q => 
                           n_1627, QN => n31274);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n8519, CK => CLK, Q => 
                           n_1628, QN => n31275);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n8520, CK => CLK, Q => 
                           n_1629, QN => n31276);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n8521, CK => CLK, Q => 
                           n_1630, QN => n31277);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n8522, CK => CLK, Q => 
                           n_1631, QN => n31278);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n8523, CK => CLK, Q => 
                           n_1632, QN => n31279);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n8524, CK => CLK, Q => 
                           n_1633, QN => n31280);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n8525, CK => CLK, Q => 
                           n_1634, QN => n31281);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n8526, CK => CLK, Q => 
                           n_1635, QN => n31282);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n8527, CK => CLK, Q => 
                           n_1636, QN => n31283);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n8528, CK => CLK, Q => 
                           n_1637, QN => n31284);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n8529, CK => CLK, Q => 
                           n_1638, QN => n31285);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n8530, CK => CLK, Q => 
                           n_1639, QN => n31286);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n8531, CK => CLK, Q => 
                           n_1640, QN => n31287);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n8532, CK => CLK, Q => 
                           n_1641, QN => n31288);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n8533, CK => CLK, Q => 
                           n_1642, QN => n31289);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n8534, CK => CLK, Q => 
                           n_1643, QN => n31290);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n8535, CK => CLK, Q => 
                           n_1644, QN => n31291);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n8536, CK => CLK, Q => 
                           n_1645, QN => n31292);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n8537, CK => CLK, Q => 
                           n_1646, QN => n31293);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n8538, CK => CLK, Q => 
                           n_1647, QN => n31294);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n8539, CK => CLK, Q => 
                           n_1648, QN => n31295);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n8540, CK => CLK, Q => 
                           n_1649, QN => n31296);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n8541, CK => CLK, Q => 
                           n_1650, QN => n31297);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n8542, CK => CLK, Q => 
                           n_1651, QN => n31298);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n8547, CK => CLK, Q => 
                           n_1652, QN => n31303);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n8548, CK => CLK, Q => 
                           n_1653, QN => n31304);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n8549, CK => CLK, Q => 
                           n_1654, QN => n31305);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n8550, CK => CLK, Q => 
                           n_1655, QN => n31306);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n8551, CK => CLK, Q => 
                           n_1656, QN => n31307);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n8552, CK => CLK, Q => 
                           n_1657, QN => n31308);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n8553, CK => CLK, Q => 
                           n_1658, QN => n31309);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n8554, CK => CLK, Q => 
                           n_1659, QN => n31310);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n8555, CK => CLK, Q => 
                           n_1660, QN => n31311);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n8556, CK => CLK, Q => 
                           n_1661, QN => n31312);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n8557, CK => CLK, Q => 
                           n_1662, QN => n31313);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n8558, CK => CLK, Q => 
                           n_1663, QN => n31314);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n8559, CK => CLK, Q => 
                           n_1664, QN => n31315);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n8560, CK => CLK, Q => 
                           n_1665, QN => n31316);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n8561, CK => CLK, Q => 
                           n_1666, QN => n31317);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n8562, CK => CLK, Q => 
                           n_1667, QN => n31318);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n8563, CK => CLK, Q => 
                           n_1668, QN => n31319);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n8564, CK => CLK, Q => 
                           n_1669, QN => n31320);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n8565, CK => CLK, Q => 
                           n_1670, QN => n31321);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n8566, CK => CLK, Q => 
                           n_1671, QN => n31322);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n8567, CK => CLK, Q => 
                           n_1672, QN => n31323);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n8568, CK => CLK, Q => 
                           n_1673, QN => n31324);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n8569, CK => CLK, Q => 
                           n_1674, QN => n31325);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n8570, CK => CLK, Q => 
                           n_1675, QN => n31326);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n8571, CK => CLK, Q => 
                           n_1676, QN => n31327);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n8572, CK => CLK, Q => 
                           n_1677, QN => n31328);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n8573, CK => CLK, Q => 
                           n_1678, QN => n31329);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n8574, CK => CLK, Q => 
                           n_1679, QN => n31330);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n8575, CK => CLK, Q => 
                           n_1680, QN => n31331);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n8576, CK => CLK, Q => 
                           n_1681, QN => n31332);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n8577, CK => CLK, Q => 
                           n_1682, QN => n31333);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n8578, CK => CLK, Q => 
                           n_1683, QN => n31334);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n8579, CK => CLK, Q => 
                           n_1684, QN => n31335);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n8580, CK => CLK, Q => 
                           n_1685, QN => n31336);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n8581, CK => CLK, Q => 
                           n_1686, QN => n31337);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n8582, CK => CLK, Q => 
                           n_1687, QN => n31338);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n8583, CK => CLK, Q => 
                           n_1688, QN => n31339);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n8584, CK => CLK, Q => 
                           n_1689, QN => n31340);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n8585, CK => CLK, Q => 
                           n_1690, QN => n31341);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n8586, CK => CLK, Q => 
                           n_1691, QN => n31342);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n8587, CK => CLK, Q => 
                           n_1692, QN => n31343);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n8588, CK => CLK, Q => 
                           n_1693, QN => n31344);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n8589, CK => CLK, Q => 
                           n_1694, QN => n31345);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n8590, CK => CLK, Q => 
                           n_1695, QN => n31346);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n8591, CK => CLK, Q => 
                           n_1696, QN => n31347);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n8592, CK => CLK, Q => 
                           n_1697, QN => n31348);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n8593, CK => CLK, Q => 
                           n_1698, QN => n31349);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n8594, CK => CLK, Q => 
                           n_1699, QN => n31350);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n8595, CK => CLK, Q => 
                           n_1700, QN => n31351);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n8596, CK => CLK, Q => 
                           n_1701, QN => n31352);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n8597, CK => CLK, Q => 
                           n_1702, QN => n31353);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n8598, CK => CLK, Q => 
                           n_1703, QN => n31354);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n8599, CK => CLK, Q => 
                           n_1704, QN => n31355);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n8600, CK => CLK, Q => 
                           n_1705, QN => n31356);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n8601, CK => CLK, Q => 
                           n_1706, QN => n31357);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n8602, CK => CLK, Q => 
                           n_1707, QN => n31358);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n8603, CK => CLK, Q => 
                           n_1708, QN => n31359);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n8604, CK => CLK, Q => 
                           n_1709, QN => n31360);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n8605, CK => CLK, Q => 
                           n_1710, QN => n31361);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n8606, CK => CLK, Q => 
                           n_1711, QN => n31362);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n8739, CK => CLK, Q => 
                           n_1712, QN => n31367);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n8740, CK => CLK, Q => 
                           n_1713, QN => n31368);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n8741, CK => CLK, Q => 
                           n_1714, QN => n31369);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n8742, CK => CLK, Q => 
                           n_1715, QN => n31370);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n8743, CK => CLK, Q => 
                           n_1716, QN => n31371);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n8744, CK => CLK, Q => 
                           n_1717, QN => n31372);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n8745, CK => CLK, Q => 
                           n_1718, QN => n31373);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n8746, CK => CLK, Q => 
                           n_1719, QN => n31374);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n8747, CK => CLK, Q => 
                           n_1720, QN => n31375);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n8748, CK => CLK, Q => 
                           n_1721, QN => n31376);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n8749, CK => CLK, Q => 
                           n_1722, QN => n31377);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n8750, CK => CLK, Q => 
                           n_1723, QN => n31378);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n8751, CK => CLK, Q => 
                           n_1724, QN => n31379);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n8752, CK => CLK, Q => 
                           n_1725, QN => n31380);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n8753, CK => CLK, Q => 
                           n_1726, QN => n31381);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n8754, CK => CLK, Q => 
                           n_1727, QN => n31382);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n8755, CK => CLK, Q => 
                           n_1728, QN => n31383);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n8756, CK => CLK, Q => 
                           n_1729, QN => n31384);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n8757, CK => CLK, Q => 
                           n_1730, QN => n31385);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n8758, CK => CLK, Q => 
                           n_1731, QN => n31386);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n8759, CK => CLK, Q => 
                           n_1732, QN => n31387);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n8760, CK => CLK, Q => 
                           n_1733, QN => n31388);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n8761, CK => CLK, Q => 
                           n_1734, QN => n31389);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n8762, CK => CLK, Q => 
                           n_1735, QN => n31390);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n8763, CK => CLK, Q => 
                           n_1736, QN => n31391);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n8764, CK => CLK, Q => 
                           n_1737, QN => n31392);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n8765, CK => CLK, Q => 
                           n_1738, QN => n31393);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n8766, CK => CLK, Q => 
                           n_1739, QN => n31394);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n8767, CK => CLK, Q => 
                           n_1740, QN => n31395);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n8768, CK => CLK, Q => 
                           n_1741, QN => n31396);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n8769, CK => CLK, Q => 
                           n_1742, QN => n31397);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n8770, CK => CLK, Q => 
                           n_1743, QN => n31398);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n8771, CK => CLK, Q => 
                           n_1744, QN => n31399);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n8772, CK => CLK, Q => 
                           n_1745, QN => n31400);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n8773, CK => CLK, Q => 
                           n_1746, QN => n31401);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n8774, CK => CLK, Q => 
                           n_1747, QN => n31402);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n8775, CK => CLK, Q => 
                           n_1748, QN => n31403);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n8776, CK => CLK, Q => 
                           n_1749, QN => n31404);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n8777, CK => CLK, Q => 
                           n_1750, QN => n31405);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n8778, CK => CLK, Q => 
                           n_1751, QN => n31406);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n8779, CK => CLK, Q => 
                           n_1752, QN => n31407);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n8780, CK => CLK, Q => 
                           n_1753, QN => n31408);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n8781, CK => CLK, Q => 
                           n_1754, QN => n31409);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n8782, CK => CLK, Q => 
                           n_1755, QN => n31410);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n8783, CK => CLK, Q => 
                           n_1756, QN => n31411);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n8784, CK => CLK, Q => 
                           n_1757, QN => n31412);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n8785, CK => CLK, Q => 
                           n_1758, QN => n31413);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n8786, CK => CLK, Q => 
                           n_1759, QN => n31414);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n8787, CK => CLK, Q => 
                           n_1760, QN => n31415);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n8788, CK => CLK, Q => 
                           n_1761, QN => n31416);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n8789, CK => CLK, Q => 
                           n_1762, QN => n31417);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n8790, CK => CLK, Q => 
                           n_1763, QN => n31418);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n8791, CK => CLK, Q => 
                           n_1764, QN => n31419);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n8792, CK => CLK, Q => 
                           n_1765, QN => n31420);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n8793, CK => CLK, Q => 
                           n_1766, QN => n31421);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n8794, CK => CLK, Q => 
                           n_1767, QN => n31422);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n8795, CK => CLK, Q => 
                           n_1768, QN => n31423);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n8796, CK => CLK, Q => 
                           n_1769, QN => n31424);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n8797, CK => CLK, Q => 
                           n_1770, QN => n31425);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n8798, CK => CLK, Q => 
                           n_1771, QN => n31426);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n8799, CK => CLK, Q => 
                           n_1772, QN => n31427);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n8800, CK => CLK, Q => 
                           n_1773, QN => n31428);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n8801, CK => CLK, Q => 
                           n_1774, QN => n31429);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n8802, CK => CLK, Q => 
                           n_1775, QN => n31430);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n8803, CK => CLK, Q => 
                           n_1776, QN => n31431);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n8804, CK => CLK, Q => 
                           n_1777, QN => n31432);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n8805, CK => CLK, Q => 
                           n_1778, QN => n31433);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n8806, CK => CLK, Q => 
                           n_1779, QN => n31434);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n8807, CK => CLK, Q => 
                           n_1780, QN => n31435);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n8808, CK => CLK, Q => 
                           n_1781, QN => n31436);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n8809, CK => CLK, Q => 
                           n_1782, QN => n31437);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n8810, CK => CLK, Q => 
                           n_1783, QN => n31438);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n8811, CK => CLK, Q => 
                           n_1784, QN => n31439);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n8812, CK => CLK, Q => 
                           n_1785, QN => n31440);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n8813, CK => CLK, Q => 
                           n_1786, QN => n31441);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n8814, CK => CLK, Q => 
                           n_1787, QN => n31442);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n8815, CK => CLK, Q => 
                           n_1788, QN => n31443);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n8816, CK => CLK, Q => 
                           n_1789, QN => n31444);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n8817, CK => CLK, Q => 
                           n_1790, QN => n31445);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n8818, CK => CLK, Q => 
                           n_1791, QN => n31446);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n8819, CK => CLK, Q => 
                           n_1792, QN => n31447);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n8820, CK => CLK, Q => 
                           n_1793, QN => n31448);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n8821, CK => CLK, Q => 
                           n_1794, QN => n31449);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n8822, CK => CLK, Q => 
                           n_1795, QN => n31450);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n8823, CK => CLK, Q => 
                           n_1796, QN => n31451);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n8824, CK => CLK, Q => 
                           n_1797, QN => n31452);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n8825, CK => CLK, Q => 
                           n_1798, QN => n31453);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n8826, CK => CLK, Q => 
                           n_1799, QN => n31454);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n8827, CK => CLK, Q => 
                           n_1800, QN => n31455);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n8828, CK => CLK, Q => 
                           n_1801, QN => n31456);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n8829, CK => CLK, Q => 
                           n_1802, QN => n31457);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n8830, CK => CLK, Q => 
                           n_1803, QN => n31458);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n8831, CK => CLK, Q => 
                           n_1804, QN => n31459);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n8832, CK => CLK, Q => 
                           n_1805, QN => n31460);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n8833, CK => CLK, Q => 
                           n_1806, QN => n31461);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n8834, CK => CLK, Q => 
                           n_1807, QN => n31462);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n8835, CK => CLK, Q => 
                           n_1808, QN => n31463);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n8836, CK => CLK, Q => 
                           n_1809, QN => n31464);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n8837, CK => CLK, Q => 
                           n_1810, QN => n31465);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n8838, CK => CLK, Q => 
                           n_1811, QN => n31466);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n8839, CK => CLK, Q => 
                           n_1812, QN => n31467);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n8840, CK => CLK, Q => 
                           n_1813, QN => n31468);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n8841, CK => CLK, Q => 
                           n_1814, QN => n31469);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n8842, CK => CLK, Q => 
                           n_1815, QN => n31470);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n8843, CK => CLK, Q => 
                           n_1816, QN => n31471);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n8844, CK => CLK, Q => 
                           n_1817, QN => n31472);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n8845, CK => CLK, Q => 
                           n_1818, QN => n31473);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n8846, CK => CLK, Q => 
                           n_1819, QN => n31474);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n8847, CK => CLK, Q => 
                           n_1820, QN => n31475);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n8848, CK => CLK, Q => 
                           n_1821, QN => n31476);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n8849, CK => CLK, Q => 
                           n_1822, QN => n31477);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n8850, CK => CLK, Q => 
                           n_1823, QN => n31478);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n8851, CK => CLK, Q => 
                           n_1824, QN => n31479);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n8852, CK => CLK, Q => 
                           n_1825, QN => n31480);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n8853, CK => CLK, Q => 
                           n_1826, QN => n31481);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n8854, CK => CLK, Q => 
                           n_1827, QN => n31482);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n8855, CK => CLK, Q => 
                           n_1828, QN => n31483);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n8856, CK => CLK, Q => 
                           n_1829, QN => n31484);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n8857, CK => CLK, Q => 
                           n_1830, QN => n31485);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n8858, CK => CLK, Q => 
                           n_1831, QN => n31486);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n8859, CK => CLK, Q => 
                           n_1832, QN => n31487);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n8860, CK => CLK, Q => 
                           n_1833, QN => n31488);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n8861, CK => CLK, Q => 
                           n_1834, QN => n31489);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n8862, CK => CLK, Q => 
                           n_1835, QN => n31490);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n8863, CK => CLK, Q => 
                           n_1836, QN => n31491);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n8864, CK => CLK, Q => 
                           n_1837, QN => n31492);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n8865, CK => CLK, Q => 
                           n_1838, QN => n31493);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n8866, CK => CLK, Q => 
                           n_1839, QN => n31494);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n8867, CK => CLK, Q => 
                           n_1840, QN => n31495);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n8868, CK => CLK, Q => 
                           n_1841, QN => n31496);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n8869, CK => CLK, Q => 
                           n_1842, QN => n31497);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n8870, CK => CLK, Q => 
                           n_1843, QN => n31498);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n8871, CK => CLK, Q => 
                           n_1844, QN => n31499);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n8872, CK => CLK, Q => 
                           n_1845, QN => n31500);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n8873, CK => CLK, Q => 
                           n_1846, QN => n31501);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n8874, CK => CLK, Q => 
                           n_1847, QN => n31502);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n8875, CK => CLK, Q => 
                           n_1848, QN => n31503);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n8876, CK => CLK, Q => 
                           n_1849, QN => n31504);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n8877, CK => CLK, Q => 
                           n_1850, QN => n31505);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n8878, CK => CLK, Q => 
                           n_1851, QN => n31506);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n8879, CK => CLK, Q => 
                           n_1852, QN => n31507);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n8880, CK => CLK, Q => 
                           n_1853, QN => n31508);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n8881, CK => CLK, Q => 
                           n_1854, QN => n31509);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n8882, CK => CLK, Q => 
                           n_1855, QN => n31510);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n8883, CK => CLK, Q => 
                           n_1856, QN => n31511);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n8884, CK => CLK, Q => 
                           n_1857, QN => n31512);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n8885, CK => CLK, Q => 
                           n_1858, QN => n31513);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n8886, CK => CLK, Q => 
                           n_1859, QN => n31514);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n8887, CK => CLK, Q => 
                           n_1860, QN => n31515);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n8888, CK => CLK, Q => 
                           n_1861, QN => n31516);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n8889, CK => CLK, Q => 
                           n_1862, QN => n31517);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n8890, CK => CLK, Q => 
                           n_1863, QN => n31518);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n8891, CK => CLK, Q => 
                           n_1864, QN => n31519);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n8892, CK => CLK, Q => 
                           n_1865, QN => n31520);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n8893, CK => CLK, Q => 
                           n_1866, QN => n31521);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n8894, CK => CLK, Q => 
                           n_1867, QN => n31522);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n8895, CK => CLK, Q => 
                           n_1868, QN => n31523);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n8896, CK => CLK, Q => 
                           n_1869, QN => n31524);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n8897, CK => CLK, Q => 
                           n_1870, QN => n31525);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n8898, CK => CLK, Q => 
                           n_1871, QN => n31526);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n8899, CK => CLK, Q => 
                           n_1872, QN => n31527);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n8900, CK => CLK, Q => 
                           n_1873, QN => n31528);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n8901, CK => CLK, Q => 
                           n_1874, QN => n31529);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n8902, CK => CLK, Q => 
                           n_1875, QN => n31530);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n8903, CK => CLK, Q => 
                           n_1876, QN => n31531);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n8904, CK => CLK, Q => 
                           n_1877, QN => n31532);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n8905, CK => CLK, Q => 
                           n_1878, QN => n31533);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n8906, CK => CLK, Q => 
                           n_1879, QN => n31534);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n8907, CK => CLK, Q => 
                           n_1880, QN => n31535);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n8908, CK => CLK, Q => 
                           n_1881, QN => n31536);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n8909, CK => CLK, Q => 
                           n_1882, QN => n31537);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n8910, CK => CLK, Q => 
                           n_1883, QN => n31538);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n8911, CK => CLK, Q => 
                           n_1884, QN => n31539);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n8912, CK => CLK, Q => 
                           n_1885, QN => n31540);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n8913, CK => CLK, Q => 
                           n_1886, QN => n31541);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n8914, CK => CLK, Q => 
                           n_1887, QN => n31542);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n8915, CK => CLK, Q => 
                           n_1888, QN => n31543);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n8916, CK => CLK, Q => 
                           n_1889, QN => n31544);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n8917, CK => CLK, Q => 
                           n_1890, QN => n31545);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n8918, CK => CLK, Q => 
                           n_1891, QN => n31546);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n8919, CK => CLK, Q => 
                           n_1892, QN => n31547);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n8920, CK => CLK, Q => 
                           n_1893, QN => n31548);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n8921, CK => CLK, Q => 
                           n_1894, QN => n31549);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n8922, CK => CLK, Q => 
                           n_1895, QN => n31550);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n8923, CK => CLK, Q => 
                           n_1896, QN => n31551);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n8924, CK => CLK, Q => 
                           n_1897, QN => n31552);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n8925, CK => CLK, Q => 
                           n_1898, QN => n31553);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n8926, CK => CLK, Q => 
                           n_1899, QN => n31554);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n8927, CK => CLK, Q => 
                           n_1900, QN => n31555);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n8928, CK => CLK, Q => 
                           n_1901, QN => n31556);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n8929, CK => CLK, Q => 
                           n_1902, QN => n31557);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n8930, CK => CLK, Q => 
                           n_1903, QN => n31558);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n9059, CK => CLK, Q => 
                           n_1904, QN => n31559);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n9060, CK => CLK, Q => 
                           n_1905, QN => n31560);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n9061, CK => CLK, Q => 
                           n_1906, QN => n31561);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n9062, CK => CLK, Q => 
                           n_1907, QN => n31562);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n9063, CK => CLK, Q => 
                           n_1908, QN => n31563);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n9064, CK => CLK, Q => 
                           n_1909, QN => n31564);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n9065, CK => CLK, Q => 
                           n_1910, QN => n31565);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n9066, CK => CLK, Q => 
                           n_1911, QN => n31566);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n9067, CK => CLK, Q => 
                           n_1912, QN => n31567);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n9068, CK => CLK, Q => 
                           n_1913, QN => n31568);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n9069, CK => CLK, Q => 
                           n_1914, QN => n31569);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n9070, CK => CLK, Q => 
                           n_1915, QN => n31570);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n9071, CK => CLK, Q => 
                           n_1916, QN => n31571);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n9072, CK => CLK, Q => 
                           n_1917, QN => n31572);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n9073, CK => CLK, Q => 
                           n_1918, QN => n31573);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n9074, CK => CLK, Q => 
                           n_1919, QN => n31574);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n9075, CK => CLK, Q => 
                           n_1920, QN => n31575);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n9076, CK => CLK, Q => 
                           n_1921, QN => n31576);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n9077, CK => CLK, Q => 
                           n_1922, QN => n31577);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n9078, CK => CLK, Q => 
                           n_1923, QN => n31578);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n9079, CK => CLK, Q => 
                           n_1924, QN => n31579);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n9080, CK => CLK, Q => 
                           n_1925, QN => n31580);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n9081, CK => CLK, Q => 
                           n_1926, QN => n31581);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n9082, CK => CLK, Q => 
                           n_1927, QN => n31582);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n9083, CK => CLK, Q => 
                           n_1928, QN => n31583);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n9084, CK => CLK, Q => 
                           n_1929, QN => n31584);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n9085, CK => CLK, Q => 
                           n_1930, QN => n31585);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n9086, CK => CLK, Q => 
                           n_1931, QN => n31586);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n9087, CK => CLK, Q => 
                           n_1932, QN => n31587);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n9088, CK => CLK, Q => 
                           n_1933, QN => n31588);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n9089, CK => CLK, Q => 
                           n_1934, QN => n31589);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n9090, CK => CLK, Q => 
                           n_1935, QN => n31590);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n9091, CK => CLK, Q => 
                           n_1936, QN => n31591);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n9092, CK => CLK, Q => 
                           n_1937, QN => n31592);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n9093, CK => CLK, Q => 
                           n_1938, QN => n31593);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n9094, CK => CLK, Q => 
                           n_1939, QN => n31594);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n9095, CK => CLK, Q => 
                           n_1940, QN => n31595);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n9096, CK => CLK, Q => 
                           n_1941, QN => n31596);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n9097, CK => CLK, Q => 
                           n_1942, QN => n31597);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n9098, CK => CLK, Q => 
                           n_1943, QN => n31598);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n9099, CK => CLK, Q => 
                           n_1944, QN => n31599);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n9100, CK => CLK, Q => 
                           n_1945, QN => n31600);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n9101, CK => CLK, Q => 
                           n_1946, QN => n31601);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n9102, CK => CLK, Q => 
                           n_1947, QN => n31602);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n9103, CK => CLK, Q => 
                           n_1948, QN => n31603);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n9104, CK => CLK, Q => 
                           n_1949, QN => n31604);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n9105, CK => CLK, Q => 
                           n_1950, QN => n31605);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n9106, CK => CLK, Q => 
                           n_1951, QN => n31606);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n9107, CK => CLK, Q => 
                           n_1952, QN => n31607);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n9108, CK => CLK, Q => 
                           n_1953, QN => n31608);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n9109, CK => CLK, Q => 
                           n_1954, QN => n31609);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n9110, CK => CLK, Q => 
                           n_1955, QN => n31610);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n9111, CK => CLK, Q => 
                           n_1956, QN => n31611);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n9112, CK => CLK, Q => 
                           n_1957, QN => n31612);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n9113, CK => CLK, Q => 
                           n_1958, QN => n31613);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n9114, CK => CLK, Q => 
                           n_1959, QN => n31614);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n9115, CK => CLK, Q => 
                           n_1960, QN => n31615);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n9116, CK => CLK, Q => 
                           n_1961, QN => n31616);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n9117, CK => CLK, Q => 
                           n_1962, QN => n31617);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n9118, CK => CLK, Q => 
                           n_1963, QN => n31618);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n9119, CK => CLK, Q => 
                           n_1964, QN => n31619);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n9120, CK => CLK, Q => 
                           n_1965, QN => n31620);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n9121, CK => CLK, Q => 
                           n_1966, QN => n31621);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n9122, CK => CLK, Q => 
                           n_1967, QN => n31622);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n9123, CK => CLK, Q => 
                           n_1968, QN => n31623);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n9124, CK => CLK, Q => 
                           n_1969, QN => n31624);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n9125, CK => CLK, Q => 
                           n_1970, QN => n31625);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n9126, CK => CLK, Q => 
                           n_1971, QN => n31626);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n9127, CK => CLK, Q => 
                           n_1972, QN => n31627);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n9128, CK => CLK, Q => 
                           n_1973, QN => n31628);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n9129, CK => CLK, Q => 
                           n_1974, QN => n31629);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n9130, CK => CLK, Q => 
                           n_1975, QN => n31630);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n9131, CK => CLK, Q => 
                           n_1976, QN => n31631);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n9132, CK => CLK, Q => 
                           n_1977, QN => n31632);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n9133, CK => CLK, Q => 
                           n_1978, QN => n31633);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n9134, CK => CLK, Q => 
                           n_1979, QN => n31634);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n9135, CK => CLK, Q => 
                           n_1980, QN => n31635);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n9136, CK => CLK, Q => 
                           n_1981, QN => n31636);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n9137, CK => CLK, Q => 
                           n_1982, QN => n31637);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n9138, CK => CLK, Q => 
                           n_1983, QN => n31638);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n9139, CK => CLK, Q => 
                           n_1984, QN => n31639);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n9140, CK => CLK, Q => 
                           n_1985, QN => n31640);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n9141, CK => CLK, Q => 
                           n_1986, QN => n31641);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n9142, CK => CLK, Q => 
                           n_1987, QN => n31642);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n9143, CK => CLK, Q => 
                           n_1988, QN => n31643);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n9144, CK => CLK, Q => 
                           n_1989, QN => n31644);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n9145, CK => CLK, Q => 
                           n_1990, QN => n31645);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n9146, CK => CLK, Q => 
                           n_1991, QN => n31646);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n9147, CK => CLK, Q => 
                           n_1992, QN => n31647);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n9148, CK => CLK, Q => 
                           n_1993, QN => n31648);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n9149, CK => CLK, Q => 
                           n_1994, QN => n31649);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n9150, CK => CLK, Q => 
                           n_1995, QN => n31650);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n9151, CK => CLK, Q => 
                           n_1996, QN => n31651);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n9152, CK => CLK, Q => 
                           n_1997, QN => n31652);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n9153, CK => CLK, Q => 
                           n_1998, QN => n31653);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n9154, CK => CLK, Q => 
                           n_1999, QN => n31654);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n9155, CK => CLK, Q => 
                           n_2000, QN => n31655);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n9156, CK => CLK, Q => 
                           n_2001, QN => n31656);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n9157, CK => CLK, Q => 
                           n_2002, QN => n31657);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n9158, CK => CLK, Q => 
                           n_2003, QN => n31658);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n9159, CK => CLK, Q => 
                           n_2004, QN => n31659);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n9160, CK => CLK, Q => 
                           n_2005, QN => n31660);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n9161, CK => CLK, Q => 
                           n_2006, QN => n31661);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n9162, CK => CLK, Q => 
                           n_2007, QN => n31662);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n9163, CK => CLK, Q => 
                           n_2008, QN => n31663);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n9164, CK => CLK, Q => 
                           n_2009, QN => n31664);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n9165, CK => CLK, Q => 
                           n_2010, QN => n31665);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n9166, CK => CLK, Q => 
                           n_2011, QN => n31666);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n9167, CK => CLK, Q => 
                           n_2012, QN => n31667);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n9168, CK => CLK, Q => 
                           n_2013, QN => n31668);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n9169, CK => CLK, Q => 
                           n_2014, QN => n31669);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n9170, CK => CLK, Q => 
                           n_2015, QN => n31670);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n9171, CK => CLK, Q => 
                           n_2016, QN => n31671);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n9172, CK => CLK, Q => 
                           n_2017, QN => n31672);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n9173, CK => CLK, Q => 
                           n_2018, QN => n31673);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n9174, CK => CLK, Q => 
                           n_2019, QN => n31674);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n9175, CK => CLK, Q => 
                           n_2020, QN => n31675);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n9176, CK => CLK, Q => 
                           n_2021, QN => n31676);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n9177, CK => CLK, Q => 
                           n_2022, QN => n31677);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n9178, CK => CLK, Q => 
                           n_2023, QN => n31678);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n9179, CK => CLK, Q => 
                           n_2024, QN => n31679);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n9180, CK => CLK, Q => 
                           n_2025, QN => n31680);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n9181, CK => CLK, Q => 
                           n_2026, QN => n31681);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n9182, CK => CLK, Q => 
                           n_2027, QN => n31682);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n9183, CK => CLK, Q => 
                           n_2028, QN => n31683);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n9184, CK => CLK, Q => 
                           n_2029, QN => n31684);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n9185, CK => CLK, Q => 
                           n_2030, QN => n31685);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n9186, CK => CLK, Q => 
                           n_2031, QN => n31686);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n9187, CK => CLK, Q => 
                           n_2032, QN => n31687);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n9188, CK => CLK, Q => 
                           n_2033, QN => n31688);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n9189, CK => CLK, Q => 
                           n_2034, QN => n31689);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n9190, CK => CLK, Q => 
                           n_2035, QN => n31690);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n9191, CK => CLK, Q => 
                           n_2036, QN => n31691);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n9192, CK => CLK, Q => 
                           n_2037, QN => n31692);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n9193, CK => CLK, Q => 
                           n_2038, QN => n31693);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n9194, CK => CLK, Q => 
                           n_2039, QN => n31694);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n9195, CK => CLK, Q => 
                           n_2040, QN => n31695);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n9196, CK => CLK, Q => 
                           n_2041, QN => n31696);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n9197, CK => CLK, Q => 
                           n_2042, QN => n31697);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n9198, CK => CLK, Q => 
                           n_2043, QN => n31698);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n9199, CK => CLK, Q => 
                           n_2044, QN => n31699);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n9200, CK => CLK, Q => 
                           n_2045, QN => n31700);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n9201, CK => CLK, Q => 
                           n_2046, QN => n31701);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n9202, CK => CLK, Q => 
                           n_2047, QN => n31702);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n9203, CK => CLK, Q => 
                           n_2048, QN => n31703);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n9204, CK => CLK, Q => 
                           n_2049, QN => n31704);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n9205, CK => CLK, Q => 
                           n_2050, QN => n31705);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n9206, CK => CLK, Q => 
                           n_2051, QN => n31706);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n9207, CK => CLK, Q => 
                           n_2052, QN => n31707);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n9208, CK => CLK, Q => 
                           n_2053, QN => n31708);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n9209, CK => CLK, Q => 
                           n_2054, QN => n31709);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n9210, CK => CLK, Q => 
                           n_2055, QN => n31710);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n9211, CK => CLK, Q => 
                           n_2056, QN => n31711);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n9212, CK => CLK, Q => 
                           n_2057, QN => n31712);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n9213, CK => CLK, Q => 
                           n_2058, QN => n31713);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n9214, CK => CLK, Q => 
                           n_2059, QN => n31714);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n9215, CK => CLK, Q => 
                           n_2060, QN => n31715);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n9216, CK => CLK, Q => 
                           n_2061, QN => n31716);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n9217, CK => CLK, Q => 
                           n_2062, QN => n31717);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n9218, CK => CLK, Q => 
                           n_2063, QN => n31718);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n9219, CK => CLK, Q => 
                           n_2064, QN => n31719);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n9220, CK => CLK, Q => 
                           n_2065, QN => n31720);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n9221, CK => CLK, Q => 
                           n_2066, QN => n31721);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n9222, CK => CLK, Q => 
                           n_2067, QN => n31722);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n9223, CK => CLK, Q => 
                           n_2068, QN => n31723);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n9224, CK => CLK, Q => 
                           n_2069, QN => n31724);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n9225, CK => CLK, Q => 
                           n_2070, QN => n31725);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n9226, CK => CLK, Q => 
                           n_2071, QN => n31726);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n9227, CK => CLK, Q => 
                           n_2072, QN => n31727);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n9228, CK => CLK, Q => 
                           n_2073, QN => n31728);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n9229, CK => CLK, Q => 
                           n_2074, QN => n31729);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n9230, CK => CLK, Q => 
                           n_2075, QN => n31730);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n9231, CK => CLK, Q => 
                           n_2076, QN => n31731);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n9232, CK => CLK, Q => 
                           n_2077, QN => n31732);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n9233, CK => CLK, Q => 
                           n_2078, QN => n31733);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n9234, CK => CLK, Q => 
                           n_2079, QN => n31734);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n9235, CK => CLK, Q => 
                           n_2080, QN => n31735);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n9236, CK => CLK, Q => 
                           n_2081, QN => n31736);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n9237, CK => CLK, Q => 
                           n_2082, QN => n31737);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n9238, CK => CLK, Q => 
                           n_2083, QN => n31738);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n9239, CK => CLK, Q => 
                           n_2084, QN => n31739);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n9240, CK => CLK, Q => 
                           n_2085, QN => n31740);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n9241, CK => CLK, Q => 
                           n_2086, QN => n31741);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n9242, CK => CLK, Q => 
                           n_2087, QN => n31742);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n9243, CK => CLK, Q => 
                           n_2088, QN => n31743);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n9244, CK => CLK, Q => 
                           n_2089, QN => n31744);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n9245, CK => CLK, Q => 
                           n_2090, QN => n31745);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n9246, CK => CLK, Q => 
                           n_2091, QN => n31746);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n9247, CK => CLK, Q => 
                           n_2092, QN => n31747);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n9248, CK => CLK, Q => 
                           n_2093, QN => n31748);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n9249, CK => CLK, Q => 
                           n_2094, QN => n31749);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n9250, CK => CLK, Q => 
                           n_2095, QN => n31750);
   REGISTERS_reg_32_63_inst : DFF_X1 port map( D => n9379, CK => CLK, Q => 
                           n_2096, QN => n31751);
   REGISTERS_reg_32_62_inst : DFF_X1 port map( D => n9380, CK => CLK, Q => 
                           n_2097, QN => n31752);
   REGISTERS_reg_32_61_inst : DFF_X1 port map( D => n9381, CK => CLK, Q => 
                           n_2098, QN => n31753);
   REGISTERS_reg_32_60_inst : DFF_X1 port map( D => n9382, CK => CLK, Q => 
                           n_2099, QN => n31754);
   REGISTERS_reg_32_59_inst : DFF_X1 port map( D => n9383, CK => CLK, Q => 
                           n_2100, QN => n31755);
   REGISTERS_reg_32_58_inst : DFF_X1 port map( D => n9384, CK => CLK, Q => 
                           n_2101, QN => n31756);
   REGISTERS_reg_32_57_inst : DFF_X1 port map( D => n9385, CK => CLK, Q => 
                           n_2102, QN => n31757);
   REGISTERS_reg_32_56_inst : DFF_X1 port map( D => n9386, CK => CLK, Q => 
                           n_2103, QN => n31758);
   REGISTERS_reg_32_55_inst : DFF_X1 port map( D => n9387, CK => CLK, Q => 
                           n_2104, QN => n31759);
   REGISTERS_reg_32_54_inst : DFF_X1 port map( D => n9388, CK => CLK, Q => 
                           n_2105, QN => n31760);
   REGISTERS_reg_32_53_inst : DFF_X1 port map( D => n9389, CK => CLK, Q => 
                           n_2106, QN => n31761);
   REGISTERS_reg_32_52_inst : DFF_X1 port map( D => n9390, CK => CLK, Q => 
                           n_2107, QN => n31762);
   REGISTERS_reg_32_51_inst : DFF_X1 port map( D => n9391, CK => CLK, Q => 
                           n_2108, QN => n31763);
   REGISTERS_reg_32_50_inst : DFF_X1 port map( D => n9392, CK => CLK, Q => 
                           n_2109, QN => n31764);
   REGISTERS_reg_32_49_inst : DFF_X1 port map( D => n9393, CK => CLK, Q => 
                           n_2110, QN => n31765);
   REGISTERS_reg_32_48_inst : DFF_X1 port map( D => n9394, CK => CLK, Q => 
                           n_2111, QN => n31766);
   REGISTERS_reg_32_47_inst : DFF_X1 port map( D => n9395, CK => CLK, Q => 
                           n_2112, QN => n31767);
   REGISTERS_reg_32_46_inst : DFF_X1 port map( D => n9396, CK => CLK, Q => 
                           n_2113, QN => n31768);
   REGISTERS_reg_32_45_inst : DFF_X1 port map( D => n9397, CK => CLK, Q => 
                           n_2114, QN => n31769);
   REGISTERS_reg_32_44_inst : DFF_X1 port map( D => n9398, CK => CLK, Q => 
                           n_2115, QN => n31770);
   REGISTERS_reg_32_43_inst : DFF_X1 port map( D => n9399, CK => CLK, Q => 
                           n_2116, QN => n31771);
   REGISTERS_reg_32_42_inst : DFF_X1 port map( D => n9400, CK => CLK, Q => 
                           n_2117, QN => n31772);
   REGISTERS_reg_32_41_inst : DFF_X1 port map( D => n9401, CK => CLK, Q => 
                           n_2118, QN => n31773);
   REGISTERS_reg_32_40_inst : DFF_X1 port map( D => n9402, CK => CLK, Q => 
                           n_2119, QN => n31774);
   REGISTERS_reg_32_39_inst : DFF_X1 port map( D => n9403, CK => CLK, Q => 
                           n_2120, QN => n31775);
   REGISTERS_reg_32_38_inst : DFF_X1 port map( D => n9404, CK => CLK, Q => 
                           n_2121, QN => n31776);
   REGISTERS_reg_32_37_inst : DFF_X1 port map( D => n9405, CK => CLK, Q => 
                           n_2122, QN => n31777);
   REGISTERS_reg_32_36_inst : DFF_X1 port map( D => n9406, CK => CLK, Q => 
                           n_2123, QN => n31778);
   REGISTERS_reg_32_35_inst : DFF_X1 port map( D => n9407, CK => CLK, Q => 
                           n_2124, QN => n31779);
   REGISTERS_reg_32_34_inst : DFF_X1 port map( D => n9408, CK => CLK, Q => 
                           n_2125, QN => n31780);
   REGISTERS_reg_32_33_inst : DFF_X1 port map( D => n9409, CK => CLK, Q => 
                           n_2126, QN => n31781);
   REGISTERS_reg_32_32_inst : DFF_X1 port map( D => n9410, CK => CLK, Q => 
                           n_2127, QN => n31782);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n9411, CK => CLK, Q => 
                           n_2128, QN => n31783);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n9412, CK => CLK, Q => 
                           n_2129, QN => n31784);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n9413, CK => CLK, Q => 
                           n_2130, QN => n31785);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n9414, CK => CLK, Q => 
                           n_2131, QN => n31786);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n9415, CK => CLK, Q => 
                           n_2132, QN => n31787);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n9416, CK => CLK, Q => 
                           n_2133, QN => n31788);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n9417, CK => CLK, Q => 
                           n_2134, QN => n31789);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n9418, CK => CLK, Q => 
                           n_2135, QN => n31790);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n9419, CK => CLK, Q => 
                           n_2136, QN => n31791);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n9420, CK => CLK, Q => 
                           n_2137, QN => n31792);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n9421, CK => CLK, Q => 
                           n_2138, QN => n31793);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n9422, CK => CLK, Q => 
                           n_2139, QN => n31794);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n9423, CK => CLK, Q => 
                           n_2140, QN => n31795);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n9424, CK => CLK, Q => 
                           n_2141, QN => n31796);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n9425, CK => CLK, Q => 
                           n_2142, QN => n31797);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n9426, CK => CLK, Q => 
                           n_2143, QN => n31798);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n9427, CK => CLK, Q => 
                           n_2144, QN => n31799);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n9428, CK => CLK, Q => 
                           n_2145, QN => n31800);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n9429, CK => CLK, Q => 
                           n_2146, QN => n31801);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n9430, CK => CLK, Q => 
                           n_2147, QN => n31802);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n9431, CK => CLK, Q => 
                           n_2148, QN => n31803);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n9432, CK => CLK, Q => 
                           n_2149, QN => n31804);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n9433, CK => CLK, Q => 
                           n_2150, QN => n31805);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n9434, CK => CLK, Q => 
                           n_2151, QN => n31806);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n9435, CK => CLK, Q => 
                           n_2152, QN => n31807);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n9436, CK => CLK, Q => 
                           n_2153, QN => n31808);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n9437, CK => CLK, Q => 
                           n_2154, QN => n31809);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n9438, CK => CLK, Q => 
                           n_2155, QN => n31810);
   REGISTERS_reg_33_63_inst : DFF_X1 port map( D => n9443, CK => CLK, Q => 
                           n_2156, QN => n31811);
   REGISTERS_reg_33_62_inst : DFF_X1 port map( D => n9444, CK => CLK, Q => 
                           n_2157, QN => n31812);
   REGISTERS_reg_33_61_inst : DFF_X1 port map( D => n9445, CK => CLK, Q => 
                           n_2158, QN => n31813);
   REGISTERS_reg_33_60_inst : DFF_X1 port map( D => n9446, CK => CLK, Q => 
                           n_2159, QN => n31814);
   REGISTERS_reg_33_59_inst : DFF_X1 port map( D => n9447, CK => CLK, Q => 
                           n_2160, QN => n31815);
   REGISTERS_reg_33_58_inst : DFF_X1 port map( D => n9448, CK => CLK, Q => 
                           n_2161, QN => n31816);
   REGISTERS_reg_33_57_inst : DFF_X1 port map( D => n9449, CK => CLK, Q => 
                           n_2162, QN => n31817);
   REGISTERS_reg_33_56_inst : DFF_X1 port map( D => n9450, CK => CLK, Q => 
                           n_2163, QN => n31818);
   REGISTERS_reg_33_55_inst : DFF_X1 port map( D => n9451, CK => CLK, Q => 
                           n_2164, QN => n31819);
   REGISTERS_reg_33_54_inst : DFF_X1 port map( D => n9452, CK => CLK, Q => 
                           n_2165, QN => n31820);
   REGISTERS_reg_33_53_inst : DFF_X1 port map( D => n9453, CK => CLK, Q => 
                           n_2166, QN => n31821);
   REGISTERS_reg_33_52_inst : DFF_X1 port map( D => n9454, CK => CLK, Q => 
                           n_2167, QN => n31822);
   REGISTERS_reg_33_51_inst : DFF_X1 port map( D => n9455, CK => CLK, Q => 
                           n_2168, QN => n31823);
   REGISTERS_reg_33_50_inst : DFF_X1 port map( D => n9456, CK => CLK, Q => 
                           n_2169, QN => n31824);
   REGISTERS_reg_33_49_inst : DFF_X1 port map( D => n9457, CK => CLK, Q => 
                           n_2170, QN => n31825);
   REGISTERS_reg_33_48_inst : DFF_X1 port map( D => n9458, CK => CLK, Q => 
                           n_2171, QN => n31826);
   REGISTERS_reg_33_47_inst : DFF_X1 port map( D => n9459, CK => CLK, Q => 
                           n_2172, QN => n31827);
   REGISTERS_reg_33_46_inst : DFF_X1 port map( D => n9460, CK => CLK, Q => 
                           n_2173, QN => n31828);
   REGISTERS_reg_33_45_inst : DFF_X1 port map( D => n9461, CK => CLK, Q => 
                           n_2174, QN => n31829);
   REGISTERS_reg_33_44_inst : DFF_X1 port map( D => n9462, CK => CLK, Q => 
                           n_2175, QN => n31830);
   REGISTERS_reg_33_43_inst : DFF_X1 port map( D => n9463, CK => CLK, Q => 
                           n_2176, QN => n31831);
   REGISTERS_reg_33_42_inst : DFF_X1 port map( D => n9464, CK => CLK, Q => 
                           n_2177, QN => n31832);
   REGISTERS_reg_33_41_inst : DFF_X1 port map( D => n9465, CK => CLK, Q => 
                           n_2178, QN => n31833);
   REGISTERS_reg_33_40_inst : DFF_X1 port map( D => n9466, CK => CLK, Q => 
                           n_2179, QN => n31834);
   REGISTERS_reg_33_39_inst : DFF_X1 port map( D => n9467, CK => CLK, Q => 
                           n_2180, QN => n31835);
   REGISTERS_reg_33_38_inst : DFF_X1 port map( D => n9468, CK => CLK, Q => 
                           n_2181, QN => n31836);
   REGISTERS_reg_33_37_inst : DFF_X1 port map( D => n9469, CK => CLK, Q => 
                           n_2182, QN => n31837);
   REGISTERS_reg_33_36_inst : DFF_X1 port map( D => n9470, CK => CLK, Q => 
                           n_2183, QN => n31838);
   REGISTERS_reg_33_35_inst : DFF_X1 port map( D => n9471, CK => CLK, Q => 
                           n_2184, QN => n31839);
   REGISTERS_reg_33_34_inst : DFF_X1 port map( D => n9472, CK => CLK, Q => 
                           n_2185, QN => n31840);
   REGISTERS_reg_33_33_inst : DFF_X1 port map( D => n9473, CK => CLK, Q => 
                           n_2186, QN => n31841);
   REGISTERS_reg_33_32_inst : DFF_X1 port map( D => n9474, CK => CLK, Q => 
                           n_2187, QN => n31842);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n9475, CK => CLK, Q => 
                           n_2188, QN => n31843);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n9476, CK => CLK, Q => 
                           n_2189, QN => n31844);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n9477, CK => CLK, Q => 
                           n_2190, QN => n31845);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n9478, CK => CLK, Q => 
                           n_2191, QN => n31846);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n9479, CK => CLK, Q => 
                           n_2192, QN => n31847);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n9480, CK => CLK, Q => 
                           n_2193, QN => n31848);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n9481, CK => CLK, Q => 
                           n_2194, QN => n31849);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n9482, CK => CLK, Q => 
                           n_2195, QN => n31850);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n9483, CK => CLK, Q => 
                           n_2196, QN => n31851);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n9484, CK => CLK, Q => 
                           n_2197, QN => n31852);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n9485, CK => CLK, Q => 
                           n_2198, QN => n31853);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n9486, CK => CLK, Q => 
                           n_2199, QN => n31854);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n9487, CK => CLK, Q => 
                           n_2200, QN => n31855);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n9488, CK => CLK, Q => 
                           n_2201, QN => n31856);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n9489, CK => CLK, Q => 
                           n_2202, QN => n31857);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n9490, CK => CLK, Q => 
                           n_2203, QN => n31858);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n9491, CK => CLK, Q => 
                           n_2204, QN => n31859);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n9492, CK => CLK, Q => 
                           n_2205, QN => n31860);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n9493, CK => CLK, Q => 
                           n_2206, QN => n31861);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n9494, CK => CLK, Q => 
                           n_2207, QN => n31862);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n9495, CK => CLK, Q => 
                           n_2208, QN => n31863);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n9496, CK => CLK, Q => 
                           n_2209, QN => n31864);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n9497, CK => CLK, Q => 
                           n_2210, QN => n31865);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n9498, CK => CLK, Q => 
                           n_2211, QN => n31866);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n9499, CK => CLK, Q => 
                           n_2212, QN => n31867);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n9500, CK => CLK, Q => 
                           n_2213, QN => n31868);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n9501, CK => CLK, Q => 
                           n_2214, QN => n31869);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n9502, CK => CLK, Q => 
                           n_2215, QN => n31870);
   REGISTERS_reg_34_63_inst : DFF_X1 port map( D => n9507, CK => CLK, Q => 
                           n_2216, QN => n31871);
   REGISTERS_reg_34_62_inst : DFF_X1 port map( D => n9508, CK => CLK, Q => 
                           n_2217, QN => n31872);
   REGISTERS_reg_34_61_inst : DFF_X1 port map( D => n9509, CK => CLK, Q => 
                           n_2218, QN => n31873);
   REGISTERS_reg_34_60_inst : DFF_X1 port map( D => n9510, CK => CLK, Q => 
                           n_2219, QN => n31874);
   REGISTERS_reg_34_59_inst : DFF_X1 port map( D => n9511, CK => CLK, Q => 
                           n_2220, QN => n31875);
   REGISTERS_reg_34_58_inst : DFF_X1 port map( D => n9512, CK => CLK, Q => 
                           n_2221, QN => n31876);
   REGISTERS_reg_34_57_inst : DFF_X1 port map( D => n9513, CK => CLK, Q => 
                           n_2222, QN => n31877);
   REGISTERS_reg_34_56_inst : DFF_X1 port map( D => n9514, CK => CLK, Q => 
                           n_2223, QN => n31878);
   REGISTERS_reg_34_55_inst : DFF_X1 port map( D => n9515, CK => CLK, Q => 
                           n_2224, QN => n31879);
   REGISTERS_reg_34_54_inst : DFF_X1 port map( D => n9516, CK => CLK, Q => 
                           n_2225, QN => n31880);
   REGISTERS_reg_34_53_inst : DFF_X1 port map( D => n9517, CK => CLK, Q => 
                           n_2226, QN => n31881);
   REGISTERS_reg_34_52_inst : DFF_X1 port map( D => n9518, CK => CLK, Q => 
                           n_2227, QN => n31882);
   REGISTERS_reg_34_51_inst : DFF_X1 port map( D => n9519, CK => CLK, Q => 
                           n_2228, QN => n31883);
   REGISTERS_reg_34_50_inst : DFF_X1 port map( D => n9520, CK => CLK, Q => 
                           n_2229, QN => n31884);
   REGISTERS_reg_34_49_inst : DFF_X1 port map( D => n9521, CK => CLK, Q => 
                           n_2230, QN => n31885);
   REGISTERS_reg_34_48_inst : DFF_X1 port map( D => n9522, CK => CLK, Q => 
                           n_2231, QN => n31886);
   REGISTERS_reg_34_47_inst : DFF_X1 port map( D => n9523, CK => CLK, Q => 
                           n_2232, QN => n31887);
   REGISTERS_reg_34_46_inst : DFF_X1 port map( D => n9524, CK => CLK, Q => 
                           n_2233, QN => n31888);
   REGISTERS_reg_34_45_inst : DFF_X1 port map( D => n9525, CK => CLK, Q => 
                           n_2234, QN => n31889);
   REGISTERS_reg_34_44_inst : DFF_X1 port map( D => n9526, CK => CLK, Q => 
                           n_2235, QN => n31890);
   REGISTERS_reg_34_43_inst : DFF_X1 port map( D => n9527, CK => CLK, Q => 
                           n_2236, QN => n31891);
   REGISTERS_reg_34_42_inst : DFF_X1 port map( D => n9528, CK => CLK, Q => 
                           n_2237, QN => n31892);
   REGISTERS_reg_34_41_inst : DFF_X1 port map( D => n9529, CK => CLK, Q => 
                           n_2238, QN => n31893);
   REGISTERS_reg_34_40_inst : DFF_X1 port map( D => n9530, CK => CLK, Q => 
                           n_2239, QN => n31894);
   REGISTERS_reg_34_39_inst : DFF_X1 port map( D => n9531, CK => CLK, Q => 
                           n_2240, QN => n31895);
   REGISTERS_reg_34_38_inst : DFF_X1 port map( D => n9532, CK => CLK, Q => 
                           n_2241, QN => n31896);
   REGISTERS_reg_34_37_inst : DFF_X1 port map( D => n9533, CK => CLK, Q => 
                           n_2242, QN => n31897);
   REGISTERS_reg_34_36_inst : DFF_X1 port map( D => n9534, CK => CLK, Q => 
                           n_2243, QN => n31898);
   REGISTERS_reg_34_35_inst : DFF_X1 port map( D => n9535, CK => CLK, Q => 
                           n_2244, QN => n31899);
   REGISTERS_reg_34_34_inst : DFF_X1 port map( D => n9536, CK => CLK, Q => 
                           n_2245, QN => n31900);
   REGISTERS_reg_34_33_inst : DFF_X1 port map( D => n9537, CK => CLK, Q => 
                           n_2246, QN => n31901);
   REGISTERS_reg_34_32_inst : DFF_X1 port map( D => n9538, CK => CLK, Q => 
                           n_2247, QN => n31902);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n9539, CK => CLK, Q => 
                           n_2248, QN => n31903);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n9540, CK => CLK, Q => 
                           n_2249, QN => n31904);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n9541, CK => CLK, Q => 
                           n_2250, QN => n31905);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n9542, CK => CLK, Q => 
                           n_2251, QN => n31906);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n9543, CK => CLK, Q => 
                           n_2252, QN => n31907);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n9544, CK => CLK, Q => 
                           n_2253, QN => n31908);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n9545, CK => CLK, Q => 
                           n_2254, QN => n31909);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n9546, CK => CLK, Q => 
                           n_2255, QN => n31910);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n9547, CK => CLK, Q => 
                           n_2256, QN => n31911);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n9548, CK => CLK, Q => 
                           n_2257, QN => n31912);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n9549, CK => CLK, Q => 
                           n_2258, QN => n31913);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n9550, CK => CLK, Q => 
                           n_2259, QN => n31914);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n9551, CK => CLK, Q => 
                           n_2260, QN => n31915);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n9552, CK => CLK, Q => 
                           n_2261, QN => n31916);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n9553, CK => CLK, Q => 
                           n_2262, QN => n31917);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n9554, CK => CLK, Q => 
                           n_2263, QN => n31918);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n9555, CK => CLK, Q => 
                           n_2264, QN => n31919);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n9556, CK => CLK, Q => 
                           n_2265, QN => n31920);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n9557, CK => CLK, Q => 
                           n_2266, QN => n31921);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n9558, CK => CLK, Q => 
                           n_2267, QN => n31922);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n9559, CK => CLK, Q => 
                           n_2268, QN => n31923);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n9560, CK => CLK, Q => 
                           n_2269, QN => n31924);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n9561, CK => CLK, Q => 
                           n_2270, QN => n31925);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n9562, CK => CLK, Q => 
                           n_2271, QN => n31926);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n9563, CK => CLK, Q => 
                           n_2272, QN => n31927);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n9564, CK => CLK, Q => 
                           n_2273, QN => n31928);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n9565, CK => CLK, Q => 
                           n_2274, QN => n31929);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n9566, CK => CLK, Q => 
                           n_2275, QN => n31930);
   REGISTERS_reg_37_63_inst : DFF_X1 port map( D => n9699, CK => CLK, Q => 
                           n_2276, QN => n31931);
   REGISTERS_reg_37_62_inst : DFF_X1 port map( D => n9700, CK => CLK, Q => 
                           n_2277, QN => n31932);
   REGISTERS_reg_37_61_inst : DFF_X1 port map( D => n9701, CK => CLK, Q => 
                           n_2278, QN => n31933);
   REGISTERS_reg_37_60_inst : DFF_X1 port map( D => n9702, CK => CLK, Q => 
                           n_2279, QN => n31934);
   REGISTERS_reg_37_59_inst : DFF_X1 port map( D => n9703, CK => CLK, Q => 
                           n_2280, QN => n31935);
   REGISTERS_reg_37_58_inst : DFF_X1 port map( D => n9704, CK => CLK, Q => 
                           n_2281, QN => n31936);
   REGISTERS_reg_37_57_inst : DFF_X1 port map( D => n9705, CK => CLK, Q => 
                           n_2282, QN => n31937);
   REGISTERS_reg_37_56_inst : DFF_X1 port map( D => n9706, CK => CLK, Q => 
                           n_2283, QN => n31938);
   REGISTERS_reg_37_55_inst : DFF_X1 port map( D => n9707, CK => CLK, Q => 
                           n_2284, QN => n31939);
   REGISTERS_reg_37_54_inst : DFF_X1 port map( D => n9708, CK => CLK, Q => 
                           n_2285, QN => n31940);
   REGISTERS_reg_37_53_inst : DFF_X1 port map( D => n9709, CK => CLK, Q => 
                           n_2286, QN => n31941);
   REGISTERS_reg_37_52_inst : DFF_X1 port map( D => n9710, CK => CLK, Q => 
                           n_2287, QN => n31942);
   REGISTERS_reg_37_51_inst : DFF_X1 port map( D => n9711, CK => CLK, Q => 
                           n_2288, QN => n31943);
   REGISTERS_reg_37_50_inst : DFF_X1 port map( D => n9712, CK => CLK, Q => 
                           n_2289, QN => n31944);
   REGISTERS_reg_37_49_inst : DFF_X1 port map( D => n9713, CK => CLK, Q => 
                           n_2290, QN => n31945);
   REGISTERS_reg_37_48_inst : DFF_X1 port map( D => n9714, CK => CLK, Q => 
                           n_2291, QN => n31946);
   REGISTERS_reg_37_47_inst : DFF_X1 port map( D => n9715, CK => CLK, Q => 
                           n_2292, QN => n31947);
   REGISTERS_reg_37_46_inst : DFF_X1 port map( D => n9716, CK => CLK, Q => 
                           n_2293, QN => n31948);
   REGISTERS_reg_37_45_inst : DFF_X1 port map( D => n9717, CK => CLK, Q => 
                           n_2294, QN => n31949);
   REGISTERS_reg_37_44_inst : DFF_X1 port map( D => n9718, CK => CLK, Q => 
                           n_2295, QN => n31950);
   REGISTERS_reg_37_43_inst : DFF_X1 port map( D => n9719, CK => CLK, Q => 
                           n_2296, QN => n31951);
   REGISTERS_reg_37_42_inst : DFF_X1 port map( D => n9720, CK => CLK, Q => 
                           n_2297, QN => n31952);
   REGISTERS_reg_37_41_inst : DFF_X1 port map( D => n9721, CK => CLK, Q => 
                           n_2298, QN => n31953);
   REGISTERS_reg_37_40_inst : DFF_X1 port map( D => n9722, CK => CLK, Q => 
                           n_2299, QN => n31954);
   REGISTERS_reg_37_39_inst : DFF_X1 port map( D => n9723, CK => CLK, Q => 
                           n_2300, QN => n31955);
   REGISTERS_reg_37_38_inst : DFF_X1 port map( D => n9724, CK => CLK, Q => 
                           n_2301, QN => n31956);
   REGISTERS_reg_37_37_inst : DFF_X1 port map( D => n9725, CK => CLK, Q => 
                           n_2302, QN => n31957);
   REGISTERS_reg_37_36_inst : DFF_X1 port map( D => n9726, CK => CLK, Q => 
                           n_2303, QN => n31958);
   REGISTERS_reg_37_35_inst : DFF_X1 port map( D => n9727, CK => CLK, Q => 
                           n_2304, QN => n31959);
   REGISTERS_reg_37_34_inst : DFF_X1 port map( D => n9728, CK => CLK, Q => 
                           n_2305, QN => n31960);
   REGISTERS_reg_37_33_inst : DFF_X1 port map( D => n9729, CK => CLK, Q => 
                           n_2306, QN => n31961);
   REGISTERS_reg_37_32_inst : DFF_X1 port map( D => n9730, CK => CLK, Q => 
                           n_2307, QN => n31962);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n9731, CK => CLK, Q => 
                           n_2308, QN => n31963);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n9732, CK => CLK, Q => 
                           n_2309, QN => n31964);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n9733, CK => CLK, Q => 
                           n_2310, QN => n31965);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n9734, CK => CLK, Q => 
                           n_2311, QN => n31966);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n9735, CK => CLK, Q => 
                           n_2312, QN => n31967);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n9736, CK => CLK, Q => 
                           n_2313, QN => n31968);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n9737, CK => CLK, Q => 
                           n_2314, QN => n31969);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n9738, CK => CLK, Q => 
                           n_2315, QN => n31970);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n9739, CK => CLK, Q => 
                           n_2316, QN => n31971);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n9740, CK => CLK, Q => 
                           n_2317, QN => n31972);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n9741, CK => CLK, Q => 
                           n_2318, QN => n31973);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n9742, CK => CLK, Q => 
                           n_2319, QN => n31974);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n9743, CK => CLK, Q => 
                           n_2320, QN => n31975);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n9744, CK => CLK, Q => 
                           n_2321, QN => n31976);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n9745, CK => CLK, Q => 
                           n_2322, QN => n31977);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n9746, CK => CLK, Q => 
                           n_2323, QN => n31978);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n9747, CK => CLK, Q => 
                           n_2324, QN => n31979);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n9748, CK => CLK, Q => 
                           n_2325, QN => n31980);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n9749, CK => CLK, Q => 
                           n_2326, QN => n31981);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n9750, CK => CLK, Q => 
                           n_2327, QN => n31982);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n9751, CK => CLK, Q => 
                           n_2328, QN => n31983);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n9752, CK => CLK, Q => 
                           n_2329, QN => n31984);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n9753, CK => CLK, Q => 
                           n_2330, QN => n31985);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n9754, CK => CLK, Q => 
                           n_2331, QN => n31986);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n9755, CK => CLK, Q => 
                           n_2332, QN => n31987);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n9756, CK => CLK, Q => 
                           n_2333, QN => n31988);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n9757, CK => CLK, Q => 
                           n_2334, QN => n31989);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n9758, CK => CLK, Q => 
                           n_2335, QN => n31990);
   REGISTERS_reg_38_63_inst : DFF_X1 port map( D => n9763, CK => CLK, Q => 
                           n_2336, QN => n31991);
   REGISTERS_reg_38_62_inst : DFF_X1 port map( D => n9764, CK => CLK, Q => 
                           n_2337, QN => n31992);
   REGISTERS_reg_38_61_inst : DFF_X1 port map( D => n9765, CK => CLK, Q => 
                           n_2338, QN => n31993);
   REGISTERS_reg_38_60_inst : DFF_X1 port map( D => n9766, CK => CLK, Q => 
                           n_2339, QN => n31994);
   REGISTERS_reg_38_59_inst : DFF_X1 port map( D => n9767, CK => CLK, Q => 
                           n_2340, QN => n31995);
   REGISTERS_reg_38_58_inst : DFF_X1 port map( D => n9768, CK => CLK, Q => 
                           n_2341, QN => n31996);
   REGISTERS_reg_38_57_inst : DFF_X1 port map( D => n9769, CK => CLK, Q => 
                           n_2342, QN => n31997);
   REGISTERS_reg_38_56_inst : DFF_X1 port map( D => n9770, CK => CLK, Q => 
                           n_2343, QN => n31998);
   REGISTERS_reg_38_55_inst : DFF_X1 port map( D => n9771, CK => CLK, Q => 
                           n_2344, QN => n31999);
   REGISTERS_reg_38_54_inst : DFF_X1 port map( D => n9772, CK => CLK, Q => 
                           n_2345, QN => n32000);
   REGISTERS_reg_38_53_inst : DFF_X1 port map( D => n9773, CK => CLK, Q => 
                           n_2346, QN => n32001);
   REGISTERS_reg_38_52_inst : DFF_X1 port map( D => n9774, CK => CLK, Q => 
                           n_2347, QN => n32002);
   REGISTERS_reg_38_51_inst : DFF_X1 port map( D => n9775, CK => CLK, Q => 
                           n_2348, QN => n32003);
   REGISTERS_reg_38_50_inst : DFF_X1 port map( D => n9776, CK => CLK, Q => 
                           n_2349, QN => n32004);
   REGISTERS_reg_38_49_inst : DFF_X1 port map( D => n9777, CK => CLK, Q => 
                           n_2350, QN => n32005);
   REGISTERS_reg_38_48_inst : DFF_X1 port map( D => n9778, CK => CLK, Q => 
                           n_2351, QN => n32006);
   REGISTERS_reg_38_47_inst : DFF_X1 port map( D => n9779, CK => CLK, Q => 
                           n_2352, QN => n32007);
   REGISTERS_reg_38_46_inst : DFF_X1 port map( D => n9780, CK => CLK, Q => 
                           n_2353, QN => n32008);
   REGISTERS_reg_38_45_inst : DFF_X1 port map( D => n9781, CK => CLK, Q => 
                           n_2354, QN => n32009);
   REGISTERS_reg_38_44_inst : DFF_X1 port map( D => n9782, CK => CLK, Q => 
                           n_2355, QN => n32010);
   REGISTERS_reg_38_43_inst : DFF_X1 port map( D => n9783, CK => CLK, Q => 
                           n_2356, QN => n32011);
   REGISTERS_reg_38_42_inst : DFF_X1 port map( D => n9784, CK => CLK, Q => 
                           n_2357, QN => n32012);
   REGISTERS_reg_38_41_inst : DFF_X1 port map( D => n9785, CK => CLK, Q => 
                           n_2358, QN => n32013);
   REGISTERS_reg_38_40_inst : DFF_X1 port map( D => n9786, CK => CLK, Q => 
                           n_2359, QN => n32014);
   REGISTERS_reg_38_39_inst : DFF_X1 port map( D => n9787, CK => CLK, Q => 
                           n_2360, QN => n32015);
   REGISTERS_reg_38_38_inst : DFF_X1 port map( D => n9788, CK => CLK, Q => 
                           n_2361, QN => n32016);
   REGISTERS_reg_38_37_inst : DFF_X1 port map( D => n9789, CK => CLK, Q => 
                           n_2362, QN => n32017);
   REGISTERS_reg_38_36_inst : DFF_X1 port map( D => n9790, CK => CLK, Q => 
                           n_2363, QN => n32018);
   REGISTERS_reg_38_35_inst : DFF_X1 port map( D => n9791, CK => CLK, Q => 
                           n_2364, QN => n32019);
   REGISTERS_reg_38_34_inst : DFF_X1 port map( D => n9792, CK => CLK, Q => 
                           n_2365, QN => n32020);
   REGISTERS_reg_38_33_inst : DFF_X1 port map( D => n9793, CK => CLK, Q => 
                           n_2366, QN => n32021);
   REGISTERS_reg_38_32_inst : DFF_X1 port map( D => n9794, CK => CLK, Q => 
                           n_2367, QN => n32022);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n9795, CK => CLK, Q => 
                           n_2368, QN => n32023);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n9796, CK => CLK, Q => 
                           n_2369, QN => n32024);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n9797, CK => CLK, Q => 
                           n_2370, QN => n32025);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n9798, CK => CLK, Q => 
                           n_2371, QN => n32026);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n9799, CK => CLK, Q => 
                           n_2372, QN => n32027);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n9800, CK => CLK, Q => 
                           n_2373, QN => n32028);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n9801, CK => CLK, Q => 
                           n_2374, QN => n32029);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n9802, CK => CLK, Q => 
                           n_2375, QN => n32030);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n9803, CK => CLK, Q => 
                           n_2376, QN => n32031);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n9804, CK => CLK, Q => 
                           n_2377, QN => n32032);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n9805, CK => CLK, Q => 
                           n_2378, QN => n32033);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n9806, CK => CLK, Q => 
                           n_2379, QN => n32034);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n9807, CK => CLK, Q => 
                           n_2380, QN => n32035);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n9808, CK => CLK, Q => 
                           n_2381, QN => n32036);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n9809, CK => CLK, Q => 
                           n_2382, QN => n32037);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n9810, CK => CLK, Q => 
                           n_2383, QN => n32038);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n9811, CK => CLK, Q => 
                           n_2384, QN => n32039);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n9812, CK => CLK, Q => 
                           n_2385, QN => n32040);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n9813, CK => CLK, Q => 
                           n_2386, QN => n32041);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n9814, CK => CLK, Q => 
                           n_2387, QN => n32042);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n9815, CK => CLK, Q => 
                           n_2388, QN => n32043);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n9816, CK => CLK, Q => 
                           n_2389, QN => n32044);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n9817, CK => CLK, Q => 
                           n_2390, QN => n32045);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n9818, CK => CLK, Q => 
                           n_2391, QN => n32046);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n9819, CK => CLK, Q => 
                           n_2392, QN => n32047);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n9820, CK => CLK, Q => 
                           n_2393, QN => n32048);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n9821, CK => CLK, Q => 
                           n_2394, QN => n32049);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n9822, CK => CLK, Q => 
                           n_2395, QN => n32050);
   REGISTERS_reg_39_63_inst : DFF_X1 port map( D => n9827, CK => CLK, Q => 
                           n_2396, QN => n32051);
   OUT2_reg_63_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => OUT2(63), QN
                           => n16942);
   OUT1_reg_63_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => OUT1(63), QN
                           => n17006);
   REGISTERS_reg_39_62_inst : DFF_X1 port map( D => n9828, CK => CLK, Q => 
                           n_2397, QN => n32052);
   OUT2_reg_62_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => OUT2(62), QN
                           => n16943);
   OUT1_reg_62_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => OUT1(62), QN
                           => n17007);
   REGISTERS_reg_39_61_inst : DFF_X1 port map( D => n9829, CK => CLK, Q => 
                           n_2398, QN => n32053);
   OUT2_reg_61_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => OUT2(61), QN
                           => n16944);
   OUT1_reg_61_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => OUT1(61), QN
                           => n17008);
   OUT2_reg_60_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => OUT2(60), QN
                           => n16945);
   OUT1_reg_60_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => OUT1(60), QN
                           => n17009);
   REGISTERS_reg_39_59_inst : DFF_X1 port map( D => n9831, CK => CLK, Q => 
                           n_2399, QN => n32054);
   OUT2_reg_59_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => OUT2(59), QN
                           => n16946);
   OUT1_reg_59_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => OUT1(59), QN
                           => n17010);
   OUT2_reg_58_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => OUT2(58), QN
                           => n16947);
   OUT1_reg_58_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => OUT1(58), QN
                           => n17011);
   OUT2_reg_57_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => OUT2(57), QN
                           => n16948);
   OUT1_reg_57_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => OUT1(57), QN
                           => n17012);
   OUT2_reg_56_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => OUT2(56), QN
                           => n16949);
   OUT1_reg_56_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => OUT1(56), QN
                           => n17013);
   OUT2_reg_55_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => OUT2(55), QN
                           => n16950);
   OUT1_reg_55_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => OUT1(55), QN
                           => n17014);
   OUT2_reg_54_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => OUT2(54), QN
                           => n16951);
   OUT1_reg_54_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => OUT1(54), QN
                           => n17015);
   OUT2_reg_53_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => OUT2(53), QN
                           => n16952);
   OUT1_reg_53_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => OUT1(53), QN
                           => n17016);
   OUT2_reg_52_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => OUT2(52), QN
                           => n16953);
   OUT1_reg_52_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => OUT1(52), QN
                           => n17017);
   OUT2_reg_51_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => OUT2(51), QN
                           => n16954);
   OUT1_reg_51_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => OUT1(51), QN
                           => n17018);
   OUT2_reg_50_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => OUT2(50), QN
                           => n16955);
   OUT1_reg_50_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => OUT1(50), QN
                           => n17019);
   OUT2_reg_49_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => OUT2(49), QN
                           => n16956);
   OUT1_reg_49_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => OUT1(49), QN
                           => n17020);
   OUT2_reg_48_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => OUT2(48), QN
                           => n16957);
   OUT1_reg_48_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => OUT1(48), QN
                           => n17021);
   OUT2_reg_47_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => OUT2(47), QN
                           => n16958);
   OUT1_reg_47_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => OUT1(47), QN
                           => n17022);
   OUT2_reg_46_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => OUT2(46), QN
                           => n16959);
   OUT1_reg_46_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => OUT1(46), QN
                           => n17023);
   OUT2_reg_45_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => OUT2(45), QN
                           => n16960);
   OUT1_reg_45_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => OUT1(45), QN
                           => n17024);
   OUT2_reg_44_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => OUT2(44), QN
                           => n16961);
   OUT1_reg_44_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => OUT1(44), QN
                           => n17025);
   OUT2_reg_43_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => OUT2(43), QN
                           => n16962);
   OUT1_reg_43_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => OUT1(43), QN
                           => n17026);
   OUT2_reg_42_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => OUT2(42), QN
                           => n16963);
   OUT1_reg_42_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => OUT1(42), QN
                           => n17027);
   OUT2_reg_41_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => OUT2(41), QN
                           => n16964);
   OUT1_reg_41_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => OUT1(41), QN
                           => n17028);
   OUT2_reg_40_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => OUT2(40), QN
                           => n16965);
   OUT1_reg_40_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => OUT1(40), QN
                           => n17029);
   OUT2_reg_39_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => OUT2(39), QN
                           => n16966);
   OUT1_reg_39_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => OUT1(39), QN
                           => n17030);
   OUT2_reg_38_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => OUT2(38), QN
                           => n16967);
   OUT1_reg_38_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => OUT1(38), QN
                           => n17031);
   OUT2_reg_37_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => OUT2(37), QN
                           => n16968);
   OUT1_reg_37_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => OUT1(37), QN
                           => n17032);
   OUT2_reg_36_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => OUT2(36), QN
                           => n16969);
   OUT1_reg_36_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => OUT1(36), QN
                           => n17033);
   OUT2_reg_35_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => OUT2(35), QN
                           => n16970);
   OUT1_reg_35_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => OUT1(35), QN
                           => n17034);
   OUT2_reg_34_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => OUT2(34), QN
                           => n16971);
   OUT1_reg_34_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => OUT1(34), QN
                           => n17035);
   OUT2_reg_33_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => OUT2(33), QN
                           => n16972);
   OUT1_reg_33_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => OUT1(33), QN
                           => n17036);
   OUT2_reg_32_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => OUT2(32), QN
                           => n16973);
   OUT1_reg_32_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => OUT1(32), QN
                           => n17037);
   OUT2_reg_31_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => OUT2(31), QN
                           => n16974);
   OUT1_reg_31_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => OUT1(31), QN
                           => n17038);
   OUT2_reg_30_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => OUT2(30), QN
                           => n16975);
   OUT1_reg_30_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => OUT1(30), QN
                           => n17039);
   OUT2_reg_29_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => OUT2(29), QN
                           => n16976);
   OUT1_reg_29_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => OUT1(29), QN
                           => n17040);
   OUT2_reg_28_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => OUT2(28), QN
                           => n16977);
   OUT1_reg_28_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => OUT1(28), QN
                           => n17041);
   OUT2_reg_27_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => OUT2(27), QN
                           => n16978);
   OUT1_reg_27_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => OUT1(27), QN
                           => n17042);
   OUT2_reg_26_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => OUT2(26), QN
                           => n16979);
   OUT1_reg_26_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => OUT1(26), QN
                           => n17043);
   OUT2_reg_25_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => OUT2(25), QN
                           => n16980);
   OUT1_reg_25_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => OUT1(25), QN
                           => n17044);
   OUT2_reg_24_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => OUT2(24), QN
                           => n16981);
   OUT1_reg_24_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => OUT1(24), QN
                           => n17045);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n9867, CK => CLK, Q => 
                           n_2400, QN => n32055);
   OUT2_reg_23_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => OUT2(23), QN
                           => n16982);
   OUT1_reg_23_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => OUT1(23), QN
                           => n17046);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n9868, CK => CLK, Q => 
                           n_2401, QN => n32056);
   OUT2_reg_22_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => OUT2(22), QN
                           => n16983);
   OUT1_reg_22_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => OUT1(22), QN
                           => n17047);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n9869, CK => CLK, Q => 
                           n_2402, QN => n32057);
   OUT2_reg_21_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => OUT2(21), QN
                           => n16984);
   OUT1_reg_21_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => OUT1(21), QN
                           => n17048);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n9870, CK => CLK, Q => 
                           n_2403, QN => n32058);
   OUT2_reg_20_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => OUT2(20), QN
                           => n16985);
   OUT1_reg_20_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => OUT1(20), QN
                           => n17049);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n9871, CK => CLK, Q => 
                           n_2404, QN => n32059);
   OUT2_reg_19_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => OUT2(19), QN
                           => n16986);
   OUT1_reg_19_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => OUT1(19), QN
                           => n17050);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n9872, CK => CLK, Q => 
                           n_2405, QN => n32060);
   OUT2_reg_18_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => OUT2(18), QN
                           => n16987);
   OUT1_reg_18_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => OUT1(18), QN
                           => n17051);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n9873, CK => CLK, Q => 
                           n_2406, QN => n32061);
   OUT2_reg_17_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => OUT2(17), QN
                           => n16988);
   OUT1_reg_17_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => OUT1(17), QN
                           => n17052);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n9874, CK => CLK, Q => 
                           n_2407, QN => n32062);
   OUT2_reg_16_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => OUT2(16), QN
                           => n16989);
   OUT1_reg_16_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => OUT1(16), QN
                           => n17053);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n9875, CK => CLK, Q => 
                           n_2408, QN => n32063);
   OUT2_reg_15_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => OUT2(15), QN
                           => n16990);
   OUT1_reg_15_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => OUT1(15), QN
                           => n17054);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n9876, CK => CLK, Q => 
                           n_2409, QN => n32064);
   OUT2_reg_14_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => OUT2(14), QN
                           => n16991);
   OUT1_reg_14_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => OUT1(14), QN
                           => n17055);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n9877, CK => CLK, Q => 
                           n_2410, QN => n32065);
   OUT2_reg_13_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => OUT2(13), QN
                           => n16992);
   OUT1_reg_13_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => OUT1(13), QN
                           => n17056);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n9878, CK => CLK, Q => 
                           n_2411, QN => n32066);
   OUT2_reg_12_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => OUT2(12), QN
                           => n16993);
   OUT1_reg_12_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => OUT1(12), QN
                           => n17057);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n9879, CK => CLK, Q => 
                           n_2412, QN => n32067);
   OUT2_reg_11_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => OUT2(11), QN
                           => n16994);
   OUT1_reg_11_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => OUT1(11), QN
                           => n17058);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n9880, CK => CLK, Q => 
                           n_2413, QN => n32068);
   OUT2_reg_10_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => OUT2(10), QN
                           => n16995);
   OUT1_reg_10_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => OUT1(10), QN
                           => n17059);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n9881, CK => CLK, Q => 
                           n_2414, QN => n32069);
   OUT2_reg_9_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => OUT2(9), QN 
                           => n16996);
   OUT1_reg_9_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => OUT1(9), QN 
                           => n17060);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n9882, CK => CLK, Q => 
                           n_2415, QN => n32070);
   OUT2_reg_8_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => OUT2(8), QN 
                           => n16997);
   OUT1_reg_8_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => OUT1(8), QN 
                           => n17061);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n9883, CK => CLK, Q => 
                           n_2416, QN => n32071);
   OUT2_reg_7_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => OUT2(7), QN 
                           => n16998);
   OUT1_reg_7_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => OUT1(7), QN 
                           => n17062);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n9884, CK => CLK, Q => 
                           n_2417, QN => n32072);
   OUT2_reg_6_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => OUT2(6), QN 
                           => n16999);
   OUT1_reg_6_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => OUT1(6), QN 
                           => n17063);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n9885, CK => CLK, Q => 
                           n_2418, QN => n32073);
   OUT2_reg_5_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => OUT2(5), QN 
                           => n17000);
   OUT1_reg_5_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => OUT1(5), QN 
                           => n17064);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n9886, CK => CLK, Q => 
                           n_2419, QN => n32074);
   OUT2_reg_4_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => OUT2(4), QN 
                           => n17001);
   OUT1_reg_4_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => OUT1(4), QN 
                           => n17065);
   OUT2_reg_3_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => OUT2(3), QN 
                           => n17002);
   OUT1_reg_3_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => OUT1(3), QN 
                           => n17066);
   OUT2_reg_2_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => OUT2(2), QN 
                           => n17003);
   OUT1_reg_2_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => OUT1(2), QN 
                           => n17067);
   OUT2_reg_1_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => OUT2(1), QN 
                           => n17004);
   OUT1_reg_1_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => OUT1(1), QN 
                           => n17068);
   OUT2_reg_0_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => OUT2(0), QN 
                           => n17005);
   OUT1_reg_0_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => OUT1(0), QN 
                           => n17069);
   BUSout_reg_59_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => BUSout(59)
                           , QN => n16937);
   BUSout_reg_58_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => BUSout(58)
                           , QN => n16936);
   BUSout_reg_57_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => BUSout(57)
                           , QN => n16935);
   BUSout_reg_56_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => BUSout(56)
                           , QN => n16934);
   BUSout_reg_55_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => BUSout(55)
                           , QN => n16933);
   BUSout_reg_54_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => BUSout(54)
                           , QN => n16932);
   BUSout_reg_0_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => BUSout(0), 
                           QN => n16878);
   add_146_U1_1 : FA_X1 port map( A => N659, B => i_1_port, CI => n12791, CO =>
                           add_146_carry_2_port, S => N811);
   add_146_U1_2 : FA_X1 port map( A => N660, B => i_2_port, CI => 
                           add_146_carry_2_port, CO => add_146_carry_3_port, S 
                           => N812);
   add_146_U1_3 : FA_X1 port map( A => N661, B => i_3_port, CI => 
                           add_146_carry_3_port, CO => add_146_carry_4_port, S 
                           => N813);
   r510_U1_1 : FA_X1 port map( A => U3_U195_Z_1, B => ADD_RD2(1), CI => r510_n3
                           , CO => r510_carry_2_port, S => N6395);
   r510_U1_2 : FA_X1 port map( A => U3_U195_Z_2, B => ADD_RD2(2), CI => 
                           r510_carry_2_port, CO => r510_carry_3_port, S => 
                           N6396);
   r510_U1_3 : FA_X1 port map( A => U3_U195_Z_3, B => ADD_RD2(3), CI => 
                           r510_carry_3_port, CO => r510_carry_4_port, S => 
                           N6397);
   r510_U1_4 : FA_X1 port map( A => U3_U195_Z_4, B => ADD_RD2(4), CI => 
                           r510_carry_4_port, CO => r510_carry_5_port, S => 
                           N6398);
   r504_U1_1 : FA_X1 port map( A => U3_U194_Z_1, B => ADD_RD1(1), CI => r504_n3
                           , CO => r504_carry_2_port, S => N6270);
   r504_U1_2 : FA_X1 port map( A => U3_U194_Z_2, B => ADD_RD1(2), CI => 
                           r504_carry_2_port, CO => r504_carry_3_port, S => 
                           N6271);
   r504_U1_3 : FA_X1 port map( A => U3_U194_Z_3, B => ADD_RD1(3), CI => 
                           r504_carry_3_port, CO => r504_carry_4_port, S => 
                           N6272);
   r504_U1_4 : FA_X1 port map( A => U3_U194_Z_4, B => ADD_RD1(4), CI => 
                           r504_carry_4_port, CO => r504_carry_5_port, S => 
                           N6273);
   r498_U1_1 : FA_X1 port map( A => U3_U193_Z_1, B => ADD_WR(1), CI => r498_n1,
                           CO => r498_carry_2_port, S => N929);
   r498_U1_2 : FA_X1 port map( A => U3_U193_Z_2, B => ADD_WR(2), CI => 
                           r498_carry_2_port, CO => r498_carry_3_port, S => 
                           N930);
   r498_U1_3 : FA_X1 port map( A => U3_U193_Z_3, B => ADD_WR(3), CI => 
                           r498_carry_3_port, CO => r498_carry_4_port, S => 
                           N931);
   r498_U1_4 : FA_X1 port map( A => U3_U193_Z_4, B => ADD_WR(4), CI => 
                           r498_carry_4_port, CO => r498_carry_5_port, S => 
                           N932);
   add_136_U1_1 : FA_X1 port map( A => N659, B => i_1_port, CI => n12791, CO =>
                           add_136_carry_2_port, S => N688);
   add_136_U1_2 : FA_X1 port map( A => N660, B => i_2_port, CI => 
                           add_136_carry_2_port, CO => add_136_carry_3_port, S 
                           => N689);
   add_136_U1_3 : FA_X1 port map( A => N661, B => i_3_port, CI => 
                           add_136_carry_3_port, CO => add_136_carry_4_port, S 
                           => N690);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n9887, CK => CLK, Q => 
                           n_2420, QN => n32262);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n9888, CK => CLK, Q => 
                           n_2421, QN => n32263);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n9889, CK => CLK, Q => 
                           n_2422, QN => n32264);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n9890, CK => CLK, Q => 
                           n_2423, QN => n32265);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n9503, CK => CLK, Q => 
                           n_2424, QN => n32266);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n9504, CK => CLK, Q => 
                           n_2425, QN => n32267);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n9505, CK => CLK, Q => 
                           n_2426, QN => n32268);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n9506, CK => CLK, Q => 
                           n_2427, QN => n32269);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n9567, CK => CLK, Q => 
                           n_2428, QN => n32270);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n9568, CK => CLK, Q => 
                           n_2429, QN => n32271);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n9569, CK => CLK, Q => 
                           n_2430, QN => n32272);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n9570, CK => CLK, Q => 
                           n_2431, QN => n32273);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n9439, CK => CLK, Q => 
                           n_2432, QN => n32274);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n9440, CK => CLK, Q => 
                           n_2433, QN => n32275);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n9441, CK => CLK, Q => 
                           n_2434, QN => n32276);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n9442, CK => CLK, Q => 
                           n_2435, QN => n32277);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n9823, CK => CLK, Q => 
                           n_2436, QN => n32278);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n9824, CK => CLK, Q => 
                           n_2437, QN => n32279);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n9825, CK => CLK, Q => 
                           n_2438, QN => n32280);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n9826, CK => CLK, Q => 
                           n_2439, QN => n32281);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n9759, CK => CLK, Q => 
                           n_2440, QN => n32282);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n9760, CK => CLK, Q => 
                           n_2441, QN => n32283);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n9761, CK => CLK, Q => 
                           n_2442, QN => n32284);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n9762, CK => CLK, Q => 
                           n_2443, QN => n32285);
   REGISTERS_reg_39_60_inst : DFF_X1 port map( D => n9830, CK => CLK, Q => 
                           n_2444, QN => n32286);
   REGISTERS_reg_39_58_inst : DFF_X1 port map( D => n9832, CK => CLK, Q => 
                           n_2445, QN => n32287);
   REGISTERS_reg_39_57_inst : DFF_X1 port map( D => n9833, CK => CLK, Q => 
                           n_2446, QN => n32288);
   REGISTERS_reg_39_56_inst : DFF_X1 port map( D => n9834, CK => CLK, Q => 
                           n_2447, QN => n32289);
   REGISTERS_reg_39_55_inst : DFF_X1 port map( D => n9835, CK => CLK, Q => 
                           n_2448, QN => n32290);
   REGISTERS_reg_39_54_inst : DFF_X1 port map( D => n9836, CK => CLK, Q => 
                           n_2449, QN => n32291);
   REGISTERS_reg_39_53_inst : DFF_X1 port map( D => n9837, CK => CLK, Q => 
                           n_2450, QN => n32292);
   REGISTERS_reg_39_52_inst : DFF_X1 port map( D => n9838, CK => CLK, Q => 
                           n_2451, QN => n32293);
   REGISTERS_reg_39_51_inst : DFF_X1 port map( D => n9839, CK => CLK, Q => 
                           n_2452, QN => n32294);
   REGISTERS_reg_39_50_inst : DFF_X1 port map( D => n9840, CK => CLK, Q => 
                           n_2453, QN => n32295);
   REGISTERS_reg_39_49_inst : DFF_X1 port map( D => n9841, CK => CLK, Q => 
                           n_2454, QN => n32296);
   REGISTERS_reg_39_48_inst : DFF_X1 port map( D => n9842, CK => CLK, Q => 
                           n_2455, QN => n32297);
   REGISTERS_reg_39_47_inst : DFF_X1 port map( D => n9843, CK => CLK, Q => 
                           n_2456, QN => n32298);
   REGISTERS_reg_39_46_inst : DFF_X1 port map( D => n9844, CK => CLK, Q => 
                           n_2457, QN => n32299);
   REGISTERS_reg_39_45_inst : DFF_X1 port map( D => n9845, CK => CLK, Q => 
                           n_2458, QN => n32300);
   REGISTERS_reg_39_44_inst : DFF_X1 port map( D => n9846, CK => CLK, Q => 
                           n_2459, QN => n32301);
   REGISTERS_reg_39_43_inst : DFF_X1 port map( D => n9847, CK => CLK, Q => 
                           n_2460, QN => n32302);
   REGISTERS_reg_39_42_inst : DFF_X1 port map( D => n9848, CK => CLK, Q => 
                           n_2461, QN => n32303);
   REGISTERS_reg_39_41_inst : DFF_X1 port map( D => n9849, CK => CLK, Q => 
                           n_2462, QN => n32304);
   REGISTERS_reg_39_40_inst : DFF_X1 port map( D => n9850, CK => CLK, Q => 
                           n_2463, QN => n32305);
   REGISTERS_reg_39_39_inst : DFF_X1 port map( D => n9851, CK => CLK, Q => 
                           n_2464, QN => n32306);
   REGISTERS_reg_39_38_inst : DFF_X1 port map( D => n9852, CK => CLK, Q => 
                           n_2465, QN => n32307);
   REGISTERS_reg_39_37_inst : DFF_X1 port map( D => n9853, CK => CLK, Q => 
                           n_2466, QN => n32308);
   REGISTERS_reg_39_36_inst : DFF_X1 port map( D => n9854, CK => CLK, Q => 
                           n_2467, QN => n32309);
   REGISTERS_reg_39_35_inst : DFF_X1 port map( D => n9855, CK => CLK, Q => 
                           n_2468, QN => n32310);
   REGISTERS_reg_39_34_inst : DFF_X1 port map( D => n9856, CK => CLK, Q => 
                           n_2469, QN => n32311);
   REGISTERS_reg_39_33_inst : DFF_X1 port map( D => n9857, CK => CLK, Q => 
                           n_2470, QN => n32312);
   REGISTERS_reg_39_32_inst : DFF_X1 port map( D => n9858, CK => CLK, Q => 
                           n_2471, QN => n32313);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n9859, CK => CLK, Q => 
                           n_2472, QN => n32314);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n9860, CK => CLK, Q => 
                           n_2473, QN => n32315);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n9861, CK => CLK, Q => 
                           n_2474, QN => n32316);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n9862, CK => CLK, Q => 
                           n_2475, QN => n32317);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n9863, CK => CLK, Q => 
                           n_2476, QN => n32318);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n9864, CK => CLK, Q => 
                           n_2477, QN => n32319);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n9865, CK => CLK, Q => 
                           n_2478, QN => n32320);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n9866, CK => CLK, Q => 
                           n_2479, QN => n32321);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n9631, CK => CLK, Q => 
                           n30063, QN => n39046);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n9632, CK => CLK, Q => 
                           n30064, QN => n39045);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n9633, CK => CLK, Q => 
                           n30065, QN => n39044);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n9634, CK => CLK, Q => 
                           n30066, QN => n39043);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n9695, CK => CLK, Q => 
                           n30127, QN => n38923);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n9696, CK => CLK, Q => 
                           n30128, QN => n38922);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n9697, CK => CLK, Q => 
                           n30129, QN => n38921);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n9698, CK => CLK, Q => 
                           n30130, QN => n38920);
   REGISTERS_reg_35_51_inst : DFF_X1 port map( D => n9583, CK => CLK, Q => 
                           n30015, QN => n39042);
   REGISTERS_reg_35_50_inst : DFF_X1 port map( D => n9584, CK => CLK, Q => 
                           n30016, QN => n39041);
   REGISTERS_reg_35_49_inst : DFF_X1 port map( D => n9585, CK => CLK, Q => 
                           n30017, QN => n39040);
   REGISTERS_reg_35_48_inst : DFF_X1 port map( D => n9586, CK => CLK, Q => 
                           n30018, QN => n39039);
   REGISTERS_reg_35_47_inst : DFF_X1 port map( D => n9587, CK => CLK, Q => 
                           n30019, QN => n39038);
   REGISTERS_reg_35_46_inst : DFF_X1 port map( D => n9588, CK => CLK, Q => 
                           n30020, QN => n39037);
   REGISTERS_reg_35_45_inst : DFF_X1 port map( D => n9589, CK => CLK, Q => 
                           n30021, QN => n39036);
   REGISTERS_reg_35_44_inst : DFF_X1 port map( D => n9590, CK => CLK, Q => 
                           n30022, QN => n39035);
   REGISTERS_reg_35_43_inst : DFF_X1 port map( D => n9591, CK => CLK, Q => 
                           n30023, QN => n39034);
   REGISTERS_reg_35_42_inst : DFF_X1 port map( D => n9592, CK => CLK, Q => 
                           n30024, QN => n39033);
   REGISTERS_reg_35_41_inst : DFF_X1 port map( D => n9593, CK => CLK, Q => 
                           n30025, QN => n39032);
   REGISTERS_reg_35_40_inst : DFF_X1 port map( D => n9594, CK => CLK, Q => 
                           n30026, QN => n39031);
   REGISTERS_reg_35_39_inst : DFF_X1 port map( D => n9595, CK => CLK, Q => 
                           n30027, QN => n39030);
   REGISTERS_reg_35_38_inst : DFF_X1 port map( D => n9596, CK => CLK, Q => 
                           n30028, QN => n39029);
   REGISTERS_reg_35_37_inst : DFF_X1 port map( D => n9597, CK => CLK, Q => 
                           n30029, QN => n39028);
   REGISTERS_reg_35_36_inst : DFF_X1 port map( D => n9598, CK => CLK, Q => 
                           n30030, QN => n39027);
   REGISTERS_reg_35_35_inst : DFF_X1 port map( D => n9599, CK => CLK, Q => 
                           n30031, QN => n39026);
   REGISTERS_reg_35_34_inst : DFF_X1 port map( D => n9600, CK => CLK, Q => 
                           n30032, QN => n39025);
   REGISTERS_reg_35_33_inst : DFF_X1 port map( D => n9601, CK => CLK, Q => 
                           n30033, QN => n39024);
   REGISTERS_reg_35_32_inst : DFF_X1 port map( D => n9602, CK => CLK, Q => 
                           n30034, QN => n39023);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n9603, CK => CLK, Q => 
                           n30035, QN => n39022);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n9604, CK => CLK, Q => 
                           n30036, QN => n39021);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n9605, CK => CLK, Q => 
                           n30037, QN => n39020);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n9606, CK => CLK, Q => 
                           n30038, QN => n39019);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n9607, CK => CLK, Q => 
                           n30039, QN => n39018);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n9608, CK => CLK, Q => 
                           n30040, QN => n39017);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n9609, CK => CLK, Q => 
                           n30041, QN => n39016);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n9610, CK => CLK, Q => 
                           n30042, QN => n39015);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n9611, CK => CLK, Q => 
                           n30043, QN => n39014);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n9612, CK => CLK, Q => 
                           n30044, QN => n39013);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n9613, CK => CLK, Q => 
                           n30045, QN => n39012);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n9614, CK => CLK, Q => 
                           n30046, QN => n39011);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n9615, CK => CLK, Q => 
                           n30047, QN => n39010);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n9616, CK => CLK, Q => 
                           n30048, QN => n39009);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n9617, CK => CLK, Q => 
                           n30049, QN => n39008);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n9618, CK => CLK, Q => 
                           n30050, QN => n39007);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n9619, CK => CLK, Q => 
                           n30051, QN => n39006);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n9620, CK => CLK, Q => 
                           n30052, QN => n39005);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n9621, CK => CLK, Q => 
                           n30053, QN => n39004);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n9622, CK => CLK, Q => 
                           n30054, QN => n39003);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n9623, CK => CLK, Q => 
                           n30055, QN => n39002);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n9624, CK => CLK, Q => 
                           n30056, QN => n39001);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n9625, CK => CLK, Q => 
                           n30057, QN => n39000);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n9626, CK => CLK, Q => 
                           n30058, QN => n38999);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n9627, CK => CLK, Q => 
                           n30059, QN => n38998);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n9628, CK => CLK, Q => 
                           n30060, QN => n38997);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n9629, CK => CLK, Q => 
                           n30061, QN => n38996);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n9630, CK => CLK, Q => 
                           n30062, QN => n38995);
   REGISTERS_reg_35_63_inst : DFF_X1 port map( D => n9571, CK => CLK, Q => 
                           n30003, QN => n38926);
   REGISTERS_reg_35_62_inst : DFF_X1 port map( D => n9572, CK => CLK, Q => 
                           n30004, QN => n38925);
   REGISTERS_reg_35_61_inst : DFF_X1 port map( D => n9573, CK => CLK, Q => 
                           n30005, QN => n38924);
   REGISTERS_reg_35_60_inst : DFF_X1 port map( D => n9574, CK => CLK, Q => 
                           n30006, QN => n38994);
   REGISTERS_reg_35_59_inst : DFF_X1 port map( D => n9575, CK => CLK, Q => 
                           n30007, QN => n32384);
   REGISTERS_reg_35_58_inst : DFF_X1 port map( D => n9576, CK => CLK, Q => 
                           n30008, QN => n38993);
   REGISTERS_reg_35_57_inst : DFF_X1 port map( D => n9577, CK => CLK, Q => 
                           n30009, QN => n38992);
   REGISTERS_reg_35_56_inst : DFF_X1 port map( D => n9578, CK => CLK, Q => 
                           n30010, QN => n38991);
   REGISTERS_reg_35_55_inst : DFF_X1 port map( D => n9579, CK => CLK, Q => 
                           n30011, QN => n38990);
   REGISTERS_reg_35_54_inst : DFF_X1 port map( D => n9580, CK => CLK, Q => 
                           n30012, QN => n38989);
   REGISTERS_reg_35_53_inst : DFF_X1 port map( D => n9581, CK => CLK, Q => 
                           n30013, QN => n38988);
   REGISTERS_reg_35_52_inst : DFF_X1 port map( D => n9582, CK => CLK, Q => 
                           n30014, QN => n38987);
   REGISTERS_reg_36_51_inst : DFF_X1 port map( D => n9647, CK => CLK, Q => 
                           n30079, QN => n38919);
   REGISTERS_reg_36_50_inst : DFF_X1 port map( D => n9648, CK => CLK, Q => 
                           n30080, QN => n38918);
   REGISTERS_reg_36_49_inst : DFF_X1 port map( D => n9649, CK => CLK, Q => 
                           n30081, QN => n38917);
   REGISTERS_reg_36_48_inst : DFF_X1 port map( D => n9650, CK => CLK, Q => 
                           n30082, QN => n38916);
   REGISTERS_reg_36_47_inst : DFF_X1 port map( D => n9651, CK => CLK, Q => 
                           n30083, QN => n38915);
   REGISTERS_reg_36_46_inst : DFF_X1 port map( D => n9652, CK => CLK, Q => 
                           n30084, QN => n38914);
   REGISTERS_reg_36_45_inst : DFF_X1 port map( D => n9653, CK => CLK, Q => 
                           n30085, QN => n38913);
   REGISTERS_reg_36_44_inst : DFF_X1 port map( D => n9654, CK => CLK, Q => 
                           n30086, QN => n38912);
   REGISTERS_reg_36_43_inst : DFF_X1 port map( D => n9655, CK => CLK, Q => 
                           n30087, QN => n38911);
   REGISTERS_reg_36_42_inst : DFF_X1 port map( D => n9656, CK => CLK, Q => 
                           n30088, QN => n38910);
   REGISTERS_reg_36_41_inst : DFF_X1 port map( D => n9657, CK => CLK, Q => 
                           n30089, QN => n38909);
   REGISTERS_reg_36_40_inst : DFF_X1 port map( D => n9658, CK => CLK, Q => 
                           n30090, QN => n38908);
   REGISTERS_reg_36_39_inst : DFF_X1 port map( D => n9659, CK => CLK, Q => 
                           n30091, QN => n38907);
   REGISTERS_reg_36_38_inst : DFF_X1 port map( D => n9660, CK => CLK, Q => 
                           n30092, QN => n38906);
   REGISTERS_reg_36_37_inst : DFF_X1 port map( D => n9661, CK => CLK, Q => 
                           n30093, QN => n38905);
   REGISTERS_reg_36_36_inst : DFF_X1 port map( D => n9662, CK => CLK, Q => 
                           n30094, QN => n38904);
   REGISTERS_reg_36_35_inst : DFF_X1 port map( D => n9663, CK => CLK, Q => 
                           n30095, QN => n38903);
   REGISTERS_reg_36_34_inst : DFF_X1 port map( D => n9664, CK => CLK, Q => 
                           n30096, QN => n38902);
   REGISTERS_reg_36_33_inst : DFF_X1 port map( D => n9665, CK => CLK, Q => 
                           n30097, QN => n38901);
   REGISTERS_reg_36_32_inst : DFF_X1 port map( D => n9666, CK => CLK, Q => 
                           n30098, QN => n38900);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n9667, CK => CLK, Q => 
                           n30099, QN => n38899);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n9668, CK => CLK, Q => 
                           n30100, QN => n38898);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n9669, CK => CLK, Q => 
                           n30101, QN => n38897);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n9670, CK => CLK, Q => 
                           n30102, QN => n38896);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n9671, CK => CLK, Q => 
                           n30103, QN => n38895);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n9672, CK => CLK, Q => 
                           n30104, QN => n38894);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n9673, CK => CLK, Q => 
                           n30105, QN => n38893);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n9674, CK => CLK, Q => 
                           n30106, QN => n38892);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n9675, CK => CLK, Q => 
                           n30107, QN => n38891);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n9676, CK => CLK, Q => 
                           n30108, QN => n38890);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n9677, CK => CLK, Q => 
                           n30109, QN => n38889);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n9678, CK => CLK, Q => 
                           n30110, QN => n38888);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n9679, CK => CLK, Q => 
                           n30111, QN => n38887);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n9680, CK => CLK, Q => 
                           n30112, QN => n38886);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n9681, CK => CLK, Q => 
                           n30113, QN => n38885);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n9682, CK => CLK, Q => 
                           n30114, QN => n38884);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n9683, CK => CLK, Q => 
                           n30115, QN => n38883);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n9684, CK => CLK, Q => 
                           n30116, QN => n38882);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n9685, CK => CLK, Q => 
                           n30117, QN => n38881);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n9686, CK => CLK, Q => 
                           n30118, QN => n38880);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n9687, CK => CLK, Q => 
                           n30119, QN => n38879);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n9688, CK => CLK, Q => 
                           n30120, QN => n38878);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n9689, CK => CLK, Q => 
                           n30121, QN => n38877);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n9690, CK => CLK, Q => 
                           n30122, QN => n38876);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n9691, CK => CLK, Q => 
                           n30123, QN => n38875);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n9692, CK => CLK, Q => 
                           n30124, QN => n38874);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n9693, CK => CLK, Q => 
                           n30125, QN => n38873);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n9694, CK => CLK, Q => 
                           n30126, QN => n38872);
   REGISTERS_reg_36_63_inst : DFF_X1 port map( D => n9635, CK => CLK, Q => 
                           n30067, QN => n38793);
   REGISTERS_reg_36_62_inst : DFF_X1 port map( D => n9636, CK => CLK, Q => 
                           n30068, QN => n38792);
   REGISTERS_reg_36_61_inst : DFF_X1 port map( D => n9637, CK => CLK, Q => 
                           n30069, QN => n38791);
   REGISTERS_reg_36_60_inst : DFF_X1 port map( D => n9638, CK => CLK, Q => 
                           n30070, QN => n38871);
   REGISTERS_reg_36_59_inst : DFF_X1 port map( D => n9639, CK => CLK, Q => 
                           n30071, QN => n32444);
   REGISTERS_reg_36_58_inst : DFF_X1 port map( D => n9640, CK => CLK, Q => 
                           n30072, QN => n38870);
   REGISTERS_reg_36_57_inst : DFF_X1 port map( D => n9641, CK => CLK, Q => 
                           n30073, QN => n38869);
   REGISTERS_reg_36_56_inst : DFF_X1 port map( D => n9642, CK => CLK, Q => 
                           n30074, QN => n38868);
   REGISTERS_reg_36_55_inst : DFF_X1 port map( D => n9643, CK => CLK, Q => 
                           n30075, QN => n38867);
   REGISTERS_reg_36_54_inst : DFF_X1 port map( D => n9644, CK => CLK, Q => 
                           n30076, QN => n38866);
   REGISTERS_reg_36_53_inst : DFF_X1 port map( D => n9645, CK => CLK, Q => 
                           n30077, QN => n38865);
   REGISTERS_reg_36_52_inst : DFF_X1 port map( D => n9646, CK => CLK, Q => 
                           n30078, QN => n38864);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n8415, CK => CLK, Q => 
                           n28847, QN => n38863);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n8416, CK => CLK, Q => 
                           n28848, QN => n38862);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n8417, CK => CLK, Q => 
                           n28849, QN => n38861);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n8418, CK => CLK, Q => 
                           n28850, QN => n38860);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n9055, CK => CLK, Q => 
                           n29487, QN => n32460);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n9056, CK => CLK, Q => 
                           n29488, QN => n32461);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n9057, CK => CLK, Q => 
                           n29489, QN => n32462);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n9058, CK => CLK, Q => 
                           n29490, QN => n32463);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n8991, CK => CLK, Q => 
                           n29423, QN => n32464);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n8992, CK => CLK, Q => 
                           n29424, QN => n32465);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n8993, CK => CLK, Q => 
                           n29425, QN => n32466);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n8994, CK => CLK, Q => 
                           n29426, QN => n32467);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n8735, CK => CLK, Q => 
                           n29167, QN => n32476);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n8736, CK => CLK, Q => 
                           n29168, QN => n32477);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n8737, CK => CLK, Q => 
                           n29169, QN => n32478);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n8738, CK => CLK, Q => 
                           n29170, QN => n32479);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n8671, CK => CLK, Q => 
                           n29103, QN => n32480);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n8672, CK => CLK, Q => 
                           n29104, QN => n32481);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n8673, CK => CLK, Q => 
                           n29105, QN => n32482);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n8674, CK => CLK, Q => 
                           n29106, QN => n32483);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n9311, CK => CLK, Q => 
                           n29743, QN => n38986);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n9312, CK => CLK, Q => 
                           n29744, QN => n38985);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n9313, CK => CLK, Q => 
                           n29745, QN => n38984);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n9314, CK => CLK, Q => 
                           n29746, QN => n38983);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n9375, CK => CLK, Q => 
                           n29807, QN => n38859);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n9376, CK => CLK, Q => 
                           n29808, QN => n38858);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n9377, CK => CLK, Q => 
                           n29809, QN => n38857);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n9378, CK => CLK, Q => 
                           n29810, QN => n38856);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n8409, CK => CLK, Q => 
                           n28841, QN => n38855);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n8410, CK => CLK, Q => 
                           n28842, QN => n38854);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n8411, CK => CLK, Q => 
                           n28843, QN => n38853);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n8413, CK => CLK, Q => 
                           n28845, QN => n38852);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n8414, CK => CLK, Q => 
                           n28846, QN => n38851);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n8412, CK => CLK, Q => 
                           n28844, QN => n38850);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n27956, QN => n32547);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n27957, QN => n32548);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n27958, QN => n32549);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n27959, QN => n32550);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n27960, QN => n32551);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n27961, QN => n32552);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n27962, QN => n32553);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n27963, QN => n32554);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n27964, QN => n32555);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n27965, QN => n32556);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n27966, QN => n32557);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n27967, QN => n32558);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n27968, QN => n32559);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n27969, QN => n32560);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n27970, QN => n32561);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n27971, QN => n32562);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => 
                           n27972, QN => n32563);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => 
                           n27973, QN => n32564);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => 
                           n27974, QN => n32565);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => 
                           n27975, QN => n32566);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => 
                           n27976, QN => n32567);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => 
                           n27977, QN => n32568);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => 
                           n27978, QN => n32569);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => 
                           n27979, QN => n32570);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => 
                           n27980, QN => n32571);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => 
                           n27981, QN => n32572);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => 
                           n27982, QN => n32573);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => 
                           n27983, QN => n32574);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => 
                           n27984, QN => n32575);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n27985, QN => n32576);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n27986, QN => n32577);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n27987, QN => n32578);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n27988, QN => n32579);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n27989, QN => n32580);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n27990, QN => n32581);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n27991, QN => n32582);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n27992, QN => n32583);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n27993, QN => n32584);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n27994, QN => n32585);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n27995, QN => n32586);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n27996, QN => n32587);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n27997, QN => n32588);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => n27998
                           , QN => n32589);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => n27999
                           , QN => n32590);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => n28000
                           , QN => n32591);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => n28001
                           , QN => n32592);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => n28002
                           , QN => n32593);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => n28003
                           , QN => n32594);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n9007, CK => CLK, Q => 
                           n29439, QN => n32595);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n9008, CK => CLK, Q => 
                           n29440, QN => n32596);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n9009, CK => CLK, Q => 
                           n29441, QN => n32597);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n9010, CK => CLK, Q => 
                           n29442, QN => n32598);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n9011, CK => CLK, Q => 
                           n29443, QN => n32599);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n9012, CK => CLK, Q => 
                           n29444, QN => n32600);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n9013, CK => CLK, Q => 
                           n29445, QN => n32601);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n9014, CK => CLK, Q => 
                           n29446, QN => n32602);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n9015, CK => CLK, Q => 
                           n29447, QN => n32603);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n9016, CK => CLK, Q => 
                           n29448, QN => n32604);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n9017, CK => CLK, Q => 
                           n29449, QN => n32605);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n9018, CK => CLK, Q => 
                           n29450, QN => n32606);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n9019, CK => CLK, Q => 
                           n29451, QN => n32607);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n9020, CK => CLK, Q => 
                           n29452, QN => n32608);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n9021, CK => CLK, Q => 
                           n29453, QN => n32609);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n9022, CK => CLK, Q => 
                           n29454, QN => n32610);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n9023, CK => CLK, Q => 
                           n29455, QN => n32611);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n9024, CK => CLK, Q => 
                           n29456, QN => n32612);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n9025, CK => CLK, Q => 
                           n29457, QN => n32613);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n9026, CK => CLK, Q => 
                           n29458, QN => n32614);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n9027, CK => CLK, Q => 
                           n29459, QN => n32615);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n9028, CK => CLK, Q => 
                           n29460, QN => n32616);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n9029, CK => CLK, Q => 
                           n29461, QN => n32617);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n9030, CK => CLK, Q => 
                           n29462, QN => n32618);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n9031, CK => CLK, Q => 
                           n29463, QN => n32619);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n9032, CK => CLK, Q => 
                           n29464, QN => n32620);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n9033, CK => CLK, Q => 
                           n29465, QN => n32621);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n9034, CK => CLK, Q => 
                           n29466, QN => n32622);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n9035, CK => CLK, Q => 
                           n29467, QN => n32623);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n9036, CK => CLK, Q => 
                           n29468, QN => n32624);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n9037, CK => CLK, Q => 
                           n29469, QN => n32625);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n9038, CK => CLK, Q => 
                           n29470, QN => n32626);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n9039, CK => CLK, Q => 
                           n29471, QN => n32627);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n9040, CK => CLK, Q => 
                           n29472, QN => n32628);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n9041, CK => CLK, Q => 
                           n29473, QN => n32629);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n9042, CK => CLK, Q => 
                           n29474, QN => n32630);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n9043, CK => CLK, Q => 
                           n29475, QN => n32631);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n9044, CK => CLK, Q => 
                           n29476, QN => n32632);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n9045, CK => CLK, Q => 
                           n29477, QN => n32633);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n9046, CK => CLK, Q => 
                           n29478, QN => n32634);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n9047, CK => CLK, Q => 
                           n29479, QN => n32635);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n9048, CK => CLK, Q => 
                           n29480, QN => n32636);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n9049, CK => CLK, Q => 
                           n29481, QN => n32637);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n9050, CK => CLK, Q => 
                           n29482, QN => n32638);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n9051, CK => CLK, Q => 
                           n29483, QN => n32639);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n9052, CK => CLK, Q => 
                           n29484, QN => n32640);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n9053, CK => CLK, Q => 
                           n29485, QN => n32641);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n9054, CK => CLK, Q => 
                           n29486, QN => n32642);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n8943, CK => CLK, Q => 
                           n29375, QN => n32643);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n8944, CK => CLK, Q => 
                           n29376, QN => n32644);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n8945, CK => CLK, Q => 
                           n29377, QN => n32645);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n8946, CK => CLK, Q => 
                           n29378, QN => n32646);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n8947, CK => CLK, Q => 
                           n29379, QN => n32647);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n8948, CK => CLK, Q => 
                           n29380, QN => n32648);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n8949, CK => CLK, Q => 
                           n29381, QN => n32649);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n8950, CK => CLK, Q => 
                           n29382, QN => n32650);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n8951, CK => CLK, Q => 
                           n29383, QN => n32651);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n8952, CK => CLK, Q => 
                           n29384, QN => n32652);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n8953, CK => CLK, Q => 
                           n29385, QN => n32653);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n8954, CK => CLK, Q => 
                           n29386, QN => n32654);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n8955, CK => CLK, Q => 
                           n29387, QN => n32655);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n8956, CK => CLK, Q => 
                           n29388, QN => n32656);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n8957, CK => CLK, Q => 
                           n29389, QN => n32657);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n8958, CK => CLK, Q => 
                           n29390, QN => n32658);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n8959, CK => CLK, Q => 
                           n29391, QN => n32659);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n8960, CK => CLK, Q => 
                           n29392, QN => n32660);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n8961, CK => CLK, Q => 
                           n29393, QN => n32661);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n8962, CK => CLK, Q => 
                           n29394, QN => n32662);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n8963, CK => CLK, Q => 
                           n29395, QN => n32663);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n8964, CK => CLK, Q => 
                           n29396, QN => n32664);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n8965, CK => CLK, Q => 
                           n29397, QN => n32665);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n8966, CK => CLK, Q => 
                           n29398, QN => n32666);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n8967, CK => CLK, Q => 
                           n29399, QN => n32667);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n8968, CK => CLK, Q => 
                           n29400, QN => n32668);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n8969, CK => CLK, Q => 
                           n29401, QN => n32669);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n8970, CK => CLK, Q => 
                           n29402, QN => n32670);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n8971, CK => CLK, Q => 
                           n29403, QN => n32671);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n8972, CK => CLK, Q => 
                           n29404, QN => n32672);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n8973, CK => CLK, Q => 
                           n29405, QN => n32673);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n8974, CK => CLK, Q => 
                           n29406, QN => n32674);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n8975, CK => CLK, Q => 
                           n29407, QN => n32675);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n8976, CK => CLK, Q => 
                           n29408, QN => n32676);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n8977, CK => CLK, Q => 
                           n29409, QN => n32677);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n8978, CK => CLK, Q => 
                           n29410, QN => n32678);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n8979, CK => CLK, Q => 
                           n29411, QN => n32679);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n8980, CK => CLK, Q => 
                           n29412, QN => n32680);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n8981, CK => CLK, Q => 
                           n29413, QN => n32681);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n8982, CK => CLK, Q => 
                           n29414, QN => n32682);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n8983, CK => CLK, Q => 
                           n29415, QN => n32683);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n8984, CK => CLK, Q => 
                           n29416, QN => n32684);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n8985, CK => CLK, Q => 
                           n29417, QN => n32685);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n8986, CK => CLK, Q => 
                           n29418, QN => n32686);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n8987, CK => CLK, Q => 
                           n29419, QN => n32687);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n8988, CK => CLK, Q => 
                           n29420, QN => n32688);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n8989, CK => CLK, Q => 
                           n29421, QN => n32689);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n8990, CK => CLK, Q => 
                           n29422, QN => n32690);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n27944, QN => n32691);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n27945, QN => n32692);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n27946, QN => n32693);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n27947, QN => n32694);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n27948, QN => n32695);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n27949, QN => n32696);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n27950, QN => n32697);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n27951, QN => n32698);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n27952, QN => n32699);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n27953, QN => n32700);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n27954, QN => n32701);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n27955, QN => n32702);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n8995, CK => CLK, Q => 
                           n29427, QN => n32703);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n8996, CK => CLK, Q => 
                           n29428, QN => n32704);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n8997, CK => CLK, Q => 
                           n29429, QN => n32705);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n8998, CK => CLK, Q => 
                           n29430, QN => n32706);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n8999, CK => CLK, Q => 
                           n29431, QN => n32707);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n9000, CK => CLK, Q => 
                           n29432, QN => n32708);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n9001, CK => CLK, Q => 
                           n29433, QN => n32709);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n9002, CK => CLK, Q => 
                           n29434, QN => n32710);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n9003, CK => CLK, Q => 
                           n29435, QN => n32711);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n9004, CK => CLK, Q => 
                           n29436, QN => n32712);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n9005, CK => CLK, Q => 
                           n29437, QN => n32713);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n9006, CK => CLK, Q => 
                           n29438, QN => n32714);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n8931, CK => CLK, Q => 
                           n29363, QN => n32715);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n8932, CK => CLK, Q => 
                           n29364, QN => n32716);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n8933, CK => CLK, Q => 
                           n29365, QN => n32717);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n8934, CK => CLK, Q => 
                           n29366, QN => n32718);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n8935, CK => CLK, Q => 
                           n29367, QN => n32719);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n8936, CK => CLK, Q => 
                           n29368, QN => n32720);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n8937, CK => CLK, Q => 
                           n29369, QN => n32721);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n8938, CK => CLK, Q => 
                           n29370, QN => n32722);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n8939, CK => CLK, Q => 
                           n29371, QN => n32723);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n8940, CK => CLK, Q => 
                           n29372, QN => n32724);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n8941, CK => CLK, Q => 
                           n29373, QN => n32725);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n8942, CK => CLK, Q => 
                           n29374, QN => n32726);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n8687, CK => CLK, Q => 
                           n29119, QN => n32847);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n8688, CK => CLK, Q => 
                           n29120, QN => n32848);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n8689, CK => CLK, Q => 
                           n29121, QN => n32849);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n8690, CK => CLK, Q => 
                           n29122, QN => n32850);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n8691, CK => CLK, Q => 
                           n29123, QN => n32851);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n8692, CK => CLK, Q => 
                           n29124, QN => n32852);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n8693, CK => CLK, Q => 
                           n29125, QN => n32853);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n8694, CK => CLK, Q => 
                           n29126, QN => n32854);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n8695, CK => CLK, Q => 
                           n29127, QN => n32855);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n8696, CK => CLK, Q => 
                           n29128, QN => n32856);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n8697, CK => CLK, Q => 
                           n29129, QN => n32857);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n8698, CK => CLK, Q => 
                           n29130, QN => n32858);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n8699, CK => CLK, Q => 
                           n29131, QN => n32859);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n8700, CK => CLK, Q => 
                           n29132, QN => n32860);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n8701, CK => CLK, Q => 
                           n29133, QN => n32861);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n8702, CK => CLK, Q => 
                           n29134, QN => n32862);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n8703, CK => CLK, Q => 
                           n29135, QN => n32863);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n8704, CK => CLK, Q => 
                           n29136, QN => n32864);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n8705, CK => CLK, Q => 
                           n29137, QN => n32865);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n8706, CK => CLK, Q => 
                           n29138, QN => n32866);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n8707, CK => CLK, Q => 
                           n29139, QN => n32867);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n8708, CK => CLK, Q => 
                           n29140, QN => n32868);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n8709, CK => CLK, Q => 
                           n29141, QN => n32869);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n8710, CK => CLK, Q => 
                           n29142, QN => n32870);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n8711, CK => CLK, Q => 
                           n29143, QN => n32871);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n8712, CK => CLK, Q => 
                           n29144, QN => n32872);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n8713, CK => CLK, Q => 
                           n29145, QN => n32873);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n8714, CK => CLK, Q => 
                           n29146, QN => n32874);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n8715, CK => CLK, Q => 
                           n29147, QN => n32875);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n8716, CK => CLK, Q => 
                           n29148, QN => n32876);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n8717, CK => CLK, Q => 
                           n29149, QN => n32877);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n8718, CK => CLK, Q => 
                           n29150, QN => n32878);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n8719, CK => CLK, Q => 
                           n29151, QN => n32879);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n8720, CK => CLK, Q => 
                           n29152, QN => n32880);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n8721, CK => CLK, Q => 
                           n29153, QN => n32881);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n8722, CK => CLK, Q => 
                           n29154, QN => n32882);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n8723, CK => CLK, Q => 
                           n29155, QN => n32883);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n8724, CK => CLK, Q => 
                           n29156, QN => n32884);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n8725, CK => CLK, Q => 
                           n29157, QN => n32885);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n8726, CK => CLK, Q => 
                           n29158, QN => n32886);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n8727, CK => CLK, Q => 
                           n29159, QN => n32887);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n8728, CK => CLK, Q => 
                           n29160, QN => n32888);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n8729, CK => CLK, Q => 
                           n29161, QN => n32889);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n8730, CK => CLK, Q => 
                           n29162, QN => n32890);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n8731, CK => CLK, Q => 
                           n29163, QN => n32891);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n8732, CK => CLK, Q => 
                           n29164, QN => n32892);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n8733, CK => CLK, Q => 
                           n29165, QN => n32893);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n8734, CK => CLK, Q => 
                           n29166, QN => n32894);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n8623, CK => CLK, Q => 
                           n29055, QN => n32895);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n8624, CK => CLK, Q => 
                           n29056, QN => n32896);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n8625, CK => CLK, Q => 
                           n29057, QN => n32897);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n8626, CK => CLK, Q => 
                           n29058, QN => n32898);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n8627, CK => CLK, Q => 
                           n29059, QN => n32899);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n8628, CK => CLK, Q => 
                           n29060, QN => n32900);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n8629, CK => CLK, Q => 
                           n29061, QN => n32901);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n8630, CK => CLK, Q => 
                           n29062, QN => n32902);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n8631, CK => CLK, Q => 
                           n29063, QN => n32903);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n8632, CK => CLK, Q => 
                           n29064, QN => n32904);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n8633, CK => CLK, Q => 
                           n29065, QN => n32905);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n8634, CK => CLK, Q => 
                           n29066, QN => n32906);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n8635, CK => CLK, Q => 
                           n29067, QN => n32907);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n8636, CK => CLK, Q => 
                           n29068, QN => n32908);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n8637, CK => CLK, Q => 
                           n29069, QN => n32909);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n8638, CK => CLK, Q => 
                           n29070, QN => n32910);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n8639, CK => CLK, Q => 
                           n29071, QN => n32911);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n8640, CK => CLK, Q => 
                           n29072, QN => n32912);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n8641, CK => CLK, Q => 
                           n29073, QN => n32913);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n8642, CK => CLK, Q => 
                           n29074, QN => n32914);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n8643, CK => CLK, Q => 
                           n29075, QN => n32915);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n8644, CK => CLK, Q => 
                           n29076, QN => n32916);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n8645, CK => CLK, Q => 
                           n29077, QN => n32917);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n8646, CK => CLK, Q => 
                           n29078, QN => n32918);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n8647, CK => CLK, Q => 
                           n29079, QN => n32919);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n8648, CK => CLK, Q => 
                           n29080, QN => n32920);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n8649, CK => CLK, Q => 
                           n29081, QN => n32921);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n8650, CK => CLK, Q => 
                           n29082, QN => n32922);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n8651, CK => CLK, Q => 
                           n29083, QN => n32923);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n8652, CK => CLK, Q => 
                           n29084, QN => n32924);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n8653, CK => CLK, Q => 
                           n29085, QN => n32925);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n8654, CK => CLK, Q => 
                           n29086, QN => n32926);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n8655, CK => CLK, Q => 
                           n29087, QN => n32927);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n8656, CK => CLK, Q => 
                           n29088, QN => n32928);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n8657, CK => CLK, Q => 
                           n29089, QN => n32929);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n8658, CK => CLK, Q => 
                           n29090, QN => n32930);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n8659, CK => CLK, Q => 
                           n29091, QN => n32931);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n8660, CK => CLK, Q => 
                           n29092, QN => n32932);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n8661, CK => CLK, Q => 
                           n29093, QN => n32933);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n8662, CK => CLK, Q => 
                           n29094, QN => n32934);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n8663, CK => CLK, Q => 
                           n29095, QN => n32935);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n8664, CK => CLK, Q => 
                           n29096, QN => n32936);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n8665, CK => CLK, Q => 
                           n29097, QN => n32937);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n8666, CK => CLK, Q => 
                           n29098, QN => n32938);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n8667, CK => CLK, Q => 
                           n29099, QN => n32939);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n8668, CK => CLK, Q => 
                           n29100, QN => n32940);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n8669, CK => CLK, Q => 
                           n29101, QN => n32941);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n8670, CK => CLK, Q => 
                           n29102, QN => n32942);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n9263, CK => CLK, Q => 
                           n29695, QN => n38982);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n9264, CK => CLK, Q => 
                           n29696, QN => n38981);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n9265, CK => CLK, Q => 
                           n29697, QN => n38980);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n9266, CK => CLK, Q => 
                           n29698, QN => n38979);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n9267, CK => CLK, Q => 
                           n29699, QN => n38978);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n9268, CK => CLK, Q => 
                           n29700, QN => n38977);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n9269, CK => CLK, Q => 
                           n29701, QN => n38976);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n9270, CK => CLK, Q => 
                           n29702, QN => n38975);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n9271, CK => CLK, Q => 
                           n29703, QN => n38974);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n9272, CK => CLK, Q => 
                           n29704, QN => n38973);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n9273, CK => CLK, Q => 
                           n29705, QN => n38972);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n9274, CK => CLK, Q => 
                           n29706, QN => n38971);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n9275, CK => CLK, Q => 
                           n29707, QN => n38970);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n9276, CK => CLK, Q => 
                           n29708, QN => n38969);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n9277, CK => CLK, Q => 
                           n29709, QN => n38968);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n9278, CK => CLK, Q => 
                           n29710, QN => n38967);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n9279, CK => CLK, Q => 
                           n29711, QN => n38966);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n9280, CK => CLK, Q => 
                           n29712, QN => n38965);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n9281, CK => CLK, Q => 
                           n29713, QN => n38964);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n9282, CK => CLK, Q => 
                           n29714, QN => n38963);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n9283, CK => CLK, Q => 
                           n29715, QN => n38962);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n9284, CK => CLK, Q => 
                           n29716, QN => n38961);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n9285, CK => CLK, Q => 
                           n29717, QN => n38960);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n9286, CK => CLK, Q => 
                           n29718, QN => n38959);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n9287, CK => CLK, Q => 
                           n29719, QN => n38958);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n9288, CK => CLK, Q => 
                           n29720, QN => n38957);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n9289, CK => CLK, Q => 
                           n29721, QN => n38956);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n9290, CK => CLK, Q => 
                           n29722, QN => n38955);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n9291, CK => CLK, Q => 
                           n29723, QN => n38954);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n9292, CK => CLK, Q => 
                           n29724, QN => n38953);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n9293, CK => CLK, Q => 
                           n29725, QN => n38952);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n9294, CK => CLK, Q => 
                           n29726, QN => n38951);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n9295, CK => CLK, Q => 
                           n29727, QN => n38950);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n9296, CK => CLK, Q => 
                           n29728, QN => n38949);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n9297, CK => CLK, Q => 
                           n29729, QN => n38948);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n9298, CK => CLK, Q => 
                           n29730, QN => n38947);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n9299, CK => CLK, Q => 
                           n29731, QN => n38946);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n9300, CK => CLK, Q => 
                           n29732, QN => n38945);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n9301, CK => CLK, Q => 
                           n29733, QN => n38944);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n9302, CK => CLK, Q => 
                           n29734, QN => n38943);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n9303, CK => CLK, Q => 
                           n29735, QN => n38942);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n9304, CK => CLK, Q => 
                           n29736, QN => n38941);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n9305, CK => CLK, Q => 
                           n29737, QN => n38940);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n9306, CK => CLK, Q => 
                           n29738, QN => n38939);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n9307, CK => CLK, Q => 
                           n29739, QN => n38938);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n9308, CK => CLK, Q => 
                           n29740, QN => n38937);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n9309, CK => CLK, Q => 
                           n29741, QN => n38936);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n9310, CK => CLK, Q => 
                           n29742, QN => n38935);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n8675, CK => CLK, Q => 
                           n29107, QN => n33087);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n8676, CK => CLK, Q => 
                           n29108, QN => n33088);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n8677, CK => CLK, Q => 
                           n29109, QN => n33089);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n8678, CK => CLK, Q => 
                           n29110, QN => n33090);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n8679, CK => CLK, Q => 
                           n29111, QN => n33091);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n8680, CK => CLK, Q => 
                           n29112, QN => n33092);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n8681, CK => CLK, Q => 
                           n29113, QN => n33093);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n8682, CK => CLK, Q => 
                           n29114, QN => n33094);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n8683, CK => CLK, Q => 
                           n29115, QN => n33095);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n8684, CK => CLK, Q => 
                           n29116, QN => n33096);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n8685, CK => CLK, Q => 
                           n29117, QN => n33097);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n8686, CK => CLK, Q => 
                           n29118, QN => n33098);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n8611, CK => CLK, Q => 
                           n29043, QN => n33099);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n8612, CK => CLK, Q => 
                           n29044, QN => n33100);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n8613, CK => CLK, Q => 
                           n29045, QN => n33101);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n8614, CK => CLK, Q => 
                           n29046, QN => n33102);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n8615, CK => CLK, Q => 
                           n29047, QN => n33103);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n8616, CK => CLK, Q => 
                           n29048, QN => n33104);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n8617, CK => CLK, Q => 
                           n29049, QN => n33105);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n8618, CK => CLK, Q => 
                           n29050, QN => n33106);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n8619, CK => CLK, Q => 
                           n29051, QN => n33107);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n8620, CK => CLK, Q => 
                           n29052, QN => n33108);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n8621, CK => CLK, Q => 
                           n29053, QN => n33109);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n8622, CK => CLK, Q => 
                           n29054, QN => n33110);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n9251, CK => CLK, Q => 
                           n29683, QN => n33135);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n9252, CK => CLK, Q => 
                           n29684, QN => n33136);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n9253, CK => CLK, Q => 
                           n29685, QN => n33137);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n9254, CK => CLK, Q => 
                           n29686, QN => n38934);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n9255, CK => CLK, Q => 
                           n29687, QN => n33139);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n9256, CK => CLK, Q => 
                           n29688, QN => n38933);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n9257, CK => CLK, Q => 
                           n29689, QN => n38932);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n9258, CK => CLK, Q => 
                           n29690, QN => n38931);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n9259, CK => CLK, Q => 
                           n29691, QN => n38930);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n9260, CK => CLK, Q => 
                           n29692, QN => n38929);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n9261, CK => CLK, Q => 
                           n29693, QN => n38928);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n9262, CK => CLK, Q => 
                           n29694, QN => n38927);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n9327, CK => CLK, Q => 
                           n29759, QN => n38849);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n9328, CK => CLK, Q => 
                           n29760, QN => n38848);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n9329, CK => CLK, Q => 
                           n29761, QN => n38847);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n9330, CK => CLK, Q => 
                           n29762, QN => n38846);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n9331, CK => CLK, Q => 
                           n29763, QN => n38845);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n9332, CK => CLK, Q => 
                           n29764, QN => n38844);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n9333, CK => CLK, Q => 
                           n29765, QN => n38843);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n9334, CK => CLK, Q => 
                           n29766, QN => n38842);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n9335, CK => CLK, Q => 
                           n29767, QN => n38841);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n9336, CK => CLK, Q => 
                           n29768, QN => n38840);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n9337, CK => CLK, Q => 
                           n29769, QN => n38839);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n9338, CK => CLK, Q => 
                           n29770, QN => n38838);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n9339, CK => CLK, Q => 
                           n29771, QN => n38837);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n9340, CK => CLK, Q => 
                           n29772, QN => n38836);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n9341, CK => CLK, Q => 
                           n29773, QN => n38835);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n9342, CK => CLK, Q => 
                           n29774, QN => n38834);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n9343, CK => CLK, Q => 
                           n29775, QN => n38833);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n9344, CK => CLK, Q => 
                           n29776, QN => n38832);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n9345, CK => CLK, Q => 
                           n29777, QN => n38831);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n9346, CK => CLK, Q => 
                           n29778, QN => n38830);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n9347, CK => CLK, Q => 
                           n29779, QN => n38829);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n9348, CK => CLK, Q => 
                           n29780, QN => n38828);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n9349, CK => CLK, Q => 
                           n29781, QN => n38827);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n9350, CK => CLK, Q => 
                           n29782, QN => n38826);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n9351, CK => CLK, Q => 
                           n29783, QN => n38825);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n9352, CK => CLK, Q => 
                           n29784, QN => n38824);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n9353, CK => CLK, Q => 
                           n29785, QN => n38823);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n9354, CK => CLK, Q => 
                           n29786, QN => n38822);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n9355, CK => CLK, Q => 
                           n29787, QN => n38821);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n9356, CK => CLK, Q => 
                           n29788, QN => n38820);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n9357, CK => CLK, Q => 
                           n29789, QN => n38819);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n9358, CK => CLK, Q => 
                           n29790, QN => n38818);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n9359, CK => CLK, Q => 
                           n29791, QN => n38817);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n9360, CK => CLK, Q => 
                           n29792, QN => n38816);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n9361, CK => CLK, Q => 
                           n29793, QN => n38815);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n9362, CK => CLK, Q => 
                           n29794, QN => n38814);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n9363, CK => CLK, Q => 
                           n29795, QN => n38813);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n9364, CK => CLK, Q => 
                           n29796, QN => n38812);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n9365, CK => CLK, Q => 
                           n29797, QN => n38811);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n9366, CK => CLK, Q => 
                           n29798, QN => n38810);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n9367, CK => CLK, Q => 
                           n29799, QN => n38809);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n9368, CK => CLK, Q => 
                           n29800, QN => n38808);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n9369, CK => CLK, Q => 
                           n29801, QN => n38807);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n9370, CK => CLK, Q => 
                           n29802, QN => n38806);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n9371, CK => CLK, Q => 
                           n29803, QN => n38805);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n9372, CK => CLK, Q => 
                           n29804, QN => n38804);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n9373, CK => CLK, Q => 
                           n29805, QN => n38803);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n9374, CK => CLK, Q => 
                           n29806, QN => n38802);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n9315, CK => CLK, Q => 
                           n29747, QN => n33195);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n9316, CK => CLK, Q => 
                           n29748, QN => n33196);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n9317, CK => CLK, Q => 
                           n29749, QN => n33197);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n9318, CK => CLK, Q => 
                           n29750, QN => n38801);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n9319, CK => CLK, Q => 
                           n29751, QN => n33199);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n9320, CK => CLK, Q => 
                           n29752, QN => n38800);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n9321, CK => CLK, Q => 
                           n29753, QN => n38799);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n9322, CK => CLK, Q => 
                           n29754, QN => n38798);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n9323, CK => CLK, Q => 
                           n29755, QN => n38797);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n9324, CK => CLK, Q => 
                           n29756, QN => n38796);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n9325, CK => CLK, Q => 
                           n29757, QN => n38795);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n9326, CK => CLK, Q => 
                           n29758, QN => n38794);
   U26382 : NAND3_X1 port map( A1 => n33212, A2 => n41370, A3 => n2695, ZN => 
                           n33214);
   U26383 : XOR2_X1 port map( A => n32323, B => n2683, Z => n33241);
   U26384 : NAND3_X1 port map( A1 => n33249, A2 => n32255, A3 => n2709, ZN => 
                           n33248);
   U26385 : NAND3_X1 port map( A1 => n32153, A2 => n40581, A3 => n33257, ZN => 
                           n33252);
   U26386 : NAND3_X1 port map( A1 => n33257, A2 => n40561, A3 => n32154, ZN => 
                           n33261);
   U26387 : NAND3_X1 port map( A1 => n33257, A2 => n40541, A3 => n32155, ZN => 
                           n33266);
   U26388 : NAND3_X1 port map( A1 => n33257, A2 => n40521, A3 => n32156, ZN => 
                           n33271);
   U26389 : NAND3_X1 port map( A1 => n33257, A2 => n40501, A3 => n33279, ZN => 
                           n33276);
   U26390 : NAND3_X1 port map( A1 => n33257, A2 => n40481, A3 => n33284, ZN => 
                           n33281);
   U26391 : NAND3_X1 port map( A1 => n33257, A2 => n40461, A3 => n33289, ZN => 
                           n33286);
   U26392 : NAND3_X1 port map( A1 => WR, A2 => n32150, A3 => n33294, ZN => 
                           n33256);
   U26393 : NAND3_X1 port map( A1 => n33257, A2 => n40441, A3 => n33295, ZN => 
                           n33291);
   U26394 : NAND3_X1 port map( A1 => n33297, A2 => ENABLE, A3 => n33298, ZN => 
                           n33259);
   U26395 : NAND3_X1 port map( A1 => n33294, A2 => n32150, A3 => n33299, ZN => 
                           n33258);
   U26396 : NAND3_X1 port map( A1 => n32153, A2 => n40421, A3 => n33306, ZN => 
                           n33302);
   U26397 : NAND3_X1 port map( A1 => n32154, A2 => n40401, A3 => n33306, ZN => 
                           n33309);
   U26398 : NAND3_X1 port map( A1 => n32155, A2 => n40381, A3 => n33306, ZN => 
                           n33312);
   U26399 : NAND3_X1 port map( A1 => n32156, A2 => n40361, A3 => n33306, ZN => 
                           n33315);
   U26400 : NAND3_X1 port map( A1 => n33279, A2 => n40341, A3 => n33306, ZN => 
                           n33318);
   U26401 : NAND3_X1 port map( A1 => n33284, A2 => n40321, A3 => n33306, ZN => 
                           n33321);
   U26402 : NAND3_X1 port map( A1 => n33289, A2 => n40301, A3 => n33306, ZN => 
                           n33324);
   U26403 : NAND3_X1 port map( A1 => N932, A2 => N931, A3 => n33330, ZN => 
                           n33305);
   U26404 : NAND3_X1 port map( A1 => n33295, A2 => n40281, A3 => n33306, ZN => 
                           n33327);
   U26405 : NAND3_X1 port map( A1 => n32239, A2 => n33332, A3 => N813, ZN => 
                           n33308);
   U26406 : NAND3_X1 port map( A1 => N931, A2 => n33333, A3 => N932, ZN => 
                           n33307);
   U26407 : NAND3_X1 port map( A1 => n32153, A2 => n40261, A3 => n33338, ZN => 
                           n33334);
   U26408 : NAND3_X1 port map( A1 => n32154, A2 => n40241, A3 => n33338, ZN => 
                           n33341);
   U26409 : NAND3_X1 port map( A1 => n32155, A2 => n40221, A3 => n33338, ZN => 
                           n33344);
   U26410 : NAND3_X1 port map( A1 => n32156, A2 => n40201, A3 => n33338, ZN => 
                           n33347);
   U26411 : NAND3_X1 port map( A1 => n33279, A2 => n40181, A3 => n33338, ZN => 
                           n33350);
   U26412 : NAND3_X1 port map( A1 => n33284, A2 => n40161, A3 => n33338, ZN => 
                           n33353);
   U26413 : NAND3_X1 port map( A1 => n33289, A2 => n40141, A3 => n33338, ZN => 
                           n33356);
   U26414 : NAND3_X1 port map( A1 => N932, A2 => n32152, A3 => n33330, ZN => 
                           n33337);
   U26415 : NAND3_X1 port map( A1 => n33295, A2 => n40121, A3 => n33338, ZN => 
                           n33359);
   U26416 : NAND3_X1 port map( A1 => n32239, A2 => n32247, A3 => n33332, ZN => 
                           n33340);
   U26417 : NAND3_X1 port map( A1 => n33333, A2 => n32152, A3 => N932, ZN => 
                           n33339);
   U26418 : NAND3_X1 port map( A1 => n32153, A2 => n40101, A3 => n33367, ZN => 
                           n33363);
   U26419 : NAND3_X1 port map( A1 => n32154, A2 => n40082, A3 => n33367, ZN => 
                           n33370);
   U26420 : NAND3_X1 port map( A1 => n32155, A2 => n40062, A3 => n33367, ZN => 
                           n33373);
   U26421 : NAND3_X1 port map( A1 => n32156, A2 => n40042, A3 => n33367, ZN => 
                           n33376);
   U26422 : NAND3_X1 port map( A1 => n33279, A2 => n40021, A3 => n33367, ZN => 
                           n33379);
   U26423 : NAND3_X1 port map( A1 => n33284, A2 => n40002, A3 => n33367, ZN => 
                           n33382);
   U26424 : NAND3_X1 port map( A1 => n33289, A2 => n39984, A3 => n33367, ZN => 
                           n33385);
   U26425 : NAND3_X1 port map( A1 => N931, A2 => n32151, A3 => n33330, ZN => 
                           n33366);
   U26426 : NAND3_X1 port map( A1 => n33295, A2 => n39964, A3 => n33367, ZN => 
                           n33388);
   U26427 : NAND3_X1 port map( A1 => n33332, A2 => n33362, A3 => N813, ZN => 
                           n33369);
   U26428 : NAND3_X1 port map( A1 => n33333, A2 => n32151, A3 => N931, ZN => 
                           n33368);
   U26429 : NAND3_X1 port map( A1 => n32153, A2 => n39944, A3 => n33395, ZN => 
                           n33391);
   U26430 : NAND3_X1 port map( A1 => N811, A2 => n33398, A3 => N812, ZN => 
                           n33260);
   U26432 : NAND3_X1 port map( A1 => n32154, A2 => n39923, A3 => n33395, ZN => 
                           n33399);
   U26433 : NAND3_X1 port map( A1 => N812, A2 => N811, A3 => n32254, ZN => 
                           n33265);
   U26434 : NAND3_X1 port map( A1 => N930, A2 => N929, A3 => n33402, ZN => 
                           n33264);
   U26435 : NAND3_X1 port map( A1 => n32155, A2 => n39904, A3 => n33395, ZN => 
                           n33403);
   U26436 : NAND3_X1 port map( A1 => n33398, A2 => n32251, A3 => N812, ZN => 
                           n33270);
   U26437 : NAND3_X1 port map( A1 => n32163, A2 => n32161, A3 => N930, ZN => 
                           n33269);
   U26438 : NAND3_X1 port map( A1 => n32156, A2 => n39886, A3 => n33395, ZN => 
                           n33406);
   U26439 : NAND3_X1 port map( A1 => N812, A2 => n32251, A3 => n32254, ZN => 
                           n33275);
   U26440 : NAND3_X1 port map( A1 => N930, A2 => n32161, A3 => n33402, ZN => 
                           n33274);
   U26441 : NAND3_X1 port map( A1 => n33279, A2 => n39866, A3 => n33395, ZN => 
                           n33409);
   U26442 : NAND3_X1 port map( A1 => n33398, A2 => n32249, A3 => N811, ZN => 
                           n33280);
   U26443 : NAND3_X1 port map( A1 => n33284, A2 => n39846, A3 => n33395, ZN => 
                           n33412);
   U26444 : NAND3_X1 port map( A1 => N811, A2 => n32249, A3 => n32254, ZN => 
                           n33285);
   U26445 : NAND3_X1 port map( A1 => n33289, A2 => n39826, A3 => n33395, ZN => 
                           n33415);
   U26446 : NAND3_X1 port map( A1 => n32251, A2 => n32249, A3 => n33398, ZN => 
                           n33290);
   U26447 : NAND3_X1 port map( A1 => n33295, A2 => n39804, A3 => n33395, ZN => 
                           n33418);
   U26448 : NAND3_X1 port map( A1 => n33362, A2 => n32247, A3 => n33332, ZN => 
                           n33396);
   U26449 : XOR2_X1 port map( A => add_146_carry_4_port, B => n2695, Z => 
                           n33362);
   U26450 : NAND3_X1 port map( A1 => n32251, A2 => n32249, A3 => n32254, ZN => 
                           n33296);
   U26451 : XOR2_X1 port map( A => n33422, B => r498_carry_5_port, Z => n33301)
                           ;
   U26452 : XOR2_X1 port map( A => n33423, B => ADD_WR(0), Z => n33402);
   U26453 : XOR2_X1 port map( A => n34696, B => ADD_RD1(0), Z => n34694);
   U26454 : XOR2_X1 port map( A => n35970, B => ADD_RD2(0), Z => n35968);
   U26455 : XOR2_X1 port map( A => n27874, B => n2697, Z => n33243);
   U26456 : XOR2_X1 port map( A => n27871, B => n2699, Z => n33242);
   U26457 : XOR2_X1 port map( A => n27870, B => n33215, Z => n35978);
   U26458 : XOR2_X1 port map( A => n32258, B => N661, Z => n33245);
   U26459 : XOR2_X1 port map( A => n38790, B => n2698, Z => n33239);
   U26460 : XOR2_X1 port map( A => add_136_carry_4_port, B => n2695, Z => 
                           n37240);
   U26461 : NAND3_X1 port map( A1 => i_1_port, A2 => n32255, A3 => n33249, ZN 
                           => n33250);
   CWP_reg_3_inst : DFF_X1 port map( D => n9904, CK => CLK, Q => N661, QN => 
                           n2696);
   CWP_reg_2_inst : DFF_X1 port map( D => n9905, CK => CLK, Q => N660, QN => 
                           n2697);
   CWP_reg_1_inst : DFF_X1 port map( D => n9906, CK => CLK, Q => N659, QN => 
                           n2698);
   i_reg_3_inst : DFF_X1 port map( D => n25394, CK => CLK, Q => i_3_port, QN =>
                           n2706);
   i_reg_1_inst : DFF_X1 port map( D => n9892, CK => CLK, Q => i_1_port, QN => 
                           n2709);
   i_reg_2_inst : DFF_X1 port map( D => n9891, CK => CLK, Q => i_2_port, QN => 
                           n2707);
   STORE_DATA_reg : DFF_X1 port map( D => n7202, CK => CLK, Q => SPILL, QN => 
                           n2700);
   RETRIEVE_DATA_reg : DFF_X1 port map( D => n9893, CK => CLK, Q => FILL, QN =>
                           n23853);
   BUSout_reg_63_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => BUSout(63)
                           , QN => n16941);
   BUSout_reg_62_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => BUSout(62)
                           , QN => n16940);
   BUSout_reg_61_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => BUSout(61)
                           , QN => n16939);
   BUSout_reg_60_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => BUSout(60)
                           , QN => n16938);
   BUSout_reg_5_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => BUSout(5), 
                           QN => n16883);
   BUSout_reg_4_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => BUSout(4), 
                           QN => n16882);
   BUSout_reg_3_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => BUSout(3), 
                           QN => n16881);
   BUSout_reg_2_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => BUSout(2), 
                           QN => n16880);
   BUSout_reg_1_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => BUSout(1), 
                           QN => n16879);
   BUSout_reg_53_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => BUSout(53)
                           , QN => n16931);
   BUSout_reg_52_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => BUSout(52)
                           , QN => n16930);
   BUSout_reg_51_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => BUSout(51)
                           , QN => n16929);
   BUSout_reg_50_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => BUSout(50)
                           , QN => n16928);
   BUSout_reg_49_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => BUSout(49)
                           , QN => n16927);
   BUSout_reg_48_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => BUSout(48)
                           , QN => n16926);
   BUSout_reg_47_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => BUSout(47)
                           , QN => n16925);
   BUSout_reg_46_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => BUSout(46)
                           , QN => n16924);
   BUSout_reg_45_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => BUSout(45)
                           , QN => n16923);
   BUSout_reg_44_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => BUSout(44)
                           , QN => n16922);
   BUSout_reg_43_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => BUSout(43)
                           , QN => n16921);
   BUSout_reg_42_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => BUSout(42)
                           , QN => n16920);
   BUSout_reg_41_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => BUSout(41)
                           , QN => n16919);
   BUSout_reg_40_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => BUSout(40)
                           , QN => n16918);
   BUSout_reg_39_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => BUSout(39)
                           , QN => n16917);
   BUSout_reg_38_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => BUSout(38)
                           , QN => n16916);
   BUSout_reg_37_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => BUSout(37)
                           , QN => n16915);
   BUSout_reg_36_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => BUSout(36)
                           , QN => n16914);
   BUSout_reg_35_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => BUSout(35)
                           , QN => n16913);
   BUSout_reg_34_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => BUSout(34)
                           , QN => n16912);
   BUSout_reg_33_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => BUSout(33)
                           , QN => n16911);
   BUSout_reg_32_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => BUSout(32)
                           , QN => n16910);
   BUSout_reg_31_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => BUSout(31)
                           , QN => n16909);
   BUSout_reg_30_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => BUSout(30)
                           , QN => n16908);
   BUSout_reg_29_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => BUSout(29)
                           , QN => n16907);
   BUSout_reg_28_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => BUSout(28)
                           , QN => n16906);
   BUSout_reg_27_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => BUSout(27)
                           , QN => n16905);
   BUSout_reg_26_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => BUSout(26)
                           , QN => n16904);
   BUSout_reg_25_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => BUSout(25)
                           , QN => n16903);
   BUSout_reg_24_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => BUSout(24)
                           , QN => n16902);
   BUSout_reg_23_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => BUSout(23)
                           , QN => n16901);
   BUSout_reg_22_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => BUSout(22)
                           , QN => n16900);
   BUSout_reg_21_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => BUSout(21)
                           , QN => n16899);
   BUSout_reg_20_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => BUSout(20)
                           , QN => n16898);
   BUSout_reg_19_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => BUSout(19)
                           , QN => n16897);
   BUSout_reg_18_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => BUSout(18)
                           , QN => n16896);
   BUSout_reg_17_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => BUSout(17)
                           , QN => n16895);
   BUSout_reg_16_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => BUSout(16)
                           , QN => n16894);
   BUSout_reg_15_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => BUSout(15)
                           , QN => n16893);
   BUSout_reg_14_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => BUSout(14)
                           , QN => n16892);
   BUSout_reg_13_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => BUSout(13)
                           , QN => n16891);
   BUSout_reg_12_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => BUSout(12)
                           , QN => n16890);
   BUSout_reg_11_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => BUSout(11)
                           , QN => n16889);
   BUSout_reg_10_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => BUSout(10)
                           , QN => n16888);
   BUSout_reg_9_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => BUSout(9), 
                           QN => n16887);
   BUSout_reg_8_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => BUSout(8), 
                           QN => n16886);
   BUSout_reg_7_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => BUSout(7), 
                           QN => n16885);
   BUSout_reg_6_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => BUSout(6), 
                           QN => n16884);
   SWP_reg_4_inst : DFF_X1 port map( D => n9896, CK => CLK, Q => n27872, QN => 
                           n32322);
   SWP_reg_3_inst : DFF_X1 port map( D => n9897, CK => CLK, Q => n38789, QN => 
                           n32258);
   SWP_reg_1_inst : DFF_X1 port map( D => n9899, CK => CLK, Q => n38790, QN => 
                           n32260);
   SWP_reg_5_inst : DFF_X1 port map( D => n9901, CK => CLK, Q => n27870, QN => 
                           n32323);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7583, CK => CLK, Q => n_2480
                           , QN => n30605);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7584, CK => CLK, Q => n_2481
                           , QN => n30606);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7585, CK => CLK, Q => n_2482
                           , QN => n30607);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7586, CK => CLK, Q => n_2483
                           , QN => n30608);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7519, CK => CLK, Q => n_2484
                           , QN => n30541);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7520, CK => CLK, Q => n_2485
                           , QN => n30542);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7521, CK => CLK, Q => n_2486
                           , QN => n30543);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7522, CK => CLK, Q => n_2487
                           , QN => n30544);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => n28004
                           , QN => n32456);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => n28005
                           , QN => n32457);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => n28006
                           , QN => n32458);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => n28007
                           , QN => n32459);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7647, CK => CLK, Q => n_2488
                           , QN => n30669);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7648, CK => CLK, Q => n_2489
                           , QN => n30670);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7649, CK => CLK, Q => n_2490
                           , QN => n30671);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7650, CK => CLK, Q => n_2491
                           , QN => n30672);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n7839, CK => CLK, Q => n_2492
                           , QN => n30733);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n7840, CK => CLK, Q => n_2493
                           , QN => n30734);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n7841, CK => CLK, Q => n_2494
                           , QN => n30735);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n7842, CK => CLK, Q => n_2495
                           , QN => n30736);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n7967, CK => CLK, Q => n_2496
                           , QN => n30861);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n7968, CK => CLK, Q => n_2497
                           , QN => n30862);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n7969, CK => CLK, Q => n_2498
                           , QN => n30863);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n7970, CK => CLK, Q => n_2499
                           , QN => n30864);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n7903, CK => CLK, Q => n_2500
                           , QN => n30797);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n7904, CK => CLK, Q => n_2501
                           , QN => n30798);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n7905, CK => CLK, Q => n_2502
                           , QN => n30799);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n7906, CK => CLK, Q => n_2503
                           , QN => n30800);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n8607, CK => CLK, Q => 
                           n_2504, QN => n31363);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n8608, CK => CLK, Q => 
                           n_2505, QN => n31364);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n8609, CK => CLK, Q => 
                           n_2506, QN => n31365);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n8610, CK => CLK, Q => 
                           n_2507, QN => n31366);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n8543, CK => CLK, Q => 
                           n_2508, QN => n31299);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n8544, CK => CLK, Q => 
                           n_2509, QN => n31300);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n8545, CK => CLK, Q => 
                           n_2510, QN => n31301);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n8546, CK => CLK, Q => 
                           n_2511, QN => n31302);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n8479, CK => CLK, Q => 
                           n_2512, QN => n31235);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n8480, CK => CLK, Q => 
                           n_2513, QN => n31236);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n8481, CK => CLK, Q => 
                           n_2514, QN => n31237);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n8482, CK => CLK, Q => 
                           n_2515, QN => n31238);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7526, CK => CLK, Q => 
                           n_2516, QN => n30548);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7528, CK => CLK, Q => 
                           n_2517, QN => n30550);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7529, CK => CLK, Q => 
                           n_2518, QN => n30551);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7530, CK => CLK, Q => 
                           n_2519, QN => n30552);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7531, CK => CLK, Q => 
                           n_2520, QN => n30553);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7532, CK => CLK, Q => 
                           n_2521, QN => n30554);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7533, CK => CLK, Q => 
                           n_2522, QN => n30555);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7534, CK => CLK, Q => 
                           n_2523, QN => n30556);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7535, CK => CLK, Q => 
                           n_2524, QN => n30557);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7536, CK => CLK, Q => 
                           n_2525, QN => n30558);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7537, CK => CLK, Q => 
                           n_2526, QN => n30559);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7538, CK => CLK, Q => 
                           n_2527, QN => n30560);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7539, CK => CLK, Q => 
                           n_2528, QN => n30561);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7540, CK => CLK, Q => 
                           n_2529, QN => n30562);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7541, CK => CLK, Q => 
                           n_2530, QN => n30563);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7542, CK => CLK, Q => 
                           n_2531, QN => n30564);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7543, CK => CLK, Q => 
                           n_2532, QN => n30565);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7544, CK => CLK, Q => 
                           n_2533, QN => n30566);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7545, CK => CLK, Q => 
                           n_2534, QN => n30567);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7546, CK => CLK, Q => 
                           n_2535, QN => n30568);
   CWP_reg_4_inst : DFF_X1 port map( D => n9903, CK => CLK, Q => n32242, QN => 
                           n2695);
   CWP_reg_5_inst : DFF_X1 port map( D => n9902, CK => CLK, Q => n32244, QN => 
                           n2683);
   i_reg_0_inst : DFF_X1 port map( D => n9895, CK => CLK, Q => n32255, QN => 
                           n2710);
   CWP_reg_0_inst : DFF_X1 port map( D => n9907, CK => CLK, Q => n32253, QN => 
                           n2699);
   SWP_reg_2_inst : DFF_X1 port map( D => n9898, CK => CLK, Q => n32259, QN => 
                           n27874);
   SWP_reg_0_inst : DFF_X1 port map( D => n9900, CK => CLK, Q => n32261, QN => 
                           n27871);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7775, CK => CLK, Q => n32484
                           , QN => n503);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7776, CK => CLK, Q => n32485
                           , QN => n504);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7777, CK => CLK, Q => n32486
                           , QN => n505);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7778, CK => CLK, Q => n32487
                           , QN => n506);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7711, CK => CLK, Q => n32488
                           , QN => n439);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7712, CK => CLK, Q => n32489
                           , QN => n440);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7713, CK => CLK, Q => n32490
                           , QN => n441);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7714, CK => CLK, Q => n32491
                           , QN => n442);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => n30477
                           , QN => n27940);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => n30478
                           , QN => n27941);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => n30479
                           , QN => n27942);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => n30480
                           , QN => n27943);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n8095, CK => CLK, Q => 
                           n32468, QN => n823);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n8096, CK => CLK, Q => 
                           n32469, QN => n824);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n8097, CK => CLK, Q => 
                           n32470, QN => n825);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n8098, CK => CLK, Q => 
                           n32471, QN => n826);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n8031, CK => CLK, Q => 
                           n32472, QN => n759);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n8032, CK => CLK, Q => 
                           n32473, QN => n760);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n8033, CK => CLK, Q => 
                           n32474, QN => n761);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n8034, CK => CLK, Q => 
                           n32475, QN => n762);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n8351, CK => CLK, Q => 
                           n31117, QN => n25401);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n8352, CK => CLK, Q => 
                           n31118, QN => n25400);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n8353, CK => CLK, Q => 
                           n31119, QN => n25399);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n8354, CK => CLK, Q => 
                           n31120, QN => n25398);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7727, CK => CLK, Q => 
                           n32943, QN => n455);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7728, CK => CLK, Q => 
                           n32944, QN => n456);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7729, CK => CLK, Q => 
                           n32945, QN => n457);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7730, CK => CLK, Q => 
                           n32946, QN => n458);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7731, CK => CLK, Q => 
                           n32947, QN => n459);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7732, CK => CLK, Q => 
                           n32948, QN => n460);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7733, CK => CLK, Q => 
                           n32949, QN => n461);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7734, CK => CLK, Q => 
                           n32950, QN => n462);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7735, CK => CLK, Q => 
                           n32951, QN => n463);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7736, CK => CLK, Q => 
                           n32952, QN => n464);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7737, CK => CLK, Q => 
                           n32953, QN => n465);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7738, CK => CLK, Q => 
                           n32954, QN => n466);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7739, CK => CLK, Q => 
                           n32955, QN => n467);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7740, CK => CLK, Q => 
                           n32956, QN => n468);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7741, CK => CLK, Q => 
                           n32957, QN => n469);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7742, CK => CLK, Q => 
                           n32958, QN => n470);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7743, CK => CLK, Q => 
                           n32959, QN => n471);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7744, CK => CLK, Q => 
                           n32960, QN => n472);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7745, CK => CLK, Q => 
                           n32961, QN => n473);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7746, CK => CLK, Q => 
                           n32962, QN => n474);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7747, CK => CLK, Q => 
                           n32963, QN => n475);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7748, CK => CLK, Q => 
                           n32964, QN => n476);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7749, CK => CLK, Q => 
                           n32965, QN => n477);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7750, CK => CLK, Q => 
                           n32966, QN => n478);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7751, CK => CLK, Q => 
                           n32967, QN => n479);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7752, CK => CLK, Q => 
                           n32968, QN => n480);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7753, CK => CLK, Q => 
                           n32969, QN => n481);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7754, CK => CLK, Q => 
                           n32970, QN => n482);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7755, CK => CLK, Q => 
                           n32971, QN => n483);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7756, CK => CLK, Q => 
                           n32972, QN => n484);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7757, CK => CLK, Q => 
                           n32973, QN => n485);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7758, CK => CLK, Q => 
                           n32974, QN => n486);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7759, CK => CLK, Q => 
                           n32975, QN => n487);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7760, CK => CLK, Q => 
                           n32976, QN => n488);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7761, CK => CLK, Q => 
                           n32977, QN => n489);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7762, CK => CLK, Q => 
                           n32978, QN => n490);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7763, CK => CLK, Q => 
                           n32979, QN => n491);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7764, CK => CLK, Q => 
                           n32980, QN => n492);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7765, CK => CLK, Q => 
                           n32981, QN => n493);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7766, CK => CLK, Q => 
                           n32982, QN => n494);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7767, CK => CLK, Q => 
                           n32983, QN => n495);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7768, CK => CLK, Q => 
                           n32984, QN => n496);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7769, CK => CLK, Q => n32985
                           , QN => n497);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7770, CK => CLK, Q => n32986
                           , QN => n498);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7771, CK => CLK, Q => n32987
                           , QN => n499);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7772, CK => CLK, Q => n32988
                           , QN => n500);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7773, CK => CLK, Q => n32989
                           , QN => n501);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7774, CK => CLK, Q => n32990
                           , QN => n502);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7715, CK => CLK, Q => 
                           n33111, QN => n443);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7716, CK => CLK, Q => 
                           n33112, QN => n444);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7717, CK => CLK, Q => 
                           n33113, QN => n445);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7718, CK => CLK, Q => 
                           n33114, QN => n446);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7719, CK => CLK, Q => 
                           n33115, QN => n447);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7720, CK => CLK, Q => 
                           n33116, QN => n448);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7721, CK => CLK, Q => 
                           n33117, QN => n449);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7722, CK => CLK, Q => 
                           n33118, QN => n450);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7723, CK => CLK, Q => 
                           n33119, QN => n451);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7724, CK => CLK, Q => 
                           n33120, QN => n452);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7725, CK => CLK, Q => 
                           n33121, QN => n453);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7726, CK => CLK, Q => 
                           n33122, QN => n454);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7663, CK => CLK, Q => 
                           n32991, QN => n391);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7664, CK => CLK, Q => 
                           n32992, QN => n392);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7665, CK => CLK, Q => 
                           n32993, QN => n393);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7666, CK => CLK, Q => 
                           n32994, QN => n394);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7667, CK => CLK, Q => 
                           n32995, QN => n395);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7668, CK => CLK, Q => 
                           n32996, QN => n396);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7669, CK => CLK, Q => 
                           n32997, QN => n397);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7670, CK => CLK, Q => 
                           n32998, QN => n398);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7671, CK => CLK, Q => 
                           n32999, QN => n399);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7672, CK => CLK, Q => 
                           n33000, QN => n400);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7673, CK => CLK, Q => 
                           n33001, QN => n401);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7674, CK => CLK, Q => 
                           n33002, QN => n402);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7675, CK => CLK, Q => 
                           n33003, QN => n403);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7676, CK => CLK, Q => 
                           n33004, QN => n404);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7677, CK => CLK, Q => 
                           n33005, QN => n405);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7678, CK => CLK, Q => 
                           n33006, QN => n406);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7679, CK => CLK, Q => 
                           n33007, QN => n407);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7680, CK => CLK, Q => 
                           n33008, QN => n408);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7681, CK => CLK, Q => 
                           n33009, QN => n409);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7682, CK => CLK, Q => 
                           n33010, QN => n410);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7683, CK => CLK, Q => 
                           n33011, QN => n411);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7684, CK => CLK, Q => 
                           n33012, QN => n412);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7685, CK => CLK, Q => 
                           n33013, QN => n413);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7686, CK => CLK, Q => 
                           n33014, QN => n414);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7687, CK => CLK, Q => 
                           n33015, QN => n415);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7688, CK => CLK, Q => 
                           n33016, QN => n416);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7689, CK => CLK, Q => 
                           n33017, QN => n417);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7690, CK => CLK, Q => 
                           n33018, QN => n418);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7691, CK => CLK, Q => 
                           n33019, QN => n419);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7692, CK => CLK, Q => 
                           n33020, QN => n420);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7693, CK => CLK, Q => 
                           n33021, QN => n421);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7694, CK => CLK, Q => 
                           n33022, QN => n422);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7695, CK => CLK, Q => 
                           n33023, QN => n423);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7696, CK => CLK, Q => 
                           n33024, QN => n424);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7697, CK => CLK, Q => 
                           n33025, QN => n425);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7698, CK => CLK, Q => 
                           n33026, QN => n426);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7699, CK => CLK, Q => 
                           n33027, QN => n427);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7700, CK => CLK, Q => 
                           n33028, QN => n428);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7701, CK => CLK, Q => 
                           n33029, QN => n429);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7702, CK => CLK, Q => 
                           n33030, QN => n430);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7703, CK => CLK, Q => 
                           n33031, QN => n431);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7704, CK => CLK, Q => 
                           n33032, QN => n432);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7705, CK => CLK, Q => n33033
                           , QN => n433);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7706, CK => CLK, Q => n33034
                           , QN => n434);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7707, CK => CLK, Q => n33035
                           , QN => n435);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7708, CK => CLK, Q => n33036
                           , QN => n436);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7709, CK => CLK, Q => n33037
                           , QN => n437);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7710, CK => CLK, Q => n33038
                           , QN => n438);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7651, CK => CLK, Q => 
                           n33123, QN => n379);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7652, CK => CLK, Q => 
                           n33124, QN => n380);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7653, CK => CLK, Q => 
                           n33125, QN => n381);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7654, CK => CLK, Q => 
                           n33126, QN => n382);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7655, CK => CLK, Q => 
                           n33127, QN => n383);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7656, CK => CLK, Q => 
                           n33128, QN => n384);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7657, CK => CLK, Q => 
                           n33129, QN => n385);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7658, CK => CLK, Q => 
                           n33130, QN => n386);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7659, CK => CLK, Q => 
                           n33131, QN => n387);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7660, CK => CLK, Q => 
                           n33132, QN => n388);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7661, CK => CLK, Q => 
                           n33133, QN => n389);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7662, CK => CLK, Q => 
                           n33134, QN => n390);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n8357, CK => CLK, Q => 
                           n31123, QN => n25509);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n8355, CK => CLK, Q => 
                           n31121, QN => n25511);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n8356, CK => CLK, Q => 
                           n31122, QN => n25510);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n8358, CK => CLK, Q => 
                           n31124, QN => n25508);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n8359, CK => CLK, Q => 
                           n31125, QN => n25507);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n8360, CK => CLK, Q => 
                           n31126, QN => n25506);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n8361, CK => CLK, Q => 
                           n31127, QN => n25505);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n8362, CK => CLK, Q => 
                           n31128, QN => n25504);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n8363, CK => CLK, Q => 
                           n31129, QN => n25503);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n8364, CK => CLK, Q => 
                           n31130, QN => n25502);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n8365, CK => CLK, Q => 
                           n31131, QN => n25501);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n8366, CK => CLK, Q => 
                           n31132, QN => n25500);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n8367, CK => CLK, Q => 
                           n31133, QN => n25499);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n8368, CK => CLK, Q => 
                           n31134, QN => n25498);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n8369, CK => CLK, Q => 
                           n31135, QN => n25497);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n8370, CK => CLK, Q => 
                           n31136, QN => n25496);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n8371, CK => CLK, Q => 
                           n31137, QN => n25495);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n8372, CK => CLK, Q => 
                           n31138, QN => n25494);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n8373, CK => CLK, Q => 
                           n31139, QN => n25493);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n8374, CK => CLK, Q => 
                           n31140, QN => n25492);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n8375, CK => CLK, Q => 
                           n31141, QN => n25491);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n8376, CK => CLK, Q => 
                           n31142, QN => n25490);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n8377, CK => CLK, Q => 
                           n31143, QN => n25489);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n8378, CK => CLK, Q => 
                           n31144, QN => n25488);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n8379, CK => CLK, Q => 
                           n31145, QN => n25487);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n8380, CK => CLK, Q => 
                           n31146, QN => n25486);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n8381, CK => CLK, Q => 
                           n31147, QN => n25485);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n8382, CK => CLK, Q => 
                           n31148, QN => n25484);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n8383, CK => CLK, Q => 
                           n31149, QN => n25483);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n8384, CK => CLK, Q => 
                           n31150, QN => n25482);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n8385, CK => CLK, Q => 
                           n31151, QN => n25481);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n8386, CK => CLK, Q => 
                           n31152, QN => n25480);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n8387, CK => CLK, Q => 
                           n31153, QN => n25479);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n8388, CK => CLK, Q => 
                           n31154, QN => n25478);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n8389, CK => CLK, Q => 
                           n31155, QN => n25477);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n8390, CK => CLK, Q => 
                           n31156, QN => n25476);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n8391, CK => CLK, Q => 
                           n31157, QN => n25475);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n8392, CK => CLK, Q => 
                           n31158, QN => n25474);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n8393, CK => CLK, Q => 
                           n31159, QN => n25473);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n8394, CK => CLK, Q => 
                           n31160, QN => n25472);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n8395, CK => CLK, Q => 
                           n31161, QN => n25471);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n8396, CK => CLK, Q => 
                           n31162, QN => n25470);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n8397, CK => CLK, Q => 
                           n31163, QN => n25469);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n8398, CK => CLK, Q => 
                           n31164, QN => n25468);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n8399, CK => CLK, Q => 
                           n31165, QN => n25467);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n8400, CK => CLK, Q => 
                           n31166, QN => n25466);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n8401, CK => CLK, Q => 
                           n31167, QN => n25465);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n8402, CK => CLK, Q => 
                           n31168, QN => n25464);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n8403, CK => CLK, Q => 
                           n31169, QN => n25463);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n8404, CK => CLK, Q => 
                           n31170, QN => n25462);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n8405, CK => CLK, Q => 
                           n31171, QN => n25461);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n8406, CK => CLK, Q => 
                           n31172, QN => n25460);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n8407, CK => CLK, Q => 
                           n31173, QN => n25459);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n8408, CK => CLK, Q => 
                           n31174, QN => n25458);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n32518, QN => n71);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n32519, QN => n72);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n32520, QN => n73);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n32521, QN => n74);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n32522, QN => n75);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n32523, QN => n76);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n32524, QN => n77);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n32525, QN => n78);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n32526, QN => n79);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n32527, QN => n80);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n32528, QN => n81);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n32529, QN => n82);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n32530, QN => n83);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n32531, QN => n84);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => 
                           n32532, QN => n85);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => 
                           n32533, QN => n86);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => 
                           n32534, QN => n87);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => 
                           n32535, QN => n88);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => 
                           n32536, QN => n89);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => 
                           n32537, QN => n90);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => 
                           n32538, QN => n91);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => 
                           n32539, QN => n92);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => 
                           n32540, QN => n93);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => 
                           n32541, QN => n94);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => 
                           n32542, QN => n95);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => 
                           n32543, QN => n96);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => 
                           n32544, QN => n97);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => 
                           n32545, QN => n98);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => 
                           n32546, QN => n99);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => 
                           n30458, QN => n27921);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => 
                           n30459, QN => n27922);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => 
                           n30460, QN => n27923);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => 
                           n30461, QN => n27924);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => 
                           n30462, QN => n27925);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => 
                           n30463, QN => n27926);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => 
                           n30464, QN => n27927);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n30465, QN => n27928);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n30466, QN => n27929);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n30467, QN => n27930);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n30468, QN => n27931);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n30469, QN => n27932);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n30470, QN => n27933);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => n30471
                           , QN => n27934);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => n30472
                           , QN => n27935);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => n30473
                           , QN => n27936);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => n30474
                           , QN => n27937);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => n30475
                           , QN => n27938);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => n30476
                           , QN => n27939);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n32508, QN => n59);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n32509, QN => n60);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n32506, QN => n61);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n32507, QN => n62);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n32510, QN => n63);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n32511, QN => n64);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n32512, QN => n65);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n32513, QN => n66);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n32514, QN => n67);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n32515, QN => n68);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n32516, QN => n69);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n32517, QN => n70);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n8047, CK => CLK, Q => 
                           n32727, QN => n775);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n8048, CK => CLK, Q => 
                           n32728, QN => n776);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n8049, CK => CLK, Q => 
                           n32729, QN => n777);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n8050, CK => CLK, Q => 
                           n32730, QN => n778);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n8051, CK => CLK, Q => 
                           n32731, QN => n779);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n8052, CK => CLK, Q => 
                           n32732, QN => n780);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n8053, CK => CLK, Q => 
                           n32733, QN => n781);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n8054, CK => CLK, Q => 
                           n32734, QN => n782);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n8055, CK => CLK, Q => 
                           n32735, QN => n783);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n8056, CK => CLK, Q => 
                           n32736, QN => n784);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n8057, CK => CLK, Q => 
                           n32737, QN => n785);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n8058, CK => CLK, Q => 
                           n32738, QN => n786);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n8059, CK => CLK, Q => 
                           n32739, QN => n787);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n8060, CK => CLK, Q => 
                           n32740, QN => n788);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n8061, CK => CLK, Q => 
                           n32741, QN => n789);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n8062, CK => CLK, Q => 
                           n32742, QN => n790);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n8063, CK => CLK, Q => 
                           n32743, QN => n791);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n8064, CK => CLK, Q => 
                           n32744, QN => n792);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n8065, CK => CLK, Q => 
                           n32745, QN => n793);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n8066, CK => CLK, Q => 
                           n32746, QN => n794);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n8067, CK => CLK, Q => 
                           n32747, QN => n795);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n8068, CK => CLK, Q => 
                           n32748, QN => n796);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n8069, CK => CLK, Q => 
                           n32749, QN => n797);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n8070, CK => CLK, Q => 
                           n32750, QN => n798);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n8071, CK => CLK, Q => 
                           n32751, QN => n799);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n8072, CK => CLK, Q => 
                           n32752, QN => n800);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n8073, CK => CLK, Q => 
                           n32753, QN => n801);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n8074, CK => CLK, Q => 
                           n32754, QN => n802);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n8075, CK => CLK, Q => 
                           n32755, QN => n803);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n8076, CK => CLK, Q => 
                           n32756, QN => n804);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n8077, CK => CLK, Q => 
                           n32757, QN => n805);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n8078, CK => CLK, Q => 
                           n32758, QN => n806);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n8079, CK => CLK, Q => 
                           n32759, QN => n807);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n8080, CK => CLK, Q => 
                           n32760, QN => n808);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n8081, CK => CLK, Q => 
                           n32761, QN => n809);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n8082, CK => CLK, Q => 
                           n32762, QN => n810);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n8083, CK => CLK, Q => 
                           n32763, QN => n811_port);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n8084, CK => CLK, Q => 
                           n32764, QN => n812_port);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n8085, CK => CLK, Q => 
                           n32765, QN => n813_port);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n8086, CK => CLK, Q => 
                           n32766, QN => n814);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n8087, CK => CLK, Q => 
                           n32767, QN => n815);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n8088, CK => CLK, Q => 
                           n32768, QN => n816);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n8089, CK => CLK, Q => 
                           n32769, QN => n817);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n8090, CK => CLK, Q => 
                           n32770, QN => n818);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n8091, CK => CLK, Q => 
                           n32771, QN => n819);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n8092, CK => CLK, Q => 
                           n32772, QN => n820);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n8093, CK => CLK, Q => 
                           n32773, QN => n821);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n8094, CK => CLK, Q => 
                           n32774, QN => n822);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n7983, CK => CLK, Q => 
                           n32775, QN => n711);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n7984, CK => CLK, Q => 
                           n32776, QN => n712);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n7985, CK => CLK, Q => 
                           n32777, QN => n713);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n7986, CK => CLK, Q => 
                           n32778, QN => n714);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n7987, CK => CLK, Q => 
                           n32779, QN => n715);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n7988, CK => CLK, Q => 
                           n32780, QN => n716);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n7989, CK => CLK, Q => 
                           n32781, QN => n717);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n7990, CK => CLK, Q => 
                           n32782, QN => n718);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n7991, CK => CLK, Q => 
                           n32783, QN => n719);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n7992, CK => CLK, Q => 
                           n32784, QN => n720);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n7993, CK => CLK, Q => 
                           n32785, QN => n721);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n7994, CK => CLK, Q => 
                           n32786, QN => n722);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n7995, CK => CLK, Q => 
                           n32787, QN => n723);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n7996, CK => CLK, Q => 
                           n32788, QN => n724);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n7997, CK => CLK, Q => 
                           n32789, QN => n725);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n7998, CK => CLK, Q => 
                           n32790, QN => n726);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n7999, CK => CLK, Q => 
                           n32791, QN => n727);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n8000, CK => CLK, Q => 
                           n32792, QN => n728);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n8001, CK => CLK, Q => 
                           n32793, QN => n729);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n8002, CK => CLK, Q => 
                           n32794, QN => n730);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n8003, CK => CLK, Q => 
                           n32795, QN => n731);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n8004, CK => CLK, Q => 
                           n32796, QN => n732);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n8005, CK => CLK, Q => 
                           n32797, QN => n733);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n8006, CK => CLK, Q => 
                           n32798, QN => n734);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n8007, CK => CLK, Q => 
                           n32799, QN => n735);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n8008, CK => CLK, Q => 
                           n32800, QN => n736);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n8009, CK => CLK, Q => 
                           n32801, QN => n737);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n8010, CK => CLK, Q => 
                           n32802, QN => n738);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n8011, CK => CLK, Q => 
                           n32803, QN => n739);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n8012, CK => CLK, Q => 
                           n32804, QN => n740);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n8013, CK => CLK, Q => 
                           n32805, QN => n741);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n8014, CK => CLK, Q => 
                           n32806, QN => n742);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n8015, CK => CLK, Q => 
                           n32807, QN => n743);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n8016, CK => CLK, Q => 
                           n32808, QN => n744);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n8017, CK => CLK, Q => 
                           n32809, QN => n745);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n8018, CK => CLK, Q => 
                           n32810, QN => n746);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n8019, CK => CLK, Q => 
                           n32811, QN => n747);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n8020, CK => CLK, Q => 
                           n32812, QN => n748);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n8021, CK => CLK, Q => 
                           n32813, QN => n749);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n8022, CK => CLK, Q => 
                           n32814, QN => n750);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n8023, CK => CLK, Q => 
                           n32815, QN => n751);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n8024, CK => CLK, Q => 
                           n32816, QN => n752);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n8025, CK => CLK, Q => 
                           n32817, QN => n753);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n8026, CK => CLK, Q => 
                           n32818, QN => n754);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n8027, CK => CLK, Q => 
                           n32819, QN => n755);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n8028, CK => CLK, Q => 
                           n32820, QN => n756);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n8029, CK => CLK, Q => 
                           n32821, QN => n757);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n8030, CK => CLK, Q => 
                           n32822, QN => n758);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n8035, CK => CLK, Q => 
                           n32823, QN => n763);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n8036, CK => CLK, Q => 
                           n32824, QN => n764);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n8037, CK => CLK, Q => 
                           n32825, QN => n765);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n8038, CK => CLK, Q => 
                           n32826, QN => n766);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n8039, CK => CLK, Q => 
                           n32827, QN => n767);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n8040, CK => CLK, Q => 
                           n32828, QN => n768);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n8041, CK => CLK, Q => 
                           n32829, QN => n769);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n8042, CK => CLK, Q => 
                           n32830, QN => n770);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n8043, CK => CLK, Q => 
                           n32831, QN => n771);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n8044, CK => CLK, Q => 
                           n32832, QN => n772);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n8045, CK => CLK, Q => 
                           n32833, QN => n773);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n8046, CK => CLK, Q => 
                           n32834, QN => n774);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n7971, CK => CLK, Q => 
                           n32835, QN => n699);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n7972, CK => CLK, Q => 
                           n32836, QN => n700);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n7973, CK => CLK, Q => 
                           n32837, QN => n701);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n7974, CK => CLK, Q => 
                           n32838, QN => n702);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n7975, CK => CLK, Q => 
                           n32839, QN => n703);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n7976, CK => CLK, Q => 
                           n32840, QN => n704);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n7977, CK => CLK, Q => 
                           n32841, QN => n705);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n7978, CK => CLK, Q => 
                           n32842, QN => n706);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n7979, CK => CLK, Q => 
                           n32843, QN => n707);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n7980, CK => CLK, Q => 
                           n32844, QN => n708);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n7981, CK => CLK, Q => 
                           n32845, QN => n709);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n7982, CK => CLK, Q => 
                           n32846, QN => n710);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n8303, CK => CLK, Q => 
                           n31069, QN => n25449);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n8304, CK => CLK, Q => 
                           n31070, QN => n25448);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n8305, CK => CLK, Q => 
                           n31071, QN => n25447);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n8306, CK => CLK, Q => 
                           n31072, QN => n25446);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n8307, CK => CLK, Q => 
                           n31073, QN => n25445);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n8308, CK => CLK, Q => 
                           n31074, QN => n25444);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n8309, CK => CLK, Q => 
                           n31075, QN => n25443);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n8310, CK => CLK, Q => 
                           n31076, QN => n25442);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n8311, CK => CLK, Q => 
                           n31077, QN => n25441);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n8312, CK => CLK, Q => 
                           n31078, QN => n25440);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n8313, CK => CLK, Q => 
                           n31079, QN => n25439);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n8314, CK => CLK, Q => 
                           n31080, QN => n25438);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n8315, CK => CLK, Q => 
                           n31081, QN => n25437);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n8316, CK => CLK, Q => 
                           n31082, QN => n25436);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n8317, CK => CLK, Q => 
                           n31083, QN => n25435);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n8318, CK => CLK, Q => 
                           n31084, QN => n25434);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n8319, CK => CLK, Q => 
                           n31085, QN => n25433);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n8320, CK => CLK, Q => 
                           n31086, QN => n25432);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n8321, CK => CLK, Q => 
                           n31087, QN => n25431);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n8322, CK => CLK, Q => 
                           n31088, QN => n25430);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n8323, CK => CLK, Q => 
                           n31089, QN => n25429);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n8324, CK => CLK, Q => 
                           n31090, QN => n25428);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n8325, CK => CLK, Q => 
                           n31091, QN => n25427);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n8326, CK => CLK, Q => 
                           n31092, QN => n25426);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n8327, CK => CLK, Q => 
                           n31093, QN => n25425);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n8328, CK => CLK, Q => 
                           n31094, QN => n25424);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n8329, CK => CLK, Q => 
                           n31095, QN => n25423);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n8330, CK => CLK, Q => 
                           n31096, QN => n25422);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n8331, CK => CLK, Q => 
                           n31097, QN => n25421);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n8332, CK => CLK, Q => 
                           n31098, QN => n25420);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n8333, CK => CLK, Q => 
                           n31099, QN => n25419);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n8334, CK => CLK, Q => 
                           n31100, QN => n25418);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n8335, CK => CLK, Q => 
                           n31101, QN => n25417);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n8336, CK => CLK, Q => 
                           n31102, QN => n25416);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n8337, CK => CLK, Q => 
                           n31103, QN => n25415);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n8338, CK => CLK, Q => 
                           n31104, QN => n25414);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n8339, CK => CLK, Q => 
                           n31105, QN => n25413);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n8340, CK => CLK, Q => 
                           n31106, QN => n25412);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n8341, CK => CLK, Q => 
                           n31107, QN => n25411);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n8342, CK => CLK, Q => 
                           n31108, QN => n25410);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n8343, CK => CLK, Q => 
                           n31109, QN => n25409);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n8344, CK => CLK, Q => 
                           n31110, QN => n25408);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n8345, CK => CLK, Q => 
                           n31111, QN => n25407);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n8346, CK => CLK, Q => 
                           n31112, QN => n25406);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n8347, CK => CLK, Q => 
                           n31113, QN => n25405);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n8348, CK => CLK, Q => 
                           n31114, QN => n25404);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n8349, CK => CLK, Q => 
                           n31115, QN => n25403);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n8350, CK => CLK, Q => 
                           n31116, QN => n25402);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n8291, CK => CLK, Q => 
                           n31057, QN => n25397);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n8292, CK => CLK, Q => 
                           n31058, QN => n25396);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n8293, CK => CLK, Q => 
                           n31059, QN => n25395);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n8294, CK => CLK, Q => 
                           n31060, QN => n25457);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n8295, CK => CLK, Q => 
                           n31061, QN => n28840);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n8296, CK => CLK, Q => 
                           n31062, QN => n25456);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n8297, CK => CLK, Q => 
                           n31063, QN => n25455);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n8298, CK => CLK, Q => 
                           n31064, QN => n25454);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n8299, CK => CLK, Q => 
                           n31065, QN => n25453);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n8300, CK => CLK, Q => 
                           n31066, QN => n25452);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n8301, CK => CLK, Q => 
                           n31067, QN => n25451);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n8302, CK => CLK, Q => 
                           n31068, QN => n25450);
   U26462 : NOR3_X1 port map( A1 => n32243, A2 => N690, A3 => n37226, ZN => 
                           n37249);
   U26463 : NOR3_X1 port map( A1 => N6272, A2 => N6273, A3 => n34672, ZN => 
                           n34693);
   U26464 : NOR3_X1 port map( A1 => N6397, A2 => N6398, A3 => n35946, ZN => 
                           n35967);
   U26465 : XNOR2_X1 port map( A => n37251, B => n32244, ZN => n37226);
   U26466 : XNOR2_X1 port map( A => n34697, B => r504_carry_5_port, ZN => 
                           n34672);
   U26467 : XNOR2_X1 port map( A => n35971, B => r510_carry_5_port, ZN => 
                           n35946);
   U26468 : XNOR2_X1 port map( A => n32255, B => n2699, ZN => n33398);
   U26469 : BUF_X1 port map( A => n36016, Z => n39163);
   U26470 : BUF_X1 port map( A => n36016, Z => n39164);
   U26471 : BUF_X1 port map( A => n36016, Z => n39165);
   U26472 : BUF_X1 port map( A => n36016, Z => n39162);
   U26473 : BUF_X1 port map( A => n36016, Z => n39166);
   U26474 : BUF_X1 port map( A => n39913, Z => n39914);
   U26475 : BUF_X1 port map( A => n39932, Z => n39933);
   U26476 : BUF_X1 port map( A => n39913, Z => n39918);
   U26477 : BUF_X1 port map( A => n39913, Z => n39917);
   U26478 : BUF_X1 port map( A => n39913, Z => n39916);
   U26479 : BUF_X1 port map( A => n39913, Z => n39915);
   U26480 : BUF_X1 port map( A => n39932, Z => n39937);
   U26481 : BUF_X1 port map( A => n39932, Z => n39936);
   U26482 : BUF_X1 port map( A => n39932, Z => n39935);
   U26483 : BUF_X1 port map( A => n39932, Z => n39934);
   U26484 : BUF_X1 port map( A => n39952, Z => n39957);
   U26485 : BUF_X1 port map( A => n39952, Z => n39956);
   U26486 : BUF_X1 port map( A => n39952, Z => n39955);
   U26487 : BUF_X1 port map( A => n39952, Z => n39954);
   U26488 : BUF_X1 port map( A => n39952, Z => n39953);
   U26489 : BUF_X1 port map( A => n39894, Z => n39899);
   U26490 : BUF_X1 port map( A => n39894, Z => n39898);
   U26491 : BUF_X1 port map( A => n39894, Z => n39897);
   U26492 : BUF_X1 port map( A => n39894, Z => n39896);
   U26493 : BUF_X1 port map( A => n39894, Z => n39895);
   U26494 : BUF_X1 port map( A => n36028, Z => n39103);
   U26495 : BUF_X1 port map( A => n36034, Z => n39073);
   U26496 : BUF_X1 port map( A => n36028, Z => n39104);
   U26497 : BUF_X1 port map( A => n36034, Z => n39074);
   U26498 : BUF_X1 port map( A => n36028, Z => n39105);
   U26499 : BUF_X1 port map( A => n36034, Z => n39075);
   U26500 : BUF_X1 port map( A => n36028, Z => n39102);
   U26501 : BUF_X1 port map( A => n36034, Z => n39072);
   U26502 : BUF_X1 port map( A => n36028, Z => n39106);
   U26503 : BUF_X1 port map( A => n36034, Z => n39076);
   U26504 : BUF_X1 port map( A => n33473, Z => n39608);
   U26505 : BUF_X1 port map( A => n33479, Z => n39578);
   U26506 : BUF_X1 port map( A => n34747, Z => n39356);
   U26507 : BUF_X1 port map( A => n34753, Z => n39326);
   U26508 : BUF_X1 port map( A => n33473, Z => n39607);
   U26509 : BUF_X1 port map( A => n33479, Z => n39577);
   U26510 : BUF_X1 port map( A => n34747, Z => n39355);
   U26511 : BUF_X1 port map( A => n34753, Z => n39325);
   U26512 : BUF_X1 port map( A => n33473, Z => n39606);
   U26513 : BUF_X1 port map( A => n33479, Z => n39576);
   U26514 : BUF_X1 port map( A => n34747, Z => n39354);
   U26515 : BUF_X1 port map( A => n34753, Z => n39324);
   U26516 : BUF_X1 port map( A => n33473, Z => n39605);
   U26517 : BUF_X1 port map( A => n33479, Z => n39575);
   U26518 : BUF_X1 port map( A => n34747, Z => n39353);
   U26519 : BUF_X1 port map( A => n34753, Z => n39323);
   U26520 : BUF_X1 port map( A => n33473, Z => n39604);
   U26521 : BUF_X1 port map( A => n33479, Z => n39574);
   U26522 : BUF_X1 port map( A => n34747, Z => n39352);
   U26523 : BUF_X1 port map( A => n34753, Z => n39322);
   U26524 : BUF_X1 port map( A => n36022, Z => n39133);
   U26525 : BUF_X1 port map( A => n36006, Z => n39193);
   U26526 : BUF_X1 port map( A => n36000, Z => n39223);
   U26527 : BUF_X1 port map( A => n35988, Z => n39283);
   U26528 : BUF_X1 port map( A => n35994, Z => n39253);
   U26529 : BUF_X1 port map( A => n36022, Z => n39134);
   U26530 : BUF_X1 port map( A => n36006, Z => n39194);
   U26531 : BUF_X1 port map( A => n36000, Z => n39224);
   U26532 : BUF_X1 port map( A => n35988, Z => n39284);
   U26533 : BUF_X1 port map( A => n35994, Z => n39254);
   U26534 : BUF_X1 port map( A => n36022, Z => n39135);
   U26535 : BUF_X1 port map( A => n36006, Z => n39195);
   U26536 : BUF_X1 port map( A => n36000, Z => n39225);
   U26537 : BUF_X1 port map( A => n35988, Z => n39285);
   U26538 : BUF_X1 port map( A => n35994, Z => n39255);
   U26539 : BUF_X1 port map( A => n36022, Z => n39132);
   U26540 : BUF_X1 port map( A => n36006, Z => n39192);
   U26541 : BUF_X1 port map( A => n36000, Z => n39222);
   U26542 : BUF_X1 port map( A => n35988, Z => n39282);
   U26543 : BUF_X1 port map( A => n35994, Z => n39252);
   U26544 : BUF_X1 port map( A => n36022, Z => n39136);
   U26545 : BUF_X1 port map( A => n36006, Z => n39196);
   U26546 : BUF_X1 port map( A => n36000, Z => n39226);
   U26547 : BUF_X1 port map( A => n35988, Z => n39286);
   U26548 : BUF_X1 port map( A => n35994, Z => n39256);
   U26549 : BUF_X1 port map( A => n33467, Z => n39638);
   U26550 : BUF_X1 port map( A => n33461, Z => n39668);
   U26551 : BUF_X1 port map( A => n33433, Z => n39788);
   U26552 : BUF_X1 port map( A => n33439, Z => n39758);
   U26553 : BUF_X1 port map( A => n33445, Z => n39728);
   U26554 : BUF_X1 port map( A => n33451, Z => n39698);
   U26555 : BUF_X1 port map( A => n34741, Z => n39386);
   U26556 : BUF_X1 port map( A => n34735, Z => n39416);
   U26557 : BUF_X1 port map( A => n34707, Z => n39536);
   U26558 : BUF_X1 port map( A => n34713, Z => n39506);
   U26559 : BUF_X1 port map( A => n34719, Z => n39476);
   U26560 : BUF_X1 port map( A => n34725, Z => n39446);
   U26561 : BUF_X1 port map( A => n33467, Z => n39637);
   U26562 : BUF_X1 port map( A => n33461, Z => n39667);
   U26563 : BUF_X1 port map( A => n33433, Z => n39787);
   U26564 : BUF_X1 port map( A => n33439, Z => n39757);
   U26565 : BUF_X1 port map( A => n33445, Z => n39727);
   U26566 : BUF_X1 port map( A => n33451, Z => n39697);
   U26567 : BUF_X1 port map( A => n34741, Z => n39385);
   U26568 : BUF_X1 port map( A => n34735, Z => n39415);
   U26569 : BUF_X1 port map( A => n34707, Z => n39535);
   U26570 : BUF_X1 port map( A => n34713, Z => n39505);
   U26571 : BUF_X1 port map( A => n34719, Z => n39475);
   U26572 : BUF_X1 port map( A => n34725, Z => n39445);
   U26573 : BUF_X1 port map( A => n33467, Z => n39636);
   U26574 : BUF_X1 port map( A => n33461, Z => n39666);
   U26575 : BUF_X1 port map( A => n33433, Z => n39786);
   U26576 : BUF_X1 port map( A => n33439, Z => n39756);
   U26577 : BUF_X1 port map( A => n33445, Z => n39726);
   U26578 : BUF_X1 port map( A => n33451, Z => n39696);
   U26579 : BUF_X1 port map( A => n34741, Z => n39384);
   U26580 : BUF_X1 port map( A => n34735, Z => n39414);
   U26581 : BUF_X1 port map( A => n34707, Z => n39534);
   U26582 : BUF_X1 port map( A => n34713, Z => n39504);
   U26583 : BUF_X1 port map( A => n34719, Z => n39474);
   U26584 : BUF_X1 port map( A => n34725, Z => n39444);
   U26585 : BUF_X1 port map( A => n33467, Z => n39635);
   U26586 : BUF_X1 port map( A => n33461, Z => n39665);
   U26587 : BUF_X1 port map( A => n33433, Z => n39785);
   U26588 : BUF_X1 port map( A => n33439, Z => n39755);
   U26589 : BUF_X1 port map( A => n33445, Z => n39725);
   U26590 : BUF_X1 port map( A => n33451, Z => n39695);
   U26591 : BUF_X1 port map( A => n34741, Z => n39383);
   U26592 : BUF_X1 port map( A => n34735, Z => n39413);
   U26593 : BUF_X1 port map( A => n34707, Z => n39533);
   U26594 : BUF_X1 port map( A => n34713, Z => n39503);
   U26595 : BUF_X1 port map( A => n34719, Z => n39473);
   U26596 : BUF_X1 port map( A => n34725, Z => n39443);
   U26597 : BUF_X1 port map( A => n33467, Z => n39634);
   U26598 : BUF_X1 port map( A => n33461, Z => n39664);
   U26599 : BUF_X1 port map( A => n33433, Z => n39784);
   U26600 : BUF_X1 port map( A => n33439, Z => n39754);
   U26601 : BUF_X1 port map( A => n33445, Z => n39724);
   U26602 : BUF_X1 port map( A => n33451, Z => n39694);
   U26603 : BUF_X1 port map( A => n34741, Z => n39382);
   U26604 : BUF_X1 port map( A => n34735, Z => n39412);
   U26605 : BUF_X1 port map( A => n34707, Z => n39532);
   U26606 : BUF_X1 port map( A => n34713, Z => n39502);
   U26607 : BUF_X1 port map( A => n34719, Z => n39472);
   U26608 : BUF_X1 port map( A => n34725, Z => n39442);
   U26609 : BUF_X1 port map( A => n36029, Z => n39097);
   U26610 : BUF_X1 port map( A => n36035, Z => n39067);
   U26611 : BUF_X1 port map( A => n36029, Z => n39098);
   U26612 : BUF_X1 port map( A => n36035, Z => n39068);
   U26613 : BUF_X1 port map( A => n36029, Z => n39099);
   U26614 : BUF_X1 port map( A => n36035, Z => n39069);
   U26615 : BUF_X1 port map( A => n36029, Z => n39096);
   U26616 : BUF_X1 port map( A => n36035, Z => n39066);
   U26617 : BUF_X1 port map( A => n36029, Z => n39100);
   U26618 : BUF_X1 port map( A => n36035, Z => n39070);
   U26619 : BUF_X1 port map( A => n33474, Z => n39602);
   U26620 : BUF_X1 port map( A => n33480, Z => n39572);
   U26621 : BUF_X1 port map( A => n34748, Z => n39350);
   U26622 : BUF_X1 port map( A => n34754, Z => n39320);
   U26623 : BUF_X1 port map( A => n33474, Z => n39601);
   U26624 : BUF_X1 port map( A => n33480, Z => n39571);
   U26625 : BUF_X1 port map( A => n34748, Z => n39349);
   U26626 : BUF_X1 port map( A => n34754, Z => n39319);
   U26627 : BUF_X1 port map( A => n33474, Z => n39600);
   U26628 : BUF_X1 port map( A => n33480, Z => n39570);
   U26629 : BUF_X1 port map( A => n34748, Z => n39348);
   U26630 : BUF_X1 port map( A => n34754, Z => n39318);
   U26631 : BUF_X1 port map( A => n33474, Z => n39599);
   U26632 : BUF_X1 port map( A => n33480, Z => n39569);
   U26633 : BUF_X1 port map( A => n34748, Z => n39347);
   U26634 : BUF_X1 port map( A => n34754, Z => n39317);
   U26635 : BUF_X1 port map( A => n33474, Z => n39598);
   U26636 : BUF_X1 port map( A => n33480, Z => n39568);
   U26637 : BUF_X1 port map( A => n34748, Z => n39346);
   U26638 : BUF_X1 port map( A => n34754, Z => n39316);
   U26639 : BUF_X1 port map( A => n36023, Z => n39127);
   U26640 : BUF_X1 port map( A => n36017, Z => n39157);
   U26641 : BUF_X1 port map( A => n36007, Z => n39187);
   U26642 : BUF_X1 port map( A => n36001, Z => n39217);
   U26643 : BUF_X1 port map( A => n35989, Z => n39277);
   U26644 : BUF_X1 port map( A => n35995, Z => n39247);
   U26645 : BUF_X1 port map( A => n36023, Z => n39128);
   U26646 : BUF_X1 port map( A => n36017, Z => n39158);
   U26647 : BUF_X1 port map( A => n36007, Z => n39188);
   U26648 : BUF_X1 port map( A => n36001, Z => n39218);
   U26649 : BUF_X1 port map( A => n35989, Z => n39278);
   U26650 : BUF_X1 port map( A => n35995, Z => n39248);
   U26651 : BUF_X1 port map( A => n36023, Z => n39129);
   U26652 : BUF_X1 port map( A => n36017, Z => n39159);
   U26653 : BUF_X1 port map( A => n36007, Z => n39189);
   U26654 : BUF_X1 port map( A => n36001, Z => n39219);
   U26655 : BUF_X1 port map( A => n35989, Z => n39279);
   U26656 : BUF_X1 port map( A => n35995, Z => n39249);
   U26657 : BUF_X1 port map( A => n36023, Z => n39126);
   U26658 : BUF_X1 port map( A => n36017, Z => n39156);
   U26659 : BUF_X1 port map( A => n36007, Z => n39186);
   U26660 : BUF_X1 port map( A => n36001, Z => n39216);
   U26661 : BUF_X1 port map( A => n35989, Z => n39276);
   U26662 : BUF_X1 port map( A => n35995, Z => n39246);
   U26663 : BUF_X1 port map( A => n36023, Z => n39130);
   U26664 : BUF_X1 port map( A => n36017, Z => n39160);
   U26665 : BUF_X1 port map( A => n36007, Z => n39190);
   U26666 : BUF_X1 port map( A => n36001, Z => n39220);
   U26667 : BUF_X1 port map( A => n35989, Z => n39280);
   U26668 : BUF_X1 port map( A => n35995, Z => n39250);
   U26669 : BUF_X1 port map( A => n33468, Z => n39632);
   U26670 : BUF_X1 port map( A => n33462, Z => n39662);
   U26671 : BUF_X1 port map( A => n33434, Z => n39782);
   U26672 : BUF_X1 port map( A => n33440, Z => n39752);
   U26673 : BUF_X1 port map( A => n33446, Z => n39722);
   U26674 : BUF_X1 port map( A => n33452, Z => n39692);
   U26675 : BUF_X1 port map( A => n34742, Z => n39380);
   U26676 : BUF_X1 port map( A => n34736, Z => n39410);
   U26677 : BUF_X1 port map( A => n34708, Z => n39530);
   U26678 : BUF_X1 port map( A => n34714, Z => n39500);
   U26679 : BUF_X1 port map( A => n34720, Z => n39470);
   U26680 : BUF_X1 port map( A => n34726, Z => n39440);
   U26681 : BUF_X1 port map( A => n33468, Z => n39631);
   U26682 : BUF_X1 port map( A => n33462, Z => n39661);
   U26683 : BUF_X1 port map( A => n33434, Z => n39781);
   U26684 : BUF_X1 port map( A => n33440, Z => n39751);
   U26685 : BUF_X1 port map( A => n33446, Z => n39721);
   U26686 : BUF_X1 port map( A => n33452, Z => n39691);
   U26687 : BUF_X1 port map( A => n34742, Z => n39379);
   U26688 : BUF_X1 port map( A => n34736, Z => n39409);
   U26689 : BUF_X1 port map( A => n34708, Z => n39529);
   U26690 : BUF_X1 port map( A => n34714, Z => n39499);
   U26691 : BUF_X1 port map( A => n34720, Z => n39469);
   U26692 : BUF_X1 port map( A => n34726, Z => n39439);
   U26693 : BUF_X1 port map( A => n33468, Z => n39630);
   U26694 : BUF_X1 port map( A => n33462, Z => n39660);
   U26695 : BUF_X1 port map( A => n33434, Z => n39780);
   U26696 : BUF_X1 port map( A => n33440, Z => n39750);
   U26697 : BUF_X1 port map( A => n33446, Z => n39720);
   U26698 : BUF_X1 port map( A => n33452, Z => n39690);
   U26699 : BUF_X1 port map( A => n34742, Z => n39378);
   U26700 : BUF_X1 port map( A => n34736, Z => n39408);
   U26701 : BUF_X1 port map( A => n34708, Z => n39528);
   U26702 : BUF_X1 port map( A => n34714, Z => n39498);
   U26703 : BUF_X1 port map( A => n34720, Z => n39468);
   U26704 : BUF_X1 port map( A => n34726, Z => n39438);
   U26705 : BUF_X1 port map( A => n33468, Z => n39629);
   U26706 : BUF_X1 port map( A => n33462, Z => n39659);
   U26707 : BUF_X1 port map( A => n33434, Z => n39779);
   U26708 : BUF_X1 port map( A => n33440, Z => n39749);
   U26709 : BUF_X1 port map( A => n33446, Z => n39719);
   U26710 : BUF_X1 port map( A => n33452, Z => n39689);
   U26711 : BUF_X1 port map( A => n34742, Z => n39377);
   U26712 : BUF_X1 port map( A => n34736, Z => n39407);
   U26713 : BUF_X1 port map( A => n34708, Z => n39527);
   U26714 : BUF_X1 port map( A => n34714, Z => n39497);
   U26715 : BUF_X1 port map( A => n34720, Z => n39467);
   U26716 : BUF_X1 port map( A => n34726, Z => n39437);
   U26717 : BUF_X1 port map( A => n33468, Z => n39628);
   U26718 : BUF_X1 port map( A => n33462, Z => n39658);
   U26719 : BUF_X1 port map( A => n33434, Z => n39778);
   U26720 : BUF_X1 port map( A => n33440, Z => n39748);
   U26721 : BUF_X1 port map( A => n33446, Z => n39718);
   U26722 : BUF_X1 port map( A => n33452, Z => n39688);
   U26723 : BUF_X1 port map( A => n34742, Z => n39376);
   U26724 : BUF_X1 port map( A => n34736, Z => n39406);
   U26725 : BUF_X1 port map( A => n34708, Z => n39526);
   U26726 : BUF_X1 port map( A => n34714, Z => n39496);
   U26727 : BUF_X1 port map( A => n34720, Z => n39466);
   U26728 : BUF_X1 port map( A => n34726, Z => n39436);
   U26729 : BUF_X1 port map( A => n33438, Z => n39764);
   U26730 : BUF_X1 port map( A => n33444, Z => n39734);
   U26731 : BUF_X1 port map( A => n34712, Z => n39512);
   U26732 : BUF_X1 port map( A => n34718, Z => n39482);
   U26733 : BUF_X1 port map( A => n33438, Z => n39763);
   U26734 : BUF_X1 port map( A => n33444, Z => n39733);
   U26735 : BUF_X1 port map( A => n34712, Z => n39511);
   U26736 : BUF_X1 port map( A => n34718, Z => n39481);
   U26737 : BUF_X1 port map( A => n33438, Z => n39762);
   U26738 : BUF_X1 port map( A => n33444, Z => n39732);
   U26739 : BUF_X1 port map( A => n34712, Z => n39510);
   U26740 : BUF_X1 port map( A => n34718, Z => n39480);
   U26741 : BUF_X1 port map( A => n33438, Z => n39761);
   U26742 : BUF_X1 port map( A => n33444, Z => n39731);
   U26743 : BUF_X1 port map( A => n34712, Z => n39509);
   U26744 : BUF_X1 port map( A => n34718, Z => n39479);
   U26745 : BUF_X1 port map( A => n33438, Z => n39760);
   U26746 : BUF_X1 port map( A => n33444, Z => n39730);
   U26747 : BUF_X1 port map( A => n34712, Z => n39508);
   U26748 : BUF_X1 port map( A => n34718, Z => n39478);
   U26749 : BUF_X1 port map( A => n35993, Z => n39259);
   U26750 : BUF_X1 port map( A => n35999, Z => n39229);
   U26751 : BUF_X1 port map( A => n35993, Z => n39260);
   U26752 : BUF_X1 port map( A => n35999, Z => n39230);
   U26753 : BUF_X1 port map( A => n35993, Z => n39261);
   U26754 : BUF_X1 port map( A => n35999, Z => n39231);
   U26755 : BUF_X1 port map( A => n35993, Z => n39258);
   U26756 : BUF_X1 port map( A => n35999, Z => n39228);
   U26757 : BUF_X1 port map( A => n35993, Z => n39262);
   U26758 : BUF_X1 port map( A => n35999, Z => n39232);
   U26759 : BUF_X1 port map( A => n33478, Z => n39584);
   U26760 : BUF_X1 port map( A => n33450, Z => n39704);
   U26761 : BUF_X1 port map( A => n34752, Z => n39332);
   U26762 : BUF_X1 port map( A => n34724, Z => n39452);
   U26763 : BUF_X1 port map( A => n33478, Z => n39583);
   U26764 : BUF_X1 port map( A => n33450, Z => n39703);
   U26765 : BUF_X1 port map( A => n34752, Z => n39331);
   U26766 : BUF_X1 port map( A => n34724, Z => n39451);
   U26767 : BUF_X1 port map( A => n33478, Z => n39582);
   U26768 : BUF_X1 port map( A => n33450, Z => n39702);
   U26769 : BUF_X1 port map( A => n34752, Z => n39330);
   U26770 : BUF_X1 port map( A => n34724, Z => n39450);
   U26771 : BUF_X1 port map( A => n33478, Z => n39581);
   U26772 : BUF_X1 port map( A => n33450, Z => n39701);
   U26773 : BUF_X1 port map( A => n34752, Z => n39329);
   U26774 : BUF_X1 port map( A => n34724, Z => n39449);
   U26775 : BUF_X1 port map( A => n33478, Z => n39580);
   U26776 : BUF_X1 port map( A => n33450, Z => n39700);
   U26777 : BUF_X1 port map( A => n34752, Z => n39328);
   U26778 : BUF_X1 port map( A => n34724, Z => n39448);
   U26779 : BUF_X1 port map( A => n33484, Z => n39554);
   U26780 : BUF_X1 port map( A => n33484, Z => n39553);
   U26781 : BUF_X1 port map( A => n36033, Z => n39079);
   U26782 : BUF_X1 port map( A => n36039, Z => n39049);
   U26783 : BUF_X1 port map( A => n36021, Z => n39139);
   U26784 : BUF_X1 port map( A => n36011, Z => n39169);
   U26785 : BUF_X1 port map( A => n36033, Z => n39080);
   U26786 : BUF_X1 port map( A => n36039, Z => n39050);
   U26787 : BUF_X1 port map( A => n36021, Z => n39140);
   U26788 : BUF_X1 port map( A => n36011, Z => n39170);
   U26789 : BUF_X1 port map( A => n36033, Z => n39081);
   U26790 : BUF_X1 port map( A => n36039, Z => n39051);
   U26791 : BUF_X1 port map( A => n36021, Z => n39141);
   U26792 : BUF_X1 port map( A => n36011, Z => n39171);
   U26793 : BUF_X1 port map( A => n36033, Z => n39078);
   U26794 : BUF_X1 port map( A => n36039, Z => n39048);
   U26795 : BUF_X1 port map( A => n36021, Z => n39138);
   U26796 : BUF_X1 port map( A => n36011, Z => n39168);
   U26797 : BUF_X1 port map( A => n36033, Z => n39082);
   U26798 : BUF_X1 port map( A => n36039, Z => n39052);
   U26799 : BUF_X1 port map( A => n36021, Z => n39142);
   U26800 : BUF_X1 port map( A => n36011, Z => n39172);
   U26801 : BUF_X1 port map( A => n33466, Z => n39644);
   U26802 : BUF_X1 port map( A => n34758, Z => n39302);
   U26803 : BUF_X1 port map( A => n34740, Z => n39392);
   U26804 : BUF_X1 port map( A => n33466, Z => n39643);
   U26805 : BUF_X1 port map( A => n34758, Z => n39301);
   U26806 : BUF_X1 port map( A => n34740, Z => n39391);
   U26807 : BUF_X1 port map( A => n33484, Z => n39552);
   U26808 : BUF_X1 port map( A => n33466, Z => n39642);
   U26809 : BUF_X1 port map( A => n34758, Z => n39300);
   U26810 : BUF_X1 port map( A => n34740, Z => n39390);
   U26811 : BUF_X1 port map( A => n33484, Z => n39551);
   U26812 : BUF_X1 port map( A => n33466, Z => n39641);
   U26813 : BUF_X1 port map( A => n34758, Z => n39299);
   U26814 : BUF_X1 port map( A => n34740, Z => n39389);
   U26815 : BUF_X1 port map( A => n33484, Z => n39550);
   U26816 : BUF_X1 port map( A => n33466, Z => n39640);
   U26817 : BUF_X1 port map( A => n34758, Z => n39298);
   U26818 : BUF_X1 port map( A => n34740, Z => n39388);
   U26819 : BUF_X1 port map( A => n36005, Z => n39199);
   U26820 : BUF_X1 port map( A => n36005, Z => n39200);
   U26821 : BUF_X1 port map( A => n36005, Z => n39201);
   U26822 : BUF_X1 port map( A => n36005, Z => n39198);
   U26823 : BUF_X1 port map( A => n36005, Z => n39202);
   U26824 : BUF_X1 port map( A => n36027, Z => n39109);
   U26825 : BUF_X1 port map( A => n36027, Z => n39110);
   U26826 : BUF_X1 port map( A => n36027, Z => n39111);
   U26827 : BUF_X1 port map( A => n36027, Z => n39108);
   U26828 : BUF_X1 port map( A => n36027, Z => n39112);
   U26829 : BUF_X1 port map( A => n33472, Z => n39614);
   U26830 : BUF_X1 port map( A => n34746, Z => n39362);
   U26831 : BUF_X1 port map( A => n33472, Z => n39613);
   U26832 : BUF_X1 port map( A => n34746, Z => n39361);
   U26833 : BUF_X1 port map( A => n33472, Z => n39612);
   U26834 : BUF_X1 port map( A => n34746, Z => n39360);
   U26835 : BUF_X1 port map( A => n33472, Z => n39611);
   U26836 : BUF_X1 port map( A => n34746, Z => n39359);
   U26837 : BUF_X1 port map( A => n33472, Z => n39610);
   U26838 : BUF_X1 port map( A => n34746, Z => n39358);
   U26839 : BUF_X1 port map( A => n33456, Z => n39674);
   U26840 : BUF_X1 port map( A => n34730, Z => n39422);
   U26841 : BUF_X1 port map( A => n33456, Z => n39673);
   U26842 : BUF_X1 port map( A => n34730, Z => n39421);
   U26843 : BUF_X1 port map( A => n33456, Z => n39672);
   U26844 : BUF_X1 port map( A => n34730, Z => n39420);
   U26845 : BUF_X1 port map( A => n33456, Z => n39671);
   U26846 : BUF_X1 port map( A => n34730, Z => n39419);
   U26847 : BUF_X1 port map( A => n33456, Z => n39670);
   U26848 : BUF_X1 port map( A => n34730, Z => n39418);
   U26849 : BUF_X1 port map( A => n33436, Z => n39776);
   U26850 : BUF_X1 port map( A => n33442, Z => n39746);
   U26851 : BUF_X1 port map( A => n34710, Z => n39524);
   U26852 : BUF_X1 port map( A => n34716, Z => n39494);
   U26853 : BUF_X1 port map( A => n33436, Z => n39775);
   U26854 : BUF_X1 port map( A => n33442, Z => n39745);
   U26855 : BUF_X1 port map( A => n34710, Z => n39523);
   U26856 : BUF_X1 port map( A => n34716, Z => n39493);
   U26857 : BUF_X1 port map( A => n33436, Z => n39774);
   U26858 : BUF_X1 port map( A => n33442, Z => n39744);
   U26859 : BUF_X1 port map( A => n34710, Z => n39522);
   U26860 : BUF_X1 port map( A => n34716, Z => n39492);
   U26861 : BUF_X1 port map( A => n33436, Z => n39773);
   U26862 : BUF_X1 port map( A => n33442, Z => n39743);
   U26863 : BUF_X1 port map( A => n34710, Z => n39521);
   U26864 : BUF_X1 port map( A => n34716, Z => n39491);
   U26865 : BUF_X1 port map( A => n33436, Z => n39772);
   U26866 : BUF_X1 port map( A => n33442, Z => n39742);
   U26867 : BUF_X1 port map( A => n34710, Z => n39520);
   U26868 : BUF_X1 port map( A => n34716, Z => n39490);
   U26869 : BUF_X1 port map( A => n35991, Z => n39271);
   U26870 : BUF_X1 port map( A => n35997, Z => n39241);
   U26871 : BUF_X1 port map( A => n35991, Z => n39272);
   U26872 : BUF_X1 port map( A => n35997, Z => n39242);
   U26873 : BUF_X1 port map( A => n35991, Z => n39273);
   U26874 : BUF_X1 port map( A => n35997, Z => n39243);
   U26875 : BUF_X1 port map( A => n35991, Z => n39270);
   U26876 : BUF_X1 port map( A => n35997, Z => n39240);
   U26877 : BUF_X1 port map( A => n35991, Z => n39274);
   U26878 : BUF_X1 port map( A => n35997, Z => n39244);
   U26879 : BUF_X1 port map( A => n33482, Z => n39566);
   U26880 : BUF_X1 port map( A => n34756, Z => n39314);
   U26881 : BUF_X1 port map( A => n33482, Z => n39565);
   U26882 : BUF_X1 port map( A => n34756, Z => n39313);
   U26883 : BUF_X1 port map( A => n33482, Z => n39564);
   U26884 : BUF_X1 port map( A => n34756, Z => n39312);
   U26885 : BUF_X1 port map( A => n33482, Z => n39563);
   U26886 : BUF_X1 port map( A => n34756, Z => n39311);
   U26887 : BUF_X1 port map( A => n33482, Z => n39562);
   U26888 : BUF_X1 port map( A => n34756, Z => n39310);
   U26889 : BUF_X1 port map( A => n36037, Z => n39061);
   U26890 : BUF_X1 port map( A => n36019, Z => n39151);
   U26891 : BUF_X1 port map( A => n36009, Z => n39181);
   U26892 : BUF_X1 port map( A => n36037, Z => n39062);
   U26893 : BUF_X1 port map( A => n36019, Z => n39152);
   U26894 : BUF_X1 port map( A => n36009, Z => n39182);
   U26895 : BUF_X1 port map( A => n36037, Z => n39063);
   U26896 : BUF_X1 port map( A => n36019, Z => n39153);
   U26897 : BUF_X1 port map( A => n36009, Z => n39183);
   U26898 : BUF_X1 port map( A => n36037, Z => n39060);
   U26899 : BUF_X1 port map( A => n36019, Z => n39150);
   U26900 : BUF_X1 port map( A => n36009, Z => n39180);
   U26901 : BUF_X1 port map( A => n36037, Z => n39064);
   U26902 : BUF_X1 port map( A => n36019, Z => n39154);
   U26903 : BUF_X1 port map( A => n36009, Z => n39184);
   U26904 : BUF_X1 port map( A => n36003, Z => n39211);
   U26905 : BUF_X1 port map( A => n36003, Z => n39212);
   U26906 : BUF_X1 port map( A => n36003, Z => n39213);
   U26907 : BUF_X1 port map( A => n36003, Z => n39210);
   U26908 : BUF_X1 port map( A => n36003, Z => n39214);
   U26909 : BUF_X1 port map( A => n33470, Z => n39626);
   U26910 : BUF_X1 port map( A => n33454, Z => n39686);
   U26911 : BUF_X1 port map( A => n34744, Z => n39374);
   U26912 : BUF_X1 port map( A => n34728, Z => n39434);
   U26913 : BUF_X1 port map( A => n33470, Z => n39625);
   U26914 : BUF_X1 port map( A => n33454, Z => n39685);
   U26915 : BUF_X1 port map( A => n34744, Z => n39373);
   U26916 : BUF_X1 port map( A => n34728, Z => n39433);
   U26917 : BUF_X1 port map( A => n33470, Z => n39624);
   U26918 : BUF_X1 port map( A => n33454, Z => n39684);
   U26919 : BUF_X1 port map( A => n34744, Z => n39372);
   U26920 : BUF_X1 port map( A => n34728, Z => n39432);
   U26921 : BUF_X1 port map( A => n33470, Z => n39623);
   U26922 : BUF_X1 port map( A => n33454, Z => n39683);
   U26923 : BUF_X1 port map( A => n34744, Z => n39371);
   U26924 : BUF_X1 port map( A => n34728, Z => n39431);
   U26925 : BUF_X1 port map( A => n33470, Z => n39622);
   U26926 : BUF_X1 port map( A => n33454, Z => n39682);
   U26927 : BUF_X1 port map( A => n34744, Z => n39370);
   U26928 : BUF_X1 port map( A => n34728, Z => n39430);
   U26929 : BUF_X1 port map( A => n36031, Z => n39091);
   U26930 : BUF_X1 port map( A => n36031, Z => n39092);
   U26931 : BUF_X1 port map( A => n36031, Z => n39093);
   U26932 : BUF_X1 port map( A => n36031, Z => n39090);
   U26933 : BUF_X1 port map( A => n36031, Z => n39094);
   U26934 : BUF_X1 port map( A => n33476, Z => n39596);
   U26935 : BUF_X1 port map( A => n33448, Z => n39716);
   U26936 : BUF_X1 port map( A => n34750, Z => n39344);
   U26937 : BUF_X1 port map( A => n34722, Z => n39464);
   U26938 : BUF_X1 port map( A => n33476, Z => n39595);
   U26939 : BUF_X1 port map( A => n33448, Z => n39715);
   U26940 : BUF_X1 port map( A => n34750, Z => n39343);
   U26941 : BUF_X1 port map( A => n34722, Z => n39463);
   U26942 : BUF_X1 port map( A => n33476, Z => n39594);
   U26943 : BUF_X1 port map( A => n33448, Z => n39714);
   U26944 : BUF_X1 port map( A => n34750, Z => n39342);
   U26945 : BUF_X1 port map( A => n34722, Z => n39462);
   U26946 : BUF_X1 port map( A => n33476, Z => n39593);
   U26947 : BUF_X1 port map( A => n33448, Z => n39713);
   U26948 : BUF_X1 port map( A => n34750, Z => n39341);
   U26949 : BUF_X1 port map( A => n34722, Z => n39461);
   U26950 : BUF_X1 port map( A => n33476, Z => n39592);
   U26951 : BUF_X1 port map( A => n33448, Z => n39712);
   U26952 : BUF_X1 port map( A => n34750, Z => n39340);
   U26953 : BUF_X1 port map( A => n34722, Z => n39460);
   U26954 : BUF_X1 port map( A => n33437, Z => n39770);
   U26955 : BUF_X1 port map( A => n33443, Z => n39740);
   U26956 : BUF_X1 port map( A => n34711, Z => n39518);
   U26957 : BUF_X1 port map( A => n34717, Z => n39488);
   U26958 : BUF_X1 port map( A => n33437, Z => n39769);
   U26959 : BUF_X1 port map( A => n33443, Z => n39739);
   U26960 : BUF_X1 port map( A => n34711, Z => n39517);
   U26961 : BUF_X1 port map( A => n34717, Z => n39487);
   U26962 : BUF_X1 port map( A => n33437, Z => n39768);
   U26963 : BUF_X1 port map( A => n33443, Z => n39738);
   U26964 : BUF_X1 port map( A => n34711, Z => n39516);
   U26965 : BUF_X1 port map( A => n34717, Z => n39486);
   U26966 : BUF_X1 port map( A => n33437, Z => n39767);
   U26967 : BUF_X1 port map( A => n33443, Z => n39737);
   U26968 : BUF_X1 port map( A => n34711, Z => n39515);
   U26969 : BUF_X1 port map( A => n34717, Z => n39485);
   U26970 : BUF_X1 port map( A => n33437, Z => n39766);
   U26971 : BUF_X1 port map( A => n33443, Z => n39736);
   U26972 : BUF_X1 port map( A => n34711, Z => n39514);
   U26973 : BUF_X1 port map( A => n34717, Z => n39484);
   U26974 : BUF_X1 port map( A => n36025, Z => n39121);
   U26975 : BUF_X1 port map( A => n36025, Z => n39122);
   U26976 : BUF_X1 port map( A => n36025, Z => n39123);
   U26977 : BUF_X1 port map( A => n36025, Z => n39120);
   U26978 : BUF_X1 port map( A => n36025, Z => n39124);
   U26979 : BUF_X1 port map( A => n33464, Z => n39656);
   U26980 : BUF_X1 port map( A => n34738, Z => n39404);
   U26981 : BUF_X1 port map( A => n33464, Z => n39655);
   U26982 : BUF_X1 port map( A => n34738, Z => n39403);
   U26983 : BUF_X1 port map( A => n33464, Z => n39654);
   U26984 : BUF_X1 port map( A => n34738, Z => n39402);
   U26985 : BUF_X1 port map( A => n33464, Z => n39653);
   U26986 : BUF_X1 port map( A => n34738, Z => n39401);
   U26987 : BUF_X1 port map( A => n33464, Z => n39652);
   U26988 : BUF_X1 port map( A => n34738, Z => n39400);
   U26989 : BUF_X1 port map( A => n33477, Z => n39590);
   U26990 : BUF_X1 port map( A => n34751, Z => n39338);
   U26991 : BUF_X1 port map( A => n33477, Z => n39589);
   U26992 : BUF_X1 port map( A => n34751, Z => n39337);
   U26993 : BUF_X1 port map( A => n33477, Z => n39588);
   U26994 : BUF_X1 port map( A => n34751, Z => n39336);
   U26995 : BUF_X1 port map( A => n33477, Z => n39587);
   U26996 : BUF_X1 port map( A => n34751, Z => n39335);
   U26997 : BUF_X1 port map( A => n33477, Z => n39586);
   U26998 : BUF_X1 port map( A => n34751, Z => n39334);
   U26999 : BUF_X1 port map( A => n35992, Z => n39265);
   U27000 : BUF_X1 port map( A => n35998, Z => n39235);
   U27001 : BUF_X1 port map( A => n35992, Z => n39266);
   U27002 : BUF_X1 port map( A => n35998, Z => n39236);
   U27003 : BUF_X1 port map( A => n35992, Z => n39267);
   U27004 : BUF_X1 port map( A => n35998, Z => n39237);
   U27005 : BUF_X1 port map( A => n35992, Z => n39264);
   U27006 : BUF_X1 port map( A => n35998, Z => n39234);
   U27007 : BUF_X1 port map( A => n35992, Z => n39268);
   U27008 : BUF_X1 port map( A => n35998, Z => n39238);
   U27009 : BUF_X1 port map( A => n33465, Z => n39650);
   U27010 : BUF_X1 port map( A => n33449, Z => n39710);
   U27011 : BUF_X1 port map( A => n34739, Z => n39398);
   U27012 : BUF_X1 port map( A => n34723, Z => n39458);
   U27013 : BUF_X1 port map( A => n33465, Z => n39649);
   U27014 : BUF_X1 port map( A => n33449, Z => n39709);
   U27015 : BUF_X1 port map( A => n34739, Z => n39397);
   U27016 : BUF_X1 port map( A => n34723, Z => n39457);
   U27017 : BUF_X1 port map( A => n33465, Z => n39648);
   U27018 : BUF_X1 port map( A => n33449, Z => n39708);
   U27019 : BUF_X1 port map( A => n34739, Z => n39396);
   U27020 : BUF_X1 port map( A => n34723, Z => n39456);
   U27021 : BUF_X1 port map( A => n33465, Z => n39647);
   U27022 : BUF_X1 port map( A => n33449, Z => n39707);
   U27023 : BUF_X1 port map( A => n34739, Z => n39395);
   U27024 : BUF_X1 port map( A => n34723, Z => n39455);
   U27025 : BUF_X1 port map( A => n33465, Z => n39646);
   U27026 : BUF_X1 port map( A => n33449, Z => n39706);
   U27027 : BUF_X1 port map( A => n34739, Z => n39394);
   U27028 : BUF_X1 port map( A => n34723, Z => n39454);
   U27029 : BUF_X1 port map( A => n33483, Z => n39560);
   U27030 : BUF_X1 port map( A => n34757, Z => n39308);
   U27031 : BUF_X1 port map( A => n33483, Z => n39559);
   U27032 : BUF_X1 port map( A => n34757, Z => n39307);
   U27033 : BUF_X1 port map( A => n33483, Z => n39558);
   U27034 : BUF_X1 port map( A => n34757, Z => n39306);
   U27035 : BUF_X1 port map( A => n33483, Z => n39557);
   U27036 : BUF_X1 port map( A => n34757, Z => n39305);
   U27037 : BUF_X1 port map( A => n33483, Z => n39556);
   U27038 : BUF_X1 port map( A => n34757, Z => n39304);
   U27039 : BUF_X1 port map( A => n36038, Z => n39055);
   U27040 : BUF_X1 port map( A => n36010, Z => n39175);
   U27041 : BUF_X1 port map( A => n36038, Z => n39056);
   U27042 : BUF_X1 port map( A => n36010, Z => n39176);
   U27043 : BUF_X1 port map( A => n36038, Z => n39057);
   U27044 : BUF_X1 port map( A => n36010, Z => n39177);
   U27045 : BUF_X1 port map( A => n36038, Z => n39054);
   U27046 : BUF_X1 port map( A => n36010, Z => n39174);
   U27047 : BUF_X1 port map( A => n36038, Z => n39058);
   U27048 : BUF_X1 port map( A => n36010, Z => n39178);
   U27049 : BUF_X1 port map( A => n36020, Z => n39145);
   U27050 : BUF_X1 port map( A => n36020, Z => n39146);
   U27051 : BUF_X1 port map( A => n36020, Z => n39147);
   U27052 : BUF_X1 port map( A => n36020, Z => n39144);
   U27053 : BUF_X1 port map( A => n36020, Z => n39148);
   U27054 : BUF_X1 port map( A => n36004, Z => n39205);
   U27055 : BUF_X1 port map( A => n36004, Z => n39206);
   U27056 : BUF_X1 port map( A => n36004, Z => n39207);
   U27057 : BUF_X1 port map( A => n36004, Z => n39204);
   U27058 : BUF_X1 port map( A => n36004, Z => n39208);
   U27059 : BUF_X1 port map( A => n36032, Z => n39085);
   U27060 : BUF_X1 port map( A => n36026, Z => n39115);
   U27061 : BUF_X1 port map( A => n36032, Z => n39086);
   U27062 : BUF_X1 port map( A => n36026, Z => n39116);
   U27063 : BUF_X1 port map( A => n36032, Z => n39087);
   U27064 : BUF_X1 port map( A => n36026, Z => n39117);
   U27065 : BUF_X1 port map( A => n36032, Z => n39084);
   U27066 : BUF_X1 port map( A => n36026, Z => n39114);
   U27067 : BUF_X1 port map( A => n36032, Z => n39088);
   U27068 : BUF_X1 port map( A => n36026, Z => n39118);
   U27069 : BUF_X1 port map( A => n33471, Z => n39620);
   U27070 : BUF_X1 port map( A => n33455, Z => n39680);
   U27071 : BUF_X1 port map( A => n34745, Z => n39368);
   U27072 : BUF_X1 port map( A => n34729, Z => n39428);
   U27073 : BUF_X1 port map( A => n33471, Z => n39619);
   U27074 : BUF_X1 port map( A => n33455, Z => n39679);
   U27075 : BUF_X1 port map( A => n34745, Z => n39367);
   U27076 : BUF_X1 port map( A => n34729, Z => n39427);
   U27077 : BUF_X1 port map( A => n33471, Z => n39618);
   U27078 : BUF_X1 port map( A => n33455, Z => n39678);
   U27079 : BUF_X1 port map( A => n34745, Z => n39366);
   U27080 : BUF_X1 port map( A => n34729, Z => n39426);
   U27081 : BUF_X1 port map( A => n33471, Z => n39617);
   U27082 : BUF_X1 port map( A => n33455, Z => n39677);
   U27083 : BUF_X1 port map( A => n34745, Z => n39365);
   U27084 : BUF_X1 port map( A => n34729, Z => n39425);
   U27085 : BUF_X1 port map( A => n33471, Z => n39616);
   U27086 : BUF_X1 port map( A => n33455, Z => n39676);
   U27087 : BUF_X1 port map( A => n34745, Z => n39364);
   U27088 : BUF_X1 port map( A => n34729, Z => n39424);
   U27089 : BUF_X1 port map( A => n33405, Z => n39901);
   U27090 : BUF_X1 port map( A => n33401, Z => n39920);
   U27091 : BUF_X1 port map( A => n33384, Z => n39999);
   U27092 : BUF_X1 port map( A => n33381, Z => n40018);
   U27093 : BUF_X1 port map( A => n33365, Z => n40097);
   U27094 : BUF_X1 port map( A => n33420, Z => n39802);
   U27095 : BUF_X1 port map( A => n33405, Z => n39904);
   U27096 : BUF_X1 port map( A => n33405, Z => n39903);
   U27097 : BUF_X1 port map( A => n33405, Z => n39902);
   U27098 : BUF_X1 port map( A => n33401, Z => n39923);
   U27099 : BUF_X1 port map( A => n33401, Z => n39922);
   U27100 : BUF_X1 port map( A => n33401, Z => n39921);
   U27101 : BUF_X1 port map( A => n33384, Z => n40002);
   U27102 : BUF_X1 port map( A => n33384, Z => n40001);
   U27103 : BUF_X1 port map( A => n33384, Z => n40000);
   U27104 : BUF_X1 port map( A => n33381, Z => n40021);
   U27105 : BUF_X1 port map( A => n33381, Z => n40020);
   U27106 : BUF_X1 port map( A => n33381, Z => n40019);
   U27107 : BUF_X1 port map( A => n33405, Z => n39905);
   U27108 : BUF_X1 port map( A => n33401, Z => n39924);
   U27109 : BUF_X1 port map( A => n33384, Z => n40003);
   U27110 : BUF_X1 port map( A => n33381, Z => n40022);
   U27111 : BUF_X1 port map( A => n33361, Z => n40117);
   U27112 : BUF_X1 port map( A => n33361, Z => n40118);
   U27113 : BUF_X1 port map( A => n33361, Z => n40119);
   U27114 : BUF_X1 port map( A => n33361, Z => n40120);
   U27115 : BUF_X1 port map( A => n33365, Z => n40101);
   U27116 : BUF_X1 port map( A => n33365, Z => n40100);
   U27117 : BUF_X1 port map( A => n33365, Z => n40099);
   U27118 : BUF_X1 port map( A => n33365, Z => n40098);
   U27119 : BUF_X1 port map( A => n33420, Z => n39804);
   U27120 : BUF_X1 port map( A => n33420, Z => n39803);
   U27121 : BUF_X1 port map( A => n33420, Z => n39806);
   U27122 : BUF_X1 port map( A => n33420, Z => n39805);
   U27123 : BUF_X1 port map( A => n33311, Z => n40397);
   U27124 : BUF_X1 port map( A => n33311, Z => n40398);
   U27125 : BUF_X1 port map( A => n33311, Z => n40399);
   U27126 : BUF_X1 port map( A => n33311, Z => n40400);
   U27127 : BUF_X1 port map( A => n33349, Z => n40197);
   U27128 : BUF_X1 port map( A => n33349, Z => n40198);
   U27129 : BUF_X1 port map( A => n33349, Z => n40199);
   U27130 : BUF_X1 port map( A => n33349, Z => n40200);
   U27131 : BUF_X1 port map( A => n33311, Z => n40396);
   U27132 : BUF_X1 port map( A => n33349, Z => n40196);
   U27133 : BUF_X1 port map( A => n33317, Z => n40356);
   U27134 : BUF_X1 port map( A => n33317, Z => n40357);
   U27135 : BUF_X1 port map( A => n33317, Z => n40358);
   U27136 : BUF_X1 port map( A => n33317, Z => n40359);
   U27137 : BUF_X1 port map( A => n33317, Z => n40360);
   U27138 : BUF_X1 port map( A => n33343, Z => n40236);
   U27139 : BUF_X1 port map( A => n33343, Z => n40237);
   U27140 : BUF_X1 port map( A => n33343, Z => n40238);
   U27141 : BUF_X1 port map( A => n33343, Z => n40239);
   U27142 : BUF_X1 port map( A => n33343, Z => n40240);
   U27143 : BUF_X1 port map( A => n33372, Z => n40077);
   U27144 : BUF_X1 port map( A => n33372, Z => n40078);
   U27145 : BUF_X1 port map( A => n33372, Z => n40079);
   U27146 : BUF_X1 port map( A => n33372, Z => n40080);
   U27147 : BUF_X1 port map( A => n33372, Z => n40081);
   U27148 : BUF_X1 port map( A => n33378, Z => n40037);
   U27149 : BUF_X1 port map( A => n33378, Z => n40038);
   U27150 : BUF_X1 port map( A => n33378, Z => n40039);
   U27151 : BUF_X1 port map( A => n33378, Z => n40040);
   U27152 : BUF_X1 port map( A => n33378, Z => n40041);
   U27153 : BUF_X1 port map( A => n33346, Z => n40217);
   U27154 : BUF_X1 port map( A => n33346, Z => n40218);
   U27155 : BUF_X1 port map( A => n33346, Z => n40219);
   U27156 : BUF_X1 port map( A => n33346, Z => n40220);
   U27157 : BUF_X1 port map( A => n33346, Z => n40216);
   U27158 : BUF_X1 port map( A => n33314, Z => n40376);
   U27159 : BUF_X1 port map( A => n33314, Z => n40377);
   U27160 : BUF_X1 port map( A => n33314, Z => n40378);
   U27161 : BUF_X1 port map( A => n33314, Z => n40379);
   U27162 : BUF_X1 port map( A => n33314, Z => n40380);
   U27163 : BUF_X1 port map( A => n33375, Z => n40057);
   U27164 : BUF_X1 port map( A => n33375, Z => n40058);
   U27165 : BUF_X1 port map( A => n33375, Z => n40059);
   U27166 : BUF_X1 port map( A => n33375, Z => n40060);
   U27167 : BUF_X1 port map( A => n33375, Z => n40061);
   U27168 : BUF_X1 port map( A => n33304, Z => n40417);
   U27169 : BUF_X1 port map( A => n33304, Z => n40418);
   U27170 : BUF_X1 port map( A => n33304, Z => n40419);
   U27171 : BUF_X1 port map( A => n33304, Z => n40420);
   U27172 : BUF_X1 port map( A => n33326, Z => n40297);
   U27173 : BUF_X1 port map( A => n33326, Z => n40298);
   U27174 : BUF_X1 port map( A => n33326, Z => n40299);
   U27175 : BUF_X1 port map( A => n33326, Z => n40300);
   U27176 : BUF_X1 port map( A => n33323, Z => n40317);
   U27177 : BUF_X1 port map( A => n33323, Z => n40318);
   U27178 : BUF_X1 port map( A => n33323, Z => n40319);
   U27179 : BUF_X1 port map( A => n33323, Z => n40320);
   U27180 : BUF_X1 port map( A => n33417, Z => n39822);
   U27181 : BUF_X1 port map( A => n33417, Z => n39823);
   U27182 : BUF_X1 port map( A => n33417, Z => n39824);
   U27183 : BUF_X1 port map( A => n33417, Z => n39825);
   U27184 : BUF_X1 port map( A => n33304, Z => n40416);
   U27185 : BUF_X1 port map( A => n33326, Z => n40296);
   U27186 : BUF_X1 port map( A => n33323, Z => n40316);
   U27187 : BUF_X1 port map( A => n33417, Z => n39821);
   U27188 : BUF_X1 port map( A => n33320, Z => n40336);
   U27189 : BUF_X1 port map( A => n33320, Z => n40337);
   U27190 : BUF_X1 port map( A => n33320, Z => n40338);
   U27191 : BUF_X1 port map( A => n33320, Z => n40339);
   U27192 : BUF_X1 port map( A => n33320, Z => n40340);
   U27193 : BUF_X1 port map( A => n33329, Z => n40276);
   U27194 : BUF_X1 port map( A => n33329, Z => n40277);
   U27195 : BUF_X1 port map( A => n33329, Z => n40278);
   U27196 : BUF_X1 port map( A => n33329, Z => n40279);
   U27197 : BUF_X1 port map( A => n33329, Z => n40280);
   U27198 : BUF_X1 port map( A => n33336, Z => n40256);
   U27199 : BUF_X1 port map( A => n33336, Z => n40257);
   U27200 : BUF_X1 port map( A => n33336, Z => n40258);
   U27201 : BUF_X1 port map( A => n33336, Z => n40259);
   U27202 : BUF_X1 port map( A => n33336, Z => n40260);
   U27203 : BUF_X1 port map( A => n33352, Z => n40176);
   U27204 : BUF_X1 port map( A => n33352, Z => n40177);
   U27205 : BUF_X1 port map( A => n33352, Z => n40178);
   U27206 : BUF_X1 port map( A => n33352, Z => n40179);
   U27207 : BUF_X1 port map( A => n33352, Z => n40180);
   U27208 : BUF_X1 port map( A => n33355, Z => n40156);
   U27209 : BUF_X1 port map( A => n33355, Z => n40157);
   U27210 : BUF_X1 port map( A => n33355, Z => n40158);
   U27211 : BUF_X1 port map( A => n33355, Z => n40159);
   U27212 : BUF_X1 port map( A => n33355, Z => n40160);
   U27213 : BUF_X1 port map( A => n33358, Z => n40136);
   U27214 : BUF_X1 port map( A => n33358, Z => n40137);
   U27215 : BUF_X1 port map( A => n33358, Z => n40138);
   U27216 : BUF_X1 port map( A => n33358, Z => n40139);
   U27217 : BUF_X1 port map( A => n33358, Z => n40140);
   U27218 : BUF_X1 port map( A => n33387, Z => n39979);
   U27219 : BUF_X1 port map( A => n33387, Z => n39980);
   U27220 : BUF_X1 port map( A => n33387, Z => n39981);
   U27221 : BUF_X1 port map( A => n33387, Z => n39982);
   U27222 : BUF_X1 port map( A => n33387, Z => n39983);
   U27223 : BUF_X1 port map( A => n33390, Z => n39959);
   U27224 : BUF_X1 port map( A => n33390, Z => n39960);
   U27225 : BUF_X1 port map( A => n33390, Z => n39961);
   U27226 : BUF_X1 port map( A => n33390, Z => n39962);
   U27227 : BUF_X1 port map( A => n33390, Z => n39963);
   U27228 : BUF_X1 port map( A => n33393, Z => n39939);
   U27229 : BUF_X1 port map( A => n33393, Z => n39940);
   U27230 : BUF_X1 port map( A => n33393, Z => n39941);
   U27231 : BUF_X1 port map( A => n33393, Z => n39942);
   U27232 : BUF_X1 port map( A => n33393, Z => n39943);
   U27233 : BUF_X1 port map( A => n33408, Z => n39881);
   U27234 : BUF_X1 port map( A => n33408, Z => n39882);
   U27235 : BUF_X1 port map( A => n33408, Z => n39883);
   U27236 : BUF_X1 port map( A => n33408, Z => n39884);
   U27237 : BUF_X1 port map( A => n33408, Z => n39885);
   U27238 : BUF_X1 port map( A => n33411, Z => n39861);
   U27239 : BUF_X1 port map( A => n33411, Z => n39862);
   U27240 : BUF_X1 port map( A => n33411, Z => n39863);
   U27241 : BUF_X1 port map( A => n33411, Z => n39864);
   U27242 : BUF_X1 port map( A => n33411, Z => n39865);
   U27243 : BUF_X1 port map( A => n33414, Z => n39841);
   U27244 : BUF_X1 port map( A => n33414, Z => n39842);
   U27245 : BUF_X1 port map( A => n33414, Z => n39843);
   U27246 : BUF_X1 port map( A => n33414, Z => n39844);
   U27247 : BUF_X1 port map( A => n33414, Z => n39845);
   U27248 : BUF_X1 port map( A => n33361, Z => n40116);
   U27249 : BUF_X1 port map( A => n40589, Z => n40592);
   U27250 : BUF_X1 port map( A => n40589, Z => n40591);
   U27251 : BUF_X1 port map( A => n40589, Z => n40594);
   U27252 : BUF_X1 port map( A => n40589, Z => n40593);
   U27253 : BUF_X1 port map( A => n40589, Z => n40590);
   U27254 : BUF_X1 port map( A => n40429, Z => n40430);
   U27255 : BUF_X1 port map( A => n40429, Z => n40434);
   U27256 : BUF_X1 port map( A => n40429, Z => n40433);
   U27257 : BUF_X1 port map( A => n40429, Z => n40432);
   U27258 : BUF_X1 port map( A => n40429, Z => n40431);
   U27259 : BUF_X1 port map( A => n40409, Z => n40410);
   U27260 : BUF_X1 port map( A => n40209, Z => n40210);
   U27261 : BUF_X1 port map( A => n40229, Z => n40230);
   U27262 : BUF_X1 port map( A => n40409, Z => n40414);
   U27263 : BUF_X1 port map( A => n40409, Z => n40413);
   U27264 : BUF_X1 port map( A => n40409, Z => n40412);
   U27265 : BUF_X1 port map( A => n40409, Z => n40411);
   U27266 : BUF_X1 port map( A => n40209, Z => n40214);
   U27267 : BUF_X1 port map( A => n40209, Z => n40213);
   U27268 : BUF_X1 port map( A => n40209, Z => n40212);
   U27269 : BUF_X1 port map( A => n40209, Z => n40211);
   U27270 : BUF_X1 port map( A => n40229, Z => n40234);
   U27271 : BUF_X1 port map( A => n40229, Z => n40233);
   U27272 : BUF_X1 port map( A => n40229, Z => n40232);
   U27273 : BUF_X1 port map( A => n40229, Z => n40231);
   U27274 : BUF_X1 port map( A => n40011, Z => n40012);
   U27275 : BUF_X1 port map( A => n40030, Z => n40031);
   U27276 : BUF_X1 port map( A => n40011, Z => n40016);
   U27277 : BUF_X1 port map( A => n40011, Z => n40015);
   U27278 : BUF_X1 port map( A => n40011, Z => n40014);
   U27279 : BUF_X1 port map( A => n40011, Z => n40013);
   U27280 : BUF_X1 port map( A => n40030, Z => n40035);
   U27281 : BUF_X1 port map( A => n40030, Z => n40034);
   U27282 : BUF_X1 port map( A => n40030, Z => n40033);
   U27283 : BUF_X1 port map( A => n40030, Z => n40032);
   U27284 : BUF_X1 port map( A => n40309, Z => n40310);
   U27285 : BUF_X1 port map( A => n40329, Z => n40330);
   U27286 : BUF_X1 port map( A => n39834, Z => n39835);
   U27287 : BUF_X1 port map( A => n40309, Z => n40314);
   U27288 : BUF_X1 port map( A => n40309, Z => n40313);
   U27289 : BUF_X1 port map( A => n40309, Z => n40312);
   U27290 : BUF_X1 port map( A => n40309, Z => n40311);
   U27291 : BUF_X1 port map( A => n40329, Z => n40334);
   U27292 : BUF_X1 port map( A => n40329, Z => n40333);
   U27293 : BUF_X1 port map( A => n40329, Z => n40332);
   U27294 : BUF_X1 port map( A => n40329, Z => n40331);
   U27295 : BUF_X1 port map( A => n39834, Z => n39839);
   U27296 : BUF_X1 port map( A => n39834, Z => n39838);
   U27297 : BUF_X1 port map( A => n39834, Z => n39837);
   U27298 : BUF_X1 port map( A => n39834, Z => n39836);
   U27299 : BUF_X1 port map( A => n39814, Z => n39817);
   U27300 : BUF_X1 port map( A => n39814, Z => n39816);
   U27301 : BUF_X1 port map( A => n39814, Z => n39815);
   U27302 : BUF_X1 port map( A => n40529, Z => n40530);
   U27303 : BUF_X1 port map( A => n40529, Z => n40534);
   U27304 : BUF_X1 port map( A => n40529, Z => n40533);
   U27305 : BUF_X1 port map( A => n40529, Z => n40532);
   U27306 : BUF_X1 port map( A => n40529, Z => n40531);
   U27307 : BUF_X1 port map( A => n40509, Z => n40510);
   U27308 : BUF_X1 port map( A => n40509, Z => n40514);
   U27309 : BUF_X1 port map( A => n40509, Z => n40513);
   U27310 : BUF_X1 port map( A => n40509, Z => n40512);
   U27311 : BUF_X1 port map( A => n40509, Z => n40511);
   U27312 : BUF_X1 port map( A => n40569, Z => n40574);
   U27313 : BUF_X1 port map( A => n40569, Z => n40573);
   U27314 : BUF_X1 port map( A => n40569, Z => n40572);
   U27315 : BUF_X1 port map( A => n40569, Z => n40571);
   U27316 : BUF_X1 port map( A => n40569, Z => n40570);
   U27317 : BUF_X1 port map( A => n40549, Z => n40554);
   U27318 : BUF_X1 port map( A => n40549, Z => n40553);
   U27319 : BUF_X1 port map( A => n40549, Z => n40552);
   U27320 : BUF_X1 port map( A => n40549, Z => n40551);
   U27321 : BUF_X1 port map( A => n40549, Z => n40550);
   U27322 : BUF_X1 port map( A => n40489, Z => n40494);
   U27323 : BUF_X1 port map( A => n40489, Z => n40493);
   U27324 : BUF_X1 port map( A => n40489, Z => n40492);
   U27325 : BUF_X1 port map( A => n40489, Z => n40491);
   U27326 : BUF_X1 port map( A => n40489, Z => n40490);
   U27327 : BUF_X1 port map( A => n40469, Z => n40474);
   U27328 : BUF_X1 port map( A => n40469, Z => n40473);
   U27329 : BUF_X1 port map( A => n40469, Z => n40472);
   U27330 : BUF_X1 port map( A => n40469, Z => n40471);
   U27331 : BUF_X1 port map( A => n40469, Z => n40470);
   U27332 : BUF_X1 port map( A => n40449, Z => n40454);
   U27333 : BUF_X1 port map( A => n40449, Z => n40453);
   U27334 : BUF_X1 port map( A => n40449, Z => n40452);
   U27335 : BUF_X1 port map( A => n40449, Z => n40451);
   U27336 : BUF_X1 port map( A => n40449, Z => n40450);
   U27337 : BUF_X1 port map( A => n40389, Z => n40394);
   U27338 : BUF_X1 port map( A => n40389, Z => n40393);
   U27339 : BUF_X1 port map( A => n40389, Z => n40392);
   U27340 : BUF_X1 port map( A => n40389, Z => n40391);
   U27341 : BUF_X1 port map( A => n40389, Z => n40390);
   U27342 : BUF_X1 port map( A => n40369, Z => n40374);
   U27343 : BUF_X1 port map( A => n40369, Z => n40373);
   U27344 : BUF_X1 port map( A => n40369, Z => n40372);
   U27345 : BUF_X1 port map( A => n40369, Z => n40371);
   U27346 : BUF_X1 port map( A => n40369, Z => n40370);
   U27347 : BUF_X1 port map( A => n40349, Z => n40354);
   U27348 : BUF_X1 port map( A => n40349, Z => n40353);
   U27349 : BUF_X1 port map( A => n40349, Z => n40352);
   U27350 : BUF_X1 port map( A => n40349, Z => n40351);
   U27351 : BUF_X1 port map( A => n40349, Z => n40350);
   U27352 : BUF_X1 port map( A => n40289, Z => n40294);
   U27353 : BUF_X1 port map( A => n40289, Z => n40293);
   U27354 : BUF_X1 port map( A => n40289, Z => n40292);
   U27355 : BUF_X1 port map( A => n40289, Z => n40291);
   U27356 : BUF_X1 port map( A => n40289, Z => n40290);
   U27357 : BUF_X1 port map( A => n40269, Z => n40274);
   U27358 : BUF_X1 port map( A => n40269, Z => n40273);
   U27359 : BUF_X1 port map( A => n40269, Z => n40272);
   U27360 : BUF_X1 port map( A => n40269, Z => n40271);
   U27361 : BUF_X1 port map( A => n40269, Z => n40270);
   U27362 : BUF_X1 port map( A => n40249, Z => n40254);
   U27363 : BUF_X1 port map( A => n40249, Z => n40253);
   U27364 : BUF_X1 port map( A => n40249, Z => n40252);
   U27365 : BUF_X1 port map( A => n40249, Z => n40251);
   U27366 : BUF_X1 port map( A => n40249, Z => n40250);
   U27367 : BUF_X1 port map( A => n40189, Z => n40194);
   U27368 : BUF_X1 port map( A => n40189, Z => n40193);
   U27369 : BUF_X1 port map( A => n40189, Z => n40192);
   U27370 : BUF_X1 port map( A => n40189, Z => n40191);
   U27371 : BUF_X1 port map( A => n40189, Z => n40190);
   U27372 : BUF_X1 port map( A => n40169, Z => n40174);
   U27373 : BUF_X1 port map( A => n40169, Z => n40173);
   U27374 : BUF_X1 port map( A => n40169, Z => n40172);
   U27375 : BUF_X1 port map( A => n40169, Z => n40171);
   U27376 : BUF_X1 port map( A => n40169, Z => n40170);
   U27377 : BUF_X1 port map( A => n40149, Z => n40154);
   U27378 : BUF_X1 port map( A => n40149, Z => n40153);
   U27379 : BUF_X1 port map( A => n40149, Z => n40152);
   U27380 : BUF_X1 port map( A => n40149, Z => n40151);
   U27381 : BUF_X1 port map( A => n40149, Z => n40150);
   U27382 : BUF_X1 port map( A => n40129, Z => n40134);
   U27383 : BUF_X1 port map( A => n40129, Z => n40133);
   U27384 : BUF_X1 port map( A => n40129, Z => n40132);
   U27385 : BUF_X1 port map( A => n40129, Z => n40131);
   U27386 : BUF_X1 port map( A => n40129, Z => n40130);
   U27387 : BUF_X1 port map( A => n40109, Z => n40114);
   U27388 : BUF_X1 port map( A => n40109, Z => n40113);
   U27389 : BUF_X1 port map( A => n40109, Z => n40112);
   U27390 : BUF_X1 port map( A => n40109, Z => n40111);
   U27391 : BUF_X1 port map( A => n40109, Z => n40110);
   U27392 : BUF_X1 port map( A => n40090, Z => n40095);
   U27393 : BUF_X1 port map( A => n40090, Z => n40094);
   U27394 : BUF_X1 port map( A => n40090, Z => n40093);
   U27395 : BUF_X1 port map( A => n40090, Z => n40092);
   U27396 : BUF_X1 port map( A => n40090, Z => n40091);
   U27397 : BUF_X1 port map( A => n40070, Z => n40075);
   U27398 : BUF_X1 port map( A => n40070, Z => n40074);
   U27399 : BUF_X1 port map( A => n40070, Z => n40073);
   U27400 : BUF_X1 port map( A => n40070, Z => n40072);
   U27401 : BUF_X1 port map( A => n40070, Z => n40071);
   U27402 : BUF_X1 port map( A => n40050, Z => n40055);
   U27403 : BUF_X1 port map( A => n40050, Z => n40054);
   U27404 : BUF_X1 port map( A => n40050, Z => n40053);
   U27405 : BUF_X1 port map( A => n40050, Z => n40052);
   U27406 : BUF_X1 port map( A => n40050, Z => n40051);
   U27407 : BUF_X1 port map( A => n39992, Z => n39997);
   U27408 : BUF_X1 port map( A => n39992, Z => n39996);
   U27409 : BUF_X1 port map( A => n39992, Z => n39995);
   U27410 : BUF_X1 port map( A => n39992, Z => n39994);
   U27411 : BUF_X1 port map( A => n39992, Z => n39993);
   U27412 : BUF_X1 port map( A => n39972, Z => n39977);
   U27413 : BUF_X1 port map( A => n39972, Z => n39976);
   U27414 : BUF_X1 port map( A => n39972, Z => n39975);
   U27415 : BUF_X1 port map( A => n39972, Z => n39974);
   U27416 : BUF_X1 port map( A => n39972, Z => n39973);
   U27417 : BUF_X1 port map( A => n39874, Z => n39879);
   U27418 : BUF_X1 port map( A => n39874, Z => n39878);
   U27419 : BUF_X1 port map( A => n39874, Z => n39877);
   U27420 : BUF_X1 port map( A => n39874, Z => n39876);
   U27421 : BUF_X1 port map( A => n39874, Z => n39875);
   U27422 : BUF_X1 port map( A => n39854, Z => n39859);
   U27423 : BUF_X1 port map( A => n39854, Z => n39858);
   U27424 : BUF_X1 port map( A => n39854, Z => n39857);
   U27425 : BUF_X1 port map( A => n39854, Z => n39856);
   U27426 : BUF_X1 port map( A => n39854, Z => n39855);
   U27427 : BUF_X1 port map( A => n39814, Z => n39819);
   U27428 : BUF_X1 port map( A => n39814, Z => n39818);
   U27429 : BUF_X1 port map( A => n40402, Z => n40403);
   U27430 : BUF_X1 port map( A => n39906, Z => n39907);
   U27431 : BUF_X1 port map( A => n39925, Z => n39926);
   U27432 : BUF_X1 port map( A => n40202, Z => n40203);
   U27433 : BUF_X1 port map( A => n40222, Z => n40223);
   U27434 : BUF_X1 port map( A => n40402, Z => n40407);
   U27435 : BUF_X1 port map( A => n40402, Z => n40406);
   U27436 : BUF_X1 port map( A => n40402, Z => n40405);
   U27437 : BUF_X1 port map( A => n40402, Z => n40404);
   U27438 : BUF_X1 port map( A => n39906, Z => n39911);
   U27439 : BUF_X1 port map( A => n39906, Z => n39910);
   U27440 : BUF_X1 port map( A => n39906, Z => n39909);
   U27441 : BUF_X1 port map( A => n39906, Z => n39908);
   U27442 : BUF_X1 port map( A => n39925, Z => n39930);
   U27443 : BUF_X1 port map( A => n39925, Z => n39929);
   U27444 : BUF_X1 port map( A => n39925, Z => n39928);
   U27445 : BUF_X1 port map( A => n39925, Z => n39927);
   U27446 : BUF_X1 port map( A => n40202, Z => n40207);
   U27447 : BUF_X1 port map( A => n40202, Z => n40206);
   U27448 : BUF_X1 port map( A => n40202, Z => n40205);
   U27449 : BUF_X1 port map( A => n40202, Z => n40204);
   U27450 : BUF_X1 port map( A => n40222, Z => n40227);
   U27451 : BUF_X1 port map( A => n40222, Z => n40226);
   U27452 : BUF_X1 port map( A => n40222, Z => n40225);
   U27453 : BUF_X1 port map( A => n40222, Z => n40224);
   U27454 : BUF_X1 port map( A => n40043, Z => n40046);
   U27455 : BUF_X1 port map( A => n40043, Z => n40045);
   U27456 : BUF_X1 port map( A => n40043, Z => n40044);
   U27457 : BUF_X1 port map( A => n39887, Z => n39892);
   U27458 : BUF_X1 port map( A => n39887, Z => n39891);
   U27459 : BUF_X1 port map( A => n39887, Z => n39890);
   U27460 : BUF_X1 port map( A => n39887, Z => n39889);
   U27461 : BUF_X1 port map( A => n39887, Z => n39888);
   U27462 : BUF_X1 port map( A => n40422, Z => n40423);
   U27463 : BUF_X1 port map( A => n40422, Z => n40427);
   U27464 : BUF_X1 port map( A => n40422, Z => n40426);
   U27465 : BUF_X1 port map( A => n40422, Z => n40425);
   U27466 : BUF_X1 port map( A => n40422, Z => n40424);
   U27467 : BUF_X1 port map( A => n40004, Z => n40005);
   U27468 : BUF_X1 port map( A => n40023, Z => n40024);
   U27469 : BUF_X1 port map( A => n40004, Z => n40009);
   U27470 : BUF_X1 port map( A => n40004, Z => n40008);
   U27471 : BUF_X1 port map( A => n40004, Z => n40007);
   U27472 : BUF_X1 port map( A => n40004, Z => n40006);
   U27473 : BUF_X1 port map( A => n40023, Z => n40028);
   U27474 : BUF_X1 port map( A => n40023, Z => n40027);
   U27475 : BUF_X1 port map( A => n40023, Z => n40026);
   U27476 : BUF_X1 port map( A => n40023, Z => n40025);
   U27477 : BUF_X1 port map( A => n40302, Z => n40303);
   U27478 : BUF_X1 port map( A => n40322, Z => n40323);
   U27479 : BUF_X1 port map( A => n40382, Z => n40387);
   U27480 : BUF_X1 port map( A => n40382, Z => n40386);
   U27481 : BUF_X1 port map( A => n40382, Z => n40385);
   U27482 : BUF_X1 port map( A => n40382, Z => n40384);
   U27483 : BUF_X1 port map( A => n40382, Z => n40383);
   U27484 : BUF_X1 port map( A => n40362, Z => n40367);
   U27485 : BUF_X1 port map( A => n40362, Z => n40366);
   U27486 : BUF_X1 port map( A => n40362, Z => n40365);
   U27487 : BUF_X1 port map( A => n40362, Z => n40364);
   U27488 : BUF_X1 port map( A => n40362, Z => n40363);
   U27489 : BUF_X1 port map( A => n40242, Z => n40247);
   U27490 : BUF_X1 port map( A => n40242, Z => n40246);
   U27491 : BUF_X1 port map( A => n40242, Z => n40245);
   U27492 : BUF_X1 port map( A => n40242, Z => n40244);
   U27493 : BUF_X1 port map( A => n40242, Z => n40243);
   U27494 : BUF_X1 port map( A => n40083, Z => n40088);
   U27495 : BUF_X1 port map( A => n40083, Z => n40087);
   U27496 : BUF_X1 port map( A => n40083, Z => n40086);
   U27497 : BUF_X1 port map( A => n40083, Z => n40085);
   U27498 : BUF_X1 port map( A => n40083, Z => n40084);
   U27499 : BUF_X1 port map( A => n40063, Z => n40068);
   U27500 : BUF_X1 port map( A => n40063, Z => n40067);
   U27501 : BUF_X1 port map( A => n40063, Z => n40066);
   U27502 : BUF_X1 port map( A => n40063, Z => n40065);
   U27503 : BUF_X1 port map( A => n40063, Z => n40064);
   U27504 : BUF_X1 port map( A => n40043, Z => n40048);
   U27505 : BUF_X1 port map( A => n40043, Z => n40047);
   U27506 : BUF_X1 port map( A => n39827, Z => n39828);
   U27507 : BUF_X1 port map( A => n40302, Z => n40307);
   U27508 : BUF_X1 port map( A => n40302, Z => n40306);
   U27509 : BUF_X1 port map( A => n40302, Z => n40305);
   U27510 : BUF_X1 port map( A => n40302, Z => n40304);
   U27511 : BUF_X1 port map( A => n40322, Z => n40327);
   U27512 : BUF_X1 port map( A => n40322, Z => n40326);
   U27513 : BUF_X1 port map( A => n40322, Z => n40325);
   U27514 : BUF_X1 port map( A => n40322, Z => n40324);
   U27515 : BUF_X1 port map( A => n39827, Z => n39832);
   U27516 : BUF_X1 port map( A => n39827, Z => n39831);
   U27517 : BUF_X1 port map( A => n39827, Z => n39830);
   U27518 : BUF_X1 port map( A => n39827, Z => n39829);
   U27519 : BUF_X1 port map( A => n39807, Z => n39810);
   U27520 : BUF_X1 port map( A => n39807, Z => n39809);
   U27521 : BUF_X1 port map( A => n39807, Z => n39808);
   U27522 : BUF_X1 port map( A => n40342, Z => n40347);
   U27523 : BUF_X1 port map( A => n40342, Z => n40346);
   U27524 : BUF_X1 port map( A => n40342, Z => n40345);
   U27525 : BUF_X1 port map( A => n40342, Z => n40344);
   U27526 : BUF_X1 port map( A => n40342, Z => n40343);
   U27527 : BUF_X1 port map( A => n40282, Z => n40287);
   U27528 : BUF_X1 port map( A => n40282, Z => n40286);
   U27529 : BUF_X1 port map( A => n40282, Z => n40285);
   U27530 : BUF_X1 port map( A => n40282, Z => n40284);
   U27531 : BUF_X1 port map( A => n40282, Z => n40283);
   U27532 : BUF_X1 port map( A => n40262, Z => n40267);
   U27533 : BUF_X1 port map( A => n40262, Z => n40266);
   U27534 : BUF_X1 port map( A => n40262, Z => n40265);
   U27535 : BUF_X1 port map( A => n40262, Z => n40264);
   U27536 : BUF_X1 port map( A => n40262, Z => n40263);
   U27537 : BUF_X1 port map( A => n40182, Z => n40187);
   U27538 : BUF_X1 port map( A => n40182, Z => n40186);
   U27539 : BUF_X1 port map( A => n40182, Z => n40185);
   U27540 : BUF_X1 port map( A => n40182, Z => n40184);
   U27541 : BUF_X1 port map( A => n40182, Z => n40183);
   U27542 : BUF_X1 port map( A => n40162, Z => n40167);
   U27543 : BUF_X1 port map( A => n40162, Z => n40166);
   U27544 : BUF_X1 port map( A => n40162, Z => n40165);
   U27545 : BUF_X1 port map( A => n40162, Z => n40164);
   U27546 : BUF_X1 port map( A => n40162, Z => n40163);
   U27547 : BUF_X1 port map( A => n40142, Z => n40147);
   U27548 : BUF_X1 port map( A => n40142, Z => n40146);
   U27549 : BUF_X1 port map( A => n40142, Z => n40145);
   U27550 : BUF_X1 port map( A => n40142, Z => n40144);
   U27551 : BUF_X1 port map( A => n40142, Z => n40143);
   U27552 : BUF_X1 port map( A => n40122, Z => n40127);
   U27553 : BUF_X1 port map( A => n40122, Z => n40126);
   U27554 : BUF_X1 port map( A => n40122, Z => n40125);
   U27555 : BUF_X1 port map( A => n40122, Z => n40124);
   U27556 : BUF_X1 port map( A => n40122, Z => n40123);
   U27557 : BUF_X1 port map( A => n40102, Z => n40107);
   U27558 : BUF_X1 port map( A => n40102, Z => n40106);
   U27559 : BUF_X1 port map( A => n40102, Z => n40105);
   U27560 : BUF_X1 port map( A => n40102, Z => n40104);
   U27561 : BUF_X1 port map( A => n40102, Z => n40103);
   U27562 : BUF_X1 port map( A => n39985, Z => n39990);
   U27563 : BUF_X1 port map( A => n39985, Z => n39989);
   U27564 : BUF_X1 port map( A => n39985, Z => n39988);
   U27565 : BUF_X1 port map( A => n39985, Z => n39987);
   U27566 : BUF_X1 port map( A => n39985, Z => n39986);
   U27567 : BUF_X1 port map( A => n39965, Z => n39970);
   U27568 : BUF_X1 port map( A => n39965, Z => n39969);
   U27569 : BUF_X1 port map( A => n39965, Z => n39968);
   U27570 : BUF_X1 port map( A => n39965, Z => n39967);
   U27571 : BUF_X1 port map( A => n39965, Z => n39966);
   U27572 : BUF_X1 port map( A => n39945, Z => n39950);
   U27573 : BUF_X1 port map( A => n39945, Z => n39949);
   U27574 : BUF_X1 port map( A => n39945, Z => n39948);
   U27575 : BUF_X1 port map( A => n39945, Z => n39947);
   U27576 : BUF_X1 port map( A => n39945, Z => n39946);
   U27577 : BUF_X1 port map( A => n39867, Z => n39872);
   U27578 : BUF_X1 port map( A => n39867, Z => n39871);
   U27579 : BUF_X1 port map( A => n39867, Z => n39870);
   U27580 : BUF_X1 port map( A => n39867, Z => n39869);
   U27581 : BUF_X1 port map( A => n39867, Z => n39868);
   U27582 : BUF_X1 port map( A => n39847, Z => n39852);
   U27583 : BUF_X1 port map( A => n39847, Z => n39851);
   U27584 : BUF_X1 port map( A => n39847, Z => n39850);
   U27585 : BUF_X1 port map( A => n39847, Z => n39849);
   U27586 : BUF_X1 port map( A => n39847, Z => n39848);
   U27587 : BUF_X1 port map( A => n39807, Z => n39812);
   U27588 : BUF_X1 port map( A => n39807, Z => n39811);
   U27589 : BUF_X1 port map( A => n33391, Z => n39952);
   U27590 : BUF_X1 port map( A => n33406, Z => n39894);
   U27591 : BUF_X1 port map( A => n33403, Z => n39913);
   U27592 : BUF_X1 port map( A => n33399, Z => n39932);
   U27593 : AND2_X1 port map( A1 => n37228, A2 => n37246, ZN => n36016);
   U27594 : BUF_X1 port map( A => n35981, Z => n39289);
   U27595 : BUF_X1 port map( A => n35981, Z => n39290);
   U27596 : BUF_X1 port map( A => n35981, Z => n39291);
   U27597 : BUF_X1 port map( A => n35981, Z => n39288);
   U27598 : BUF_X1 port map( A => n35981, Z => n39292);
   U27599 : BUF_X1 port map( A => n33426, Z => n39794);
   U27600 : BUF_X1 port map( A => n34700, Z => n39542);
   U27601 : BUF_X1 port map( A => n33426, Z => n39793);
   U27602 : BUF_X1 port map( A => n34700, Z => n39541);
   U27603 : BUF_X1 port map( A => n33426, Z => n39792);
   U27604 : BUF_X1 port map( A => n34700, Z => n39540);
   U27605 : BUF_X1 port map( A => n33426, Z => n39791);
   U27606 : BUF_X1 port map( A => n34700, Z => n39539);
   U27607 : BUF_X1 port map( A => n33426, Z => n39790);
   U27608 : BUF_X1 port map( A => n34700, Z => n39538);
   U27609 : OAI221_X1 port map( B1 => n33264, B2 => n33307, C1 => n33265, C2 =>
                           n33308, A => n41366, ZN => n33311);
   U27610 : OAI221_X1 port map( B1 => n33274, B2 => n33339, C1 => n33275, C2 =>
                           n33340, A => n41366, ZN => n33349);
   U27611 : OAI221_X1 port map( B1 => n33274, B2 => n33307, C1 => n33275, C2 =>
                           n33308, A => n41366, ZN => n33317);
   U27612 : OAI221_X1 port map( B1 => n33264, B2 => n33339, C1 => n33265, C2 =>
                           n33340, A => n41366, ZN => n33343);
   U27613 : OAI221_X1 port map( B1 => n33264, B2 => n33368, C1 => n33265, C2 =>
                           n33369, A => n41366, ZN => n33372);
   U27614 : OAI221_X1 port map( B1 => n33274, B2 => n33368, C1 => n33275, C2 =>
                           n33369, A => n41365, ZN => n33378);
   U27615 : OAI221_X1 port map( B1 => n33269, B2 => n33339, C1 => n33270, C2 =>
                           n33340, A => n41366, ZN => n33346);
   U27616 : OAI221_X1 port map( B1 => n33269, B2 => n33307, C1 => n33270, C2 =>
                           n33308, A => n41366, ZN => n33314);
   U27617 : OAI221_X1 port map( B1 => n33269, B2 => n33368, C1 => n33270, C2 =>
                           n33369, A => n41364, ZN => n33375);
   U27618 : OAI221_X1 port map( B1 => n33270, B2 => n33396, C1 => n33269, C2 =>
                           n33397, A => n41365, ZN => n33405);
   U27619 : OAI221_X1 port map( B1 => n33265, B2 => n33396, C1 => n33264, C2 =>
                           n33397, A => n41365, ZN => n33401);
   U27620 : OAI221_X1 port map( B1 => n33290, B2 => n33396, C1 => n32159, C2 =>
                           n33397, A => n41364, ZN => n33417);
   U27621 : OAI221_X1 port map( B1 => n33260, B2 => n33396, C1 => n33255, C2 =>
                           n33397, A => n41365, ZN => n33393);
   U27622 : OAI221_X1 port map( B1 => n33275, B2 => n33396, C1 => n33274, C2 =>
                           n33397, A => n41364, ZN => n33408);
   U27623 : OAI221_X1 port map( B1 => n33280, B2 => n33396, C1 => n32157, C2 =>
                           n33397, A => n41364, ZN => n33411);
   U27624 : OAI221_X1 port map( B1 => n33285, B2 => n33396, C1 => n32158, C2 =>
                           n33397, A => n41364, ZN => n33414);
   U27625 : OAI221_X1 port map( B1 => n33255, B2 => n33307, C1 => n33260, C2 =>
                           n33308, A => n41365, ZN => n33304);
   U27626 : OAI221_X1 port map( B1 => n32158, B2 => n33368, C1 => n33285, C2 =>
                           n33369, A => n41365, ZN => n33384);
   U27627 : OAI221_X1 port map( B1 => n32157, B2 => n33368, C1 => n33280, C2 =>
                           n33369, A => n41365, ZN => n33381);
   U27628 : OAI221_X1 port map( B1 => n32159, B2 => n33307, C1 => n33290, C2 =>
                           n33308, A => n41367, ZN => n33326);
   U27629 : OAI221_X1 port map( B1 => n32158, B2 => n33307, C1 => n33285, C2 =>
                           n33308, A => n41366, ZN => n33323);
   U27630 : OAI221_X1 port map( B1 => n32157, B2 => n33307, C1 => n33280, C2 =>
                           n33308, A => n41367, ZN => n33320);
   U27631 : OAI221_X1 port map( B1 => n32160, B2 => n33307, C1 => n33296, C2 =>
                           n33308, A => n41365, ZN => n33329);
   U27632 : OAI221_X1 port map( B1 => n33255, B2 => n33339, C1 => n33260, C2 =>
                           n33340, A => n41367, ZN => n33336);
   U27633 : OAI221_X1 port map( B1 => n32157, B2 => n33339, C1 => n33280, C2 =>
                           n33340, A => n41366, ZN => n33352);
   U27634 : OAI221_X1 port map( B1 => n32158, B2 => n33339, C1 => n33285, C2 =>
                           n33340, A => n41366, ZN => n33355);
   U27635 : OAI221_X1 port map( B1 => n32159, B2 => n33339, C1 => n33290, C2 =>
                           n33340, A => n41366, ZN => n33358);
   U27636 : OAI221_X1 port map( B1 => n32160, B2 => n33339, C1 => n33296, C2 =>
                           n33340, A => n41366, ZN => n33361);
   U27637 : OAI221_X1 port map( B1 => n33255, B2 => n33368, C1 => n33260, C2 =>
                           n33369, A => n41366, ZN => n33365);
   U27638 : OAI221_X1 port map( B1 => n32159, B2 => n33368, C1 => n33290, C2 =>
                           n33369, A => n41365, ZN => n33387);
   U27639 : OAI221_X1 port map( B1 => n32160, B2 => n33368, C1 => n33296, C2 =>
                           n33369, A => n41365, ZN => n33390);
   U27640 : OAI221_X1 port map( B1 => n32160, B2 => n33397, C1 => n33296, C2 =>
                           n33396, A => n41364, ZN => n33420);
   U27641 : NOR3_X1 port map( A1 => n32251, A2 => n32254, A3 => n32248, ZN => 
                           n37228);
   U27642 : NOR2_X1 port map( A1 => n32246, A2 => n32243, ZN => n37246);
   U27643 : NOR3_X1 port map( A1 => n32168, A2 => n32166, A3 => n32165, ZN => 
                           n34674);
   U27644 : NOR3_X1 port map( A1 => n32173, A2 => n32171, A3 => n32170, ZN => 
                           n35948);
   U27645 : INV_X1 port map( A => n33295, ZN => n32160);
   U27646 : INV_X1 port map( A => n33289, ZN => n32159);
   U27647 : INV_X1 port map( A => n33279, ZN => n32157);
   U27648 : INV_X1 port map( A => n33284, ZN => n32158);
   U27649 : NAND2_X1 port map( A1 => n33333, A2 => n33294, ZN => n33397);
   U27650 : INV_X1 port map( A => n33264, ZN => n32154);
   U27651 : INV_X1 port map( A => n33274, ZN => n32156);
   U27652 : INV_X1 port map( A => n33269, ZN => n32155);
   U27653 : NAND2_X1 port map( A1 => n37249, A2 => n37228, ZN => n36033);
   U27654 : NAND2_X1 port map( A1 => n37249, A2 => n37234, ZN => n36039);
   U27655 : NAND2_X1 port map( A1 => n37249, A2 => n37230, ZN => n36038);
   U27656 : NAND2_X1 port map( A1 => n37249, A2 => n37231, ZN => n36037);
   U27657 : NAND2_X1 port map( A1 => n34693, A2 => n34673, ZN => n33478);
   U27658 : NAND2_X1 port map( A1 => n34693, A2 => n34679, ZN => n33484);
   U27659 : NAND2_X1 port map( A1 => n34693, A2 => n34675, ZN => n33483);
   U27660 : NAND2_X1 port map( A1 => n34693, A2 => n34676, ZN => n33482);
   U27661 : NAND2_X1 port map( A1 => n35967, A2 => n35947, ZN => n34752);
   U27662 : NAND2_X1 port map( A1 => n35967, A2 => n35953, ZN => n34758);
   U27663 : NAND2_X1 port map( A1 => n35967, A2 => n35949, ZN => n34757);
   U27664 : NAND2_X1 port map( A1 => n35967, A2 => n35950, ZN => n34756);
   U27665 : BUF_X1 port map( A => n33273, Z => n40517);
   U27666 : BUF_X1 port map( A => n33273, Z => n40518);
   U27667 : BUF_X1 port map( A => n33273, Z => n40519);
   U27668 : BUF_X1 port map( A => n33273, Z => n40520);
   U27669 : BUF_X1 port map( A => n33273, Z => n40516);
   U27670 : BUF_X1 port map( A => n33263, Z => n40556);
   U27671 : BUF_X1 port map( A => n33263, Z => n40557);
   U27672 : BUF_X1 port map( A => n33263, Z => n40558);
   U27673 : BUF_X1 port map( A => n33263, Z => n40559);
   U27674 : BUF_X1 port map( A => n33263, Z => n40560);
   U27675 : BUF_X1 port map( A => n33268, Z => n40536);
   U27676 : BUF_X1 port map( A => n33268, Z => n40537);
   U27677 : BUF_X1 port map( A => n33268, Z => n40538);
   U27678 : BUF_X1 port map( A => n33268, Z => n40539);
   U27679 : BUF_X1 port map( A => n33268, Z => n40540);
   U27680 : BUF_X1 port map( A => n33278, Z => n40497);
   U27681 : BUF_X1 port map( A => n33278, Z => n40498);
   U27682 : BUF_X1 port map( A => n33278, Z => n40499);
   U27683 : BUF_X1 port map( A => n33278, Z => n40500);
   U27684 : BUF_X1 port map( A => n33278, Z => n40496);
   U27685 : BUF_X1 port map( A => n33254, Z => n40579);
   U27686 : BUF_X1 port map( A => n33254, Z => n40580);
   U27687 : BUF_X1 port map( A => n33254, Z => n40576);
   U27688 : BUF_X1 port map( A => n33254, Z => n40578);
   U27689 : BUF_X1 port map( A => n33254, Z => n40577);
   U27690 : BUF_X1 port map( A => n33283, Z => n40476);
   U27691 : BUF_X1 port map( A => n33283, Z => n40477);
   U27692 : BUF_X1 port map( A => n33283, Z => n40478);
   U27693 : BUF_X1 port map( A => n33283, Z => n40479);
   U27694 : BUF_X1 port map( A => n33283, Z => n40480);
   U27695 : BUF_X1 port map( A => n33288, Z => n40456);
   U27696 : BUF_X1 port map( A => n33288, Z => n40457);
   U27697 : BUF_X1 port map( A => n33288, Z => n40458);
   U27698 : BUF_X1 port map( A => n33288, Z => n40459);
   U27699 : BUF_X1 port map( A => n33288, Z => n40460);
   U27700 : BUF_X1 port map( A => n33293, Z => n40436);
   U27701 : BUF_X1 port map( A => n33293, Z => n40437);
   U27702 : BUF_X1 port map( A => n33293, Z => n40438);
   U27703 : BUF_X1 port map( A => n33293, Z => n40439);
   U27704 : BUF_X1 port map( A => n33293, Z => n40440);
   U27705 : BUF_X1 port map( A => n40582, Z => n40585);
   U27706 : BUF_X1 port map( A => n40582, Z => n40584);
   U27707 : BUF_X1 port map( A => n40582, Z => n40587);
   U27708 : BUF_X1 port map( A => n40582, Z => n40586);
   U27709 : BUF_X1 port map( A => n40582, Z => n40583);
   U27710 : NAND2_X1 port map( A1 => n37226, A2 => n37227, ZN => n35993);
   U27711 : NAND2_X1 port map( A1 => n37226, A2 => n37228, ZN => n35992);
   U27712 : NAND2_X1 port map( A1 => n37226, A2 => n37229, ZN => n35991);
   U27713 : NAND2_X1 port map( A1 => n37226, A2 => n37233, ZN => n35999);
   U27714 : NAND2_X1 port map( A1 => n37226, A2 => n37234, ZN => n35998);
   U27715 : NAND2_X1 port map( A1 => n37226, A2 => n37235, ZN => n35997);
   U27716 : BUF_X1 port map( A => n40522, Z => n40523);
   U27717 : BUF_X1 port map( A => n40522, Z => n40527);
   U27718 : BUF_X1 port map( A => n40522, Z => n40526);
   U27719 : BUF_X1 port map( A => n40522, Z => n40525);
   U27720 : BUF_X1 port map( A => n40522, Z => n40524);
   U27721 : BUF_X1 port map( A => n40502, Z => n40503);
   U27722 : BUF_X1 port map( A => n40502, Z => n40507);
   U27723 : BUF_X1 port map( A => n40502, Z => n40506);
   U27724 : BUF_X1 port map( A => n40502, Z => n40505);
   U27725 : BUF_X1 port map( A => n40502, Z => n40504);
   U27726 : BUF_X1 port map( A => n40562, Z => n40567);
   U27727 : BUF_X1 port map( A => n40562, Z => n40566);
   U27728 : BUF_X1 port map( A => n40562, Z => n40565);
   U27729 : BUF_X1 port map( A => n40562, Z => n40564);
   U27730 : BUF_X1 port map( A => n40562, Z => n40563);
   U27731 : BUF_X1 port map( A => n40542, Z => n40547);
   U27732 : BUF_X1 port map( A => n40542, Z => n40546);
   U27733 : BUF_X1 port map( A => n40542, Z => n40545);
   U27734 : BUF_X1 port map( A => n40542, Z => n40544);
   U27735 : BUF_X1 port map( A => n40542, Z => n40543);
   U27736 : BUF_X1 port map( A => n40482, Z => n40487);
   U27737 : BUF_X1 port map( A => n40482, Z => n40486);
   U27738 : BUF_X1 port map( A => n40482, Z => n40485);
   U27739 : BUF_X1 port map( A => n40482, Z => n40484);
   U27740 : BUF_X1 port map( A => n40482, Z => n40483);
   U27741 : BUF_X1 port map( A => n40462, Z => n40467);
   U27742 : BUF_X1 port map( A => n40462, Z => n40466);
   U27743 : BUF_X1 port map( A => n40462, Z => n40465);
   U27744 : BUF_X1 port map( A => n40462, Z => n40464);
   U27745 : BUF_X1 port map( A => n40462, Z => n40463);
   U27746 : BUF_X1 port map( A => n40442, Z => n40447);
   U27747 : BUF_X1 port map( A => n40442, Z => n40446);
   U27748 : BUF_X1 port map( A => n40442, Z => n40445);
   U27749 : BUF_X1 port map( A => n40442, Z => n40444);
   U27750 : BUF_X1 port map( A => n40442, Z => n40443);
   U27751 : NAND2_X1 port map( A1 => n37235, A2 => n37239, ZN => n36021);
   U27752 : NAND2_X1 port map( A1 => n37234, A2 => n37239, ZN => n36019);
   U27753 : NAND2_X1 port map( A1 => n37228, A2 => n37239, ZN => n36009);
   U27754 : NAND2_X1 port map( A1 => n37233, A2 => n37246, ZN => n36031);
   U27755 : NAND2_X1 port map( A1 => n37230, A2 => n37246, ZN => n36027);
   U27756 : NAND2_X1 port map( A1 => n37227, A2 => n37246, ZN => n36025);
   U27757 : NAND2_X1 port map( A1 => n34675, A2 => n34690, ZN => n33472);
   U27758 : NAND2_X1 port map( A1 => n35949, A2 => n35964, ZN => n34746);
   U27759 : NAND2_X1 port map( A1 => n37229, A2 => n37246, ZN => n36026);
   U27760 : NAND2_X1 port map( A1 => n37229, A2 => n37239, ZN => n36011);
   U27761 : NAND2_X1 port map( A1 => n34680, A2 => n34684, ZN => n33466);
   U27762 : NAND2_X1 port map( A1 => n34679, A2 => n34684, ZN => n33464);
   U27763 : NAND2_X1 port map( A1 => n34679, A2 => n34672, ZN => n33443);
   U27764 : NAND2_X1 port map( A1 => n34680, A2 => n34672, ZN => n33442);
   U27765 : NAND2_X1 port map( A1 => n35954, A2 => n35958, ZN => n34740);
   U27766 : NAND2_X1 port map( A1 => n35953, A2 => n35958, ZN => n34738);
   U27767 : NAND2_X1 port map( A1 => n35953, A2 => n35946, ZN => n34717);
   U27768 : NAND2_X1 port map( A1 => n35954, A2 => n35946, ZN => n34716);
   U27769 : NAND2_X1 port map( A1 => n34678, A2 => n34690, ZN => n33476);
   U27770 : NAND2_X1 port map( A1 => n34671, A2 => n34690, ZN => n33470);
   U27771 : NAND2_X1 port map( A1 => n34671, A2 => n34672, ZN => n33438);
   U27772 : NAND2_X1 port map( A1 => n34673, A2 => n34672, ZN => n33437);
   U27773 : NAND2_X1 port map( A1 => n34678, A2 => n34672, ZN => n33444);
   U27774 : NAND2_X1 port map( A1 => n34673, A2 => n34684, ZN => n33454);
   U27775 : NAND2_X1 port map( A1 => n35952, A2 => n35964, ZN => n34750);
   U27776 : NAND2_X1 port map( A1 => n35945, A2 => n35964, ZN => n34744);
   U27777 : NAND2_X1 port map( A1 => n35945, A2 => n35946, ZN => n34712);
   U27778 : NAND2_X1 port map( A1 => n35947, A2 => n35946, ZN => n34711);
   U27779 : NAND2_X1 port map( A1 => n35952, A2 => n35946, ZN => n34718);
   U27780 : NAND2_X1 port map( A1 => n35947, A2 => n35958, ZN => n34728);
   U27781 : NAND2_X1 port map( A1 => n37239, A2 => n37231, ZN => n36020);
   U27782 : NAND2_X1 port map( A1 => n34690, A2 => n34680, ZN => n33477);
   U27783 : NAND2_X1 port map( A1 => n35964, A2 => n35954, ZN => n34751);
   U27784 : NAND2_X1 port map( A1 => n37246, A2 => n37235, ZN => n36032);
   U27785 : NAND2_X1 port map( A1 => n34674, A2 => n34690, ZN => n33471);
   U27786 : NAND2_X1 port map( A1 => n34674, A2 => n34672, ZN => n33436);
   U27787 : NAND2_X1 port map( A1 => n34674, A2 => n34684, ZN => n33456);
   U27788 : NAND2_X1 port map( A1 => n35948, A2 => n35964, ZN => n34745);
   U27789 : NAND2_X1 port map( A1 => n35948, A2 => n35946, ZN => n34710);
   U27790 : NAND2_X1 port map( A1 => n35948, A2 => n35958, ZN => n34730);
   U27791 : AND2_X1 port map( A1 => n33331, A2 => n33294, ZN => n33395);
   U27792 : INV_X1 port map( A => n33255, ZN => n32153);
   U27793 : NAND2_X1 port map( A1 => n37236, A2 => n37233, ZN => n36010);
   U27794 : NAND2_X1 port map( A1 => n37236, A2 => n37231, ZN => n36005);
   U27795 : NAND2_X1 port map( A1 => n37236, A2 => n37227, ZN => n36004);
   U27796 : NAND2_X1 port map( A1 => n37236, A2 => n37230, ZN => n36003);
   U27797 : NAND2_X1 port map( A1 => n34684, A2 => n34676, ZN => n33465);
   U27798 : NAND2_X1 port map( A1 => n34681, A2 => n34676, ZN => n33450);
   U27799 : NAND2_X1 port map( A1 => n35958, A2 => n35950, ZN => n34739);
   U27800 : NAND2_X1 port map( A1 => n35955, A2 => n35950, ZN => n34724);
   U27801 : NAND2_X1 port map( A1 => n34681, A2 => n34671, ZN => n33449);
   U27802 : NAND2_X1 port map( A1 => n35955, A2 => n35945, ZN => n34723);
   U27803 : NAND2_X1 port map( A1 => n34681, A2 => n34675, ZN => n33448);
   U27804 : NAND2_X1 port map( A1 => n35955, A2 => n35949, ZN => n34722);
   U27805 : NAND2_X1 port map( A1 => n34681, A2 => n34678, ZN => n33455);
   U27806 : NAND2_X1 port map( A1 => n35955, A2 => n35952, ZN => n34729);
   U27807 : BUF_X1 port map( A => n33310, Z => n40402);
   U27808 : OAI211_X1 port map( C1 => n33264, C2 => n33305, A => n40401, B => 
                           n41367, ZN => n33310);
   U27809 : BUF_X1 port map( A => n33400, Z => n39925);
   U27810 : OAI211_X1 port map( C1 => n33264, C2 => n33394, A => n39920, B => 
                           n41369, ZN => n33400);
   U27811 : BUF_X1 port map( A => n33348, Z => n40202);
   U27812 : OAI211_X1 port map( C1 => n33274, C2 => n33337, A => n40201, B => 
                           n41368, ZN => n33348);
   U27813 : BUF_X1 port map( A => n33316, Z => n40362);
   U27814 : OAI211_X1 port map( C1 => n33274, C2 => n33305, A => n40361, B => 
                           n41368, ZN => n33316);
   U27815 : BUF_X1 port map( A => n33342, Z => n40242);
   U27816 : OAI211_X1 port map( C1 => n33264, C2 => n33337, A => n40241, B => 
                           n41368, ZN => n33342);
   U27817 : BUF_X1 port map( A => n33371, Z => n40083);
   U27818 : OAI211_X1 port map( C1 => n33264, C2 => n33366, A => n40082, B => 
                           n41369, ZN => n33371);
   U27819 : BUF_X1 port map( A => n33377, Z => n40043);
   U27820 : OAI211_X1 port map( C1 => n33274, C2 => n33366, A => n40042, B => 
                           n41369, ZN => n33377);
   U27821 : BUF_X1 port map( A => n33407, Z => n39887);
   U27822 : OAI211_X1 port map( C1 => n33274, C2 => n33394, A => n39886, B => 
                           n41369, ZN => n33407);
   U27823 : BUF_X1 port map( A => n33404, Z => n39906);
   U27824 : OAI211_X1 port map( C1 => n33269, C2 => n33394, A => n39901, B => 
                           n41369, ZN => n33404);
   U27825 : BUF_X1 port map( A => n33345, Z => n40222);
   U27826 : OAI211_X1 port map( C1 => n33269, C2 => n33337, A => n40221, B => 
                           n41368, ZN => n33345);
   U27827 : BUF_X1 port map( A => n33313, Z => n40382);
   U27828 : OAI211_X1 port map( C1 => n33269, C2 => n33305, A => n40381, B => 
                           n41367, ZN => n33313);
   U27829 : BUF_X1 port map( A => n33374, Z => n40063);
   U27830 : OAI211_X1 port map( C1 => n33269, C2 => n33366, A => n40062, B => 
                           n41369, ZN => n33374);
   U27831 : BUF_X1 port map( A => n33303, Z => n40422);
   U27832 : OAI211_X1 port map( C1 => n33255, C2 => n33305, A => n40421, B => 
                           n41368, ZN => n33303);
   U27833 : BUF_X1 port map( A => n33383, Z => n40004);
   U27834 : OAI211_X1 port map( C1 => n32158, C2 => n33366, A => n39999, B => 
                           n41369, ZN => n33383);
   U27835 : BUF_X1 port map( A => n33380, Z => n40023);
   U27836 : OAI211_X1 port map( C1 => n32157, C2 => n33366, A => n40018, B => 
                           n41369, ZN => n33380);
   U27837 : BUF_X1 port map( A => n33325, Z => n40302);
   U27838 : OAI211_X1 port map( C1 => n32159, C2 => n33305, A => n40301, B => 
                           n41368, ZN => n33325);
   U27839 : BUF_X1 port map( A => n33322, Z => n40322);
   U27840 : OAI211_X1 port map( C1 => n32158, C2 => n33305, A => n40321, B => 
                           n41367, ZN => n33322);
   U27841 : BUF_X1 port map( A => n33319, Z => n40342);
   U27842 : OAI211_X1 port map( C1 => n32157, C2 => n33305, A => n40341, B => 
                           n41368, ZN => n33319);
   U27843 : BUF_X1 port map( A => n33328, Z => n40282);
   U27844 : OAI211_X1 port map( C1 => n32160, C2 => n33305, A => n40281, B => 
                           n41368, ZN => n33328);
   U27845 : BUF_X1 port map( A => n33335, Z => n40262);
   U27846 : OAI211_X1 port map( C1 => n33255, C2 => n33337, A => n40261, B => 
                           n41368, ZN => n33335);
   U27847 : BUF_X1 port map( A => n33351, Z => n40182);
   U27848 : OAI211_X1 port map( C1 => n32157, C2 => n33337, A => n40181, B => 
                           n41368, ZN => n33351);
   U27849 : BUF_X1 port map( A => n33354, Z => n40162);
   U27850 : OAI211_X1 port map( C1 => n32158, C2 => n33337, A => n40161, B => 
                           n41368, ZN => n33354);
   U27851 : BUF_X1 port map( A => n33357, Z => n40142);
   U27852 : OAI211_X1 port map( C1 => n32159, C2 => n33337, A => n40141, B => 
                           n41369, ZN => n33357);
   U27853 : BUF_X1 port map( A => n33360, Z => n40122);
   U27854 : OAI211_X1 port map( C1 => n32160, C2 => n33337, A => n40116, B => 
                           n41369, ZN => n33360);
   U27855 : BUF_X1 port map( A => n33364, Z => n40102);
   U27856 : OAI211_X1 port map( C1 => n33255, C2 => n33366, A => n40097, B => 
                           n41369, ZN => n33364);
   U27857 : BUF_X1 port map( A => n33386, Z => n39985);
   U27858 : OAI211_X1 port map( C1 => n32159, C2 => n33366, A => n39984, B => 
                           n41369, ZN => n33386);
   U27859 : BUF_X1 port map( A => n33389, Z => n39965);
   U27860 : OAI211_X1 port map( C1 => n32160, C2 => n33366, A => n39964, B => 
                           n41369, ZN => n33389);
   U27861 : BUF_X1 port map( A => n33392, Z => n39945);
   U27862 : OAI211_X1 port map( C1 => n33255, C2 => n33394, A => n39944, B => 
                           n41369, ZN => n33392);
   U27863 : BUF_X1 port map( A => n33416, Z => n39827);
   U27864 : OAI211_X1 port map( C1 => n32159, C2 => n33394, A => n39826, B => 
                           n41370, ZN => n33416);
   U27865 : BUF_X1 port map( A => n33410, Z => n39867);
   U27866 : OAI211_X1 port map( C1 => n32157, C2 => n33394, A => n39866, B => 
                           n41370, ZN => n33410);
   U27867 : BUF_X1 port map( A => n33413, Z => n39847);
   U27868 : OAI211_X1 port map( C1 => n32158, C2 => n33394, A => n39846, B => 
                           n41370, ZN => n33413);
   U27869 : BUF_X1 port map( A => n33419, Z => n39807);
   U27870 : OAI211_X1 port map( C1 => n32160, C2 => n33394, A => n39802, B => 
                           n41370, ZN => n33419);
   U27871 : BUF_X1 port map( A => n33302, Z => n40429);
   U27872 : BUF_X1 port map( A => n33309, Z => n40409);
   U27873 : BUF_X1 port map( A => n33347, Z => n40209);
   U27874 : BUF_X1 port map( A => n33344, Z => n40229);
   U27875 : BUF_X1 port map( A => n33324, Z => n40309);
   U27876 : BUF_X1 port map( A => n33321, Z => n40329);
   U27877 : BUF_X1 port map( A => n33415, Z => n39834);
   U27878 : BUF_X1 port map( A => n33271, Z => n40529);
   U27879 : BUF_X1 port map( A => n33276, Z => n40509);
   U27880 : BUF_X1 port map( A => n33252, Z => n40589);
   U27881 : BUF_X1 port map( A => n33261, Z => n40569);
   U27882 : BUF_X1 port map( A => n33266, Z => n40549);
   U27883 : BUF_X1 port map( A => n33281, Z => n40489);
   U27884 : BUF_X1 port map( A => n33286, Z => n40469);
   U27885 : BUF_X1 port map( A => n33291, Z => n40449);
   U27886 : BUF_X1 port map( A => n33312, Z => n40389);
   U27887 : BUF_X1 port map( A => n33315, Z => n40369);
   U27888 : BUF_X1 port map( A => n33318, Z => n40349);
   U27889 : BUF_X1 port map( A => n33327, Z => n40289);
   U27890 : BUF_X1 port map( A => n33334, Z => n40269);
   U27891 : BUF_X1 port map( A => n33341, Z => n40249);
   U27892 : BUF_X1 port map( A => n33350, Z => n40189);
   U27893 : BUF_X1 port map( A => n33353, Z => n40169);
   U27894 : BUF_X1 port map( A => n33356, Z => n40149);
   U27895 : BUF_X1 port map( A => n33370, Z => n40090);
   U27896 : BUF_X1 port map( A => n33373, Z => n40070);
   U27897 : BUF_X1 port map( A => n33376, Z => n40050);
   U27898 : BUF_X1 port map( A => n33385, Z => n39992);
   U27899 : BUF_X1 port map( A => n33388, Z => n39972);
   U27900 : BUF_X1 port map( A => n33409, Z => n39874);
   U27901 : BUF_X1 port map( A => n33412, Z => n39854);
   U27902 : BUF_X1 port map( A => n33379, Z => n40030);
   U27903 : BUF_X1 port map( A => n33382, Z => n40011);
   U27904 : BUF_X1 port map( A => n33359, Z => n40129);
   U27905 : BUF_X1 port map( A => n33363, Z => n40109);
   U27906 : BUF_X1 port map( A => n33418, Z => n39814);
   U27907 : AND2_X1 port map( A1 => n37249, A2 => n37227, ZN => n36028);
   U27908 : AND2_X1 port map( A1 => n37249, A2 => n37229, ZN => n36029);
   U27909 : AND2_X1 port map( A1 => n37249, A2 => n37233, ZN => n36034);
   U27910 : AND2_X1 port map( A1 => n37249, A2 => n37235, ZN => n36035);
   U27911 : AND2_X1 port map( A1 => n34693, A2 => n34671, ZN => n33473);
   U27912 : AND2_X1 port map( A1 => n34693, A2 => n34674, ZN => n33474);
   U27913 : AND2_X1 port map( A1 => n34693, A2 => n34678, ZN => n33479);
   U27914 : AND2_X1 port map( A1 => n34693, A2 => n34680, ZN => n33480);
   U27915 : AND2_X1 port map( A1 => n35967, A2 => n35945, ZN => n34747);
   U27916 : AND2_X1 port map( A1 => n35967, A2 => n35948, ZN => n34748);
   U27917 : AND2_X1 port map( A1 => n35967, A2 => n35952, ZN => n34753);
   U27918 : AND2_X1 port map( A1 => n35967, A2 => n35954, ZN => n34754);
   U27919 : AND2_X1 port map( A1 => n37226, A2 => n37231, ZN => n35988);
   U27920 : AND2_X1 port map( A1 => n37226, A2 => n37230, ZN => n35989);
   U27921 : AND2_X1 port map( A1 => n34676, A2 => n34672, ZN => n33433);
   U27922 : AND2_X1 port map( A1 => n35950, A2 => n35946, ZN => n34707);
   U27923 : AND2_X1 port map( A1 => n37233, A2 => n37239, ZN => n36017);
   U27924 : AND2_X1 port map( A1 => n37230, A2 => n37239, ZN => n36006);
   U27925 : AND2_X1 port map( A1 => n37227, A2 => n37239, ZN => n36007);
   U27926 : AND2_X1 port map( A1 => n34675, A2 => n34672, ZN => n33434);
   U27927 : AND2_X1 port map( A1 => n34675, A2 => n34684, ZN => n33451);
   U27928 : AND2_X1 port map( A1 => n35949, A2 => n35946, ZN => n34708);
   U27929 : AND2_X1 port map( A1 => n35949, A2 => n35958, ZN => n34725);
   U27930 : AND2_X1 port map( A1 => n34673, A2 => n34690, ZN => n33461);
   U27931 : AND2_X1 port map( A1 => n34678, A2 => n34684, ZN => n33462);
   U27932 : AND2_X1 port map( A1 => n34671, A2 => n34684, ZN => n33452);
   U27933 : AND2_X1 port map( A1 => n35947, A2 => n35964, ZN => n34735);
   U27934 : AND2_X1 port map( A1 => n35952, A2 => n35958, ZN => n34736);
   U27935 : AND2_X1 port map( A1 => n35945, A2 => n35958, ZN => n34726);
   U27936 : AND2_X1 port map( A1 => n37246, A2 => n37234, ZN => n36022);
   U27937 : AND2_X1 port map( A1 => n37246, A2 => n37231, ZN => n36023);
   U27938 : AND2_X1 port map( A1 => n34690, A2 => n34679, ZN => n33467);
   U27939 : AND2_X1 port map( A1 => n34690, A2 => n34676, ZN => n33468);
   U27940 : AND2_X1 port map( A1 => n35964, A2 => n35953, ZN => n34741);
   U27941 : AND2_X1 port map( A1 => n35964, A2 => n35950, ZN => n34742);
   U27942 : AND2_X1 port map( A1 => n37236, A2 => n37235, ZN => n36000);
   U27943 : AND2_X1 port map( A1 => n37236, A2 => n37234, ZN => n36001);
   U27944 : AND2_X1 port map( A1 => n37236, A2 => n37229, ZN => n35994);
   U27945 : AND2_X1 port map( A1 => n37236, A2 => n37228, ZN => n35995);
   U27946 : AND2_X1 port map( A1 => n34681, A2 => n34680, ZN => n33445);
   U27947 : AND2_X1 port map( A1 => n34681, A2 => n34679, ZN => n33446);
   U27948 : AND2_X1 port map( A1 => n35955, A2 => n35954, ZN => n34719);
   U27949 : AND2_X1 port map( A1 => n35955, A2 => n35953, ZN => n34720);
   U27950 : AND2_X1 port map( A1 => n34681, A2 => n34673, ZN => n33440);
   U27951 : AND2_X1 port map( A1 => n35955, A2 => n35947, ZN => n34714);
   U27952 : AND2_X1 port map( A1 => n34681, A2 => n34674, ZN => n33439);
   U27953 : AND2_X1 port map( A1 => n35955, A2 => n35948, ZN => n34713);
   U27954 : INV_X1 port map( A => n33301, ZN => n32150);
   U27955 : NAND2_X1 port map( A1 => n41370, A2 => n35972, ZN => n35981);
   U27956 : INV_X1 port map( A => n33225, ZN => n32075);
   U27957 : NAND2_X1 port map( A1 => n41370, A2 => n39796, ZN => n33426);
   U27958 : NAND2_X1 port map( A1 => n41370, A2 => n39544, ZN => n34700);
   U27959 : BUF_X1 port map( A => n40981, Z => n40984);
   U27960 : BUF_X1 port map( A => n40987, Z => n40990);
   U27961 : BUF_X1 port map( A => n40993, Z => n40996);
   U27962 : BUF_X1 port map( A => n40999, Z => n41002);
   U27963 : BUF_X1 port map( A => n41005, Z => n41008);
   U27964 : BUF_X1 port map( A => n41011, Z => n41014);
   U27965 : BUF_X1 port map( A => n41017, Z => n41020);
   U27966 : BUF_X1 port map( A => n41023, Z => n41026);
   U27967 : BUF_X1 port map( A => n41029, Z => n41032);
   U27968 : BUF_X1 port map( A => n41035, Z => n41038);
   U27969 : BUF_X1 port map( A => n41041, Z => n41044);
   U27970 : BUF_X1 port map( A => n41047, Z => n41050);
   U27971 : BUF_X1 port map( A => n41053, Z => n41056);
   U27972 : BUF_X1 port map( A => n41059, Z => n41062);
   U27973 : BUF_X1 port map( A => n41065, Z => n41068);
   U27974 : BUF_X1 port map( A => n41071, Z => n41074);
   U27975 : BUF_X1 port map( A => n41077, Z => n41080);
   U27976 : BUF_X1 port map( A => n41083, Z => n41086);
   U27977 : BUF_X1 port map( A => n41089, Z => n41092);
   U27978 : BUF_X1 port map( A => n41095, Z => n41098);
   U27979 : BUF_X1 port map( A => n41101, Z => n41104);
   U27980 : BUF_X1 port map( A => n41107, Z => n41110);
   U27981 : BUF_X1 port map( A => n41113, Z => n41116);
   U27982 : BUF_X1 port map( A => n41119, Z => n41122);
   U27983 : BUF_X1 port map( A => n41125, Z => n41128);
   U27984 : BUF_X1 port map( A => n41131, Z => n41134);
   U27985 : BUF_X1 port map( A => n41137, Z => n41140);
   U27986 : BUF_X1 port map( A => n41143, Z => n41146);
   U27987 : BUF_X1 port map( A => n41149, Z => n41152);
   U27988 : BUF_X1 port map( A => n41155, Z => n41158);
   U27989 : BUF_X1 port map( A => n41161, Z => n41164);
   U27990 : BUF_X1 port map( A => n41167, Z => n41170);
   U27991 : BUF_X1 port map( A => n41173, Z => n41176);
   U27992 : BUF_X1 port map( A => n41179, Z => n41182);
   U27993 : BUF_X1 port map( A => n41185, Z => n41188);
   U27994 : BUF_X1 port map( A => n41191, Z => n41194);
   U27995 : BUF_X1 port map( A => n41197, Z => n41200);
   U27996 : BUF_X1 port map( A => n41203, Z => n41206);
   U27997 : BUF_X1 port map( A => n41209, Z => n41212);
   U27998 : BUF_X1 port map( A => n41215, Z => n41218);
   U27999 : BUF_X1 port map( A => n41221, Z => n41224);
   U28000 : BUF_X1 port map( A => n41227, Z => n41230);
   U28001 : BUF_X1 port map( A => n41233, Z => n41236);
   U28002 : BUF_X1 port map( A => n41239, Z => n41242);
   U28003 : BUF_X1 port map( A => n41245, Z => n41248);
   U28004 : BUF_X1 port map( A => n41251, Z => n41254);
   U28005 : BUF_X1 port map( A => n41257, Z => n41260);
   U28006 : BUF_X1 port map( A => n41263, Z => n41266);
   U28007 : BUF_X1 port map( A => n41269, Z => n41272);
   U28008 : BUF_X1 port map( A => n41275, Z => n41278);
   U28009 : BUF_X1 port map( A => n41281, Z => n41284);
   U28010 : BUF_X1 port map( A => n41287, Z => n41290);
   U28011 : BUF_X1 port map( A => n41293, Z => n41296);
   U28012 : BUF_X1 port map( A => n41299, Z => n41302);
   U28013 : BUF_X1 port map( A => n41305, Z => n41308);
   U28014 : BUF_X1 port map( A => n41311, Z => n41314);
   U28015 : BUF_X1 port map( A => n41317, Z => n41320);
   U28016 : BUF_X1 port map( A => n41323, Z => n41326);
   U28017 : BUF_X1 port map( A => n41329, Z => n41332);
   U28018 : BUF_X1 port map( A => n41335, Z => n41338);
   U28019 : BUF_X1 port map( A => n41341, Z => n41344);
   U28020 : BUF_X1 port map( A => n41347, Z => n41350);
   U28021 : BUF_X1 port map( A => n41353, Z => n41356);
   U28022 : BUF_X1 port map( A => n41359, Z => n41362);
   U28023 : BUF_X1 port map( A => n40980, Z => n40983);
   U28024 : BUF_X1 port map( A => n40986, Z => n40989);
   U28025 : BUF_X1 port map( A => n40992, Z => n40995);
   U28026 : BUF_X1 port map( A => n40998, Z => n41001);
   U28027 : BUF_X1 port map( A => n41004, Z => n41007);
   U28028 : BUF_X1 port map( A => n41010, Z => n41013);
   U28029 : BUF_X1 port map( A => n41016, Z => n41019);
   U28030 : BUF_X1 port map( A => n41022, Z => n41025);
   U28031 : BUF_X1 port map( A => n41028, Z => n41031);
   U28032 : BUF_X1 port map( A => n41034, Z => n41037);
   U28033 : BUF_X1 port map( A => n41040, Z => n41043);
   U28034 : BUF_X1 port map( A => n41046, Z => n41049);
   U28035 : BUF_X1 port map( A => n41052, Z => n41055);
   U28036 : BUF_X1 port map( A => n41058, Z => n41061);
   U28037 : BUF_X1 port map( A => n41064, Z => n41067);
   U28038 : BUF_X1 port map( A => n41070, Z => n41073);
   U28039 : BUF_X1 port map( A => n41076, Z => n41079);
   U28040 : BUF_X1 port map( A => n41082, Z => n41085);
   U28041 : BUF_X1 port map( A => n41088, Z => n41091);
   U28042 : BUF_X1 port map( A => n41094, Z => n41097);
   U28043 : BUF_X1 port map( A => n41100, Z => n41103);
   U28044 : BUF_X1 port map( A => n41106, Z => n41109);
   U28045 : BUF_X1 port map( A => n41112, Z => n41115);
   U28046 : BUF_X1 port map( A => n41118, Z => n41121);
   U28047 : BUF_X1 port map( A => n41124, Z => n41127);
   U28048 : BUF_X1 port map( A => n41130, Z => n41133);
   U28049 : BUF_X1 port map( A => n41136, Z => n41139);
   U28050 : BUF_X1 port map( A => n41142, Z => n41145);
   U28051 : BUF_X1 port map( A => n41148, Z => n41151);
   U28052 : BUF_X1 port map( A => n41154, Z => n41157);
   U28053 : BUF_X1 port map( A => n41160, Z => n41163);
   U28054 : BUF_X1 port map( A => n41166, Z => n41169);
   U28055 : BUF_X1 port map( A => n41172, Z => n41175);
   U28056 : BUF_X1 port map( A => n41178, Z => n41181);
   U28057 : BUF_X1 port map( A => n41184, Z => n41187);
   U28058 : BUF_X1 port map( A => n41190, Z => n41193);
   U28059 : BUF_X1 port map( A => n41196, Z => n41199);
   U28060 : BUF_X1 port map( A => n41202, Z => n41205);
   U28061 : BUF_X1 port map( A => n41208, Z => n41211);
   U28062 : BUF_X1 port map( A => n41214, Z => n41217);
   U28063 : BUF_X1 port map( A => n41220, Z => n41223);
   U28064 : BUF_X1 port map( A => n41226, Z => n41229);
   U28065 : BUF_X1 port map( A => n41232, Z => n41235);
   U28066 : BUF_X1 port map( A => n41238, Z => n41241);
   U28067 : BUF_X1 port map( A => n41244, Z => n41247);
   U28068 : BUF_X1 port map( A => n41250, Z => n41253);
   U28069 : BUF_X1 port map( A => n41256, Z => n41259);
   U28070 : BUF_X1 port map( A => n41262, Z => n41265);
   U28071 : BUF_X1 port map( A => n41268, Z => n41271);
   U28072 : BUF_X1 port map( A => n41274, Z => n41277);
   U28073 : BUF_X1 port map( A => n41280, Z => n41283);
   U28074 : BUF_X1 port map( A => n41286, Z => n41289);
   U28075 : BUF_X1 port map( A => n41292, Z => n41295);
   U28076 : BUF_X1 port map( A => n41298, Z => n41301);
   U28077 : BUF_X1 port map( A => n41304, Z => n41307);
   U28078 : BUF_X1 port map( A => n41310, Z => n41313);
   U28079 : BUF_X1 port map( A => n41316, Z => n41319);
   U28080 : BUF_X1 port map( A => n41322, Z => n41325);
   U28081 : BUF_X1 port map( A => n41328, Z => n41331);
   U28082 : BUF_X1 port map( A => n41334, Z => n41337);
   U28083 : BUF_X1 port map( A => n41340, Z => n41343);
   U28084 : BUF_X1 port map( A => n41346, Z => n41349);
   U28085 : BUF_X1 port map( A => n41352, Z => n41355);
   U28086 : BUF_X1 port map( A => n41358, Z => n41361);
   U28087 : BUF_X1 port map( A => n41118, Z => n41120);
   U28088 : BUF_X1 port map( A => n41124, Z => n41126);
   U28089 : BUF_X1 port map( A => n41130, Z => n41132);
   U28090 : BUF_X1 port map( A => n41136, Z => n41138);
   U28091 : BUF_X1 port map( A => n41142, Z => n41144);
   U28092 : BUF_X1 port map( A => n41148, Z => n41150);
   U28093 : BUF_X1 port map( A => n41154, Z => n41156);
   U28094 : BUF_X1 port map( A => n41160, Z => n41162);
   U28095 : BUF_X1 port map( A => n41166, Z => n41168);
   U28096 : BUF_X1 port map( A => n41172, Z => n41174);
   U28097 : BUF_X1 port map( A => n41178, Z => n41180);
   U28098 : BUF_X1 port map( A => n41184, Z => n41186);
   U28099 : BUF_X1 port map( A => n41190, Z => n41192);
   U28100 : BUF_X1 port map( A => n41196, Z => n41198);
   U28101 : BUF_X1 port map( A => n41202, Z => n41204);
   U28102 : BUF_X1 port map( A => n41208, Z => n41210);
   U28103 : BUF_X1 port map( A => n41214, Z => n41216);
   U28104 : BUF_X1 port map( A => n41220, Z => n41222);
   U28105 : BUF_X1 port map( A => n41226, Z => n41228);
   U28106 : BUF_X1 port map( A => n41232, Z => n41234);
   U28107 : BUF_X1 port map( A => n41238, Z => n41240);
   U28108 : BUF_X1 port map( A => n41244, Z => n41246);
   U28109 : BUF_X1 port map( A => n41250, Z => n41252);
   U28110 : BUF_X1 port map( A => n41256, Z => n41258);
   U28111 : BUF_X1 port map( A => n41262, Z => n41264);
   U28112 : BUF_X1 port map( A => n41268, Z => n41270);
   U28113 : BUF_X1 port map( A => n41274, Z => n41276);
   U28114 : BUF_X1 port map( A => n41280, Z => n41282);
   U28115 : BUF_X1 port map( A => n41286, Z => n41288);
   U28116 : BUF_X1 port map( A => n41292, Z => n41294);
   U28117 : BUF_X1 port map( A => n41298, Z => n41300);
   U28118 : BUF_X1 port map( A => n41304, Z => n41306);
   U28119 : BUF_X1 port map( A => n41310, Z => n41312);
   U28120 : BUF_X1 port map( A => n41316, Z => n41318);
   U28121 : BUF_X1 port map( A => n41322, Z => n41324);
   U28122 : BUF_X1 port map( A => n41328, Z => n41330);
   U28123 : BUF_X1 port map( A => n41334, Z => n41336);
   U28124 : BUF_X1 port map( A => n41340, Z => n41342);
   U28125 : BUF_X1 port map( A => n41346, Z => n41348);
   U28126 : BUF_X1 port map( A => n41352, Z => n41354);
   U28127 : BUF_X1 port map( A => n41358, Z => n41360);
   U28128 : BUF_X1 port map( A => n40980, Z => n40982);
   U28129 : BUF_X1 port map( A => n40986, Z => n40988);
   U28130 : BUF_X1 port map( A => n40992, Z => n40994);
   U28131 : BUF_X1 port map( A => n40998, Z => n41000);
   U28132 : BUF_X1 port map( A => n41004, Z => n41006);
   U28133 : BUF_X1 port map( A => n41010, Z => n41012);
   U28134 : BUF_X1 port map( A => n41016, Z => n41018);
   U28135 : BUF_X1 port map( A => n41022, Z => n41024);
   U28136 : BUF_X1 port map( A => n41028, Z => n41030);
   U28137 : BUF_X1 port map( A => n41034, Z => n41036);
   U28138 : BUF_X1 port map( A => n41040, Z => n41042);
   U28139 : BUF_X1 port map( A => n41046, Z => n41048);
   U28140 : BUF_X1 port map( A => n41052, Z => n41054);
   U28141 : BUF_X1 port map( A => n41058, Z => n41060);
   U28142 : BUF_X1 port map( A => n41064, Z => n41066);
   U28143 : BUF_X1 port map( A => n41070, Z => n41072);
   U28144 : BUF_X1 port map( A => n41076, Z => n41078);
   U28145 : BUF_X1 port map( A => n41082, Z => n41084);
   U28146 : BUF_X1 port map( A => n41088, Z => n41090);
   U28147 : BUF_X1 port map( A => n41094, Z => n41096);
   U28148 : BUF_X1 port map( A => n41100, Z => n41102);
   U28149 : BUF_X1 port map( A => n41106, Z => n41108);
   U28150 : BUF_X1 port map( A => n41112, Z => n41114);
   U28151 : BUF_X1 port map( A => n40597, Z => n40600);
   U28152 : BUF_X1 port map( A => n40603, Z => n40606);
   U28153 : BUF_X1 port map( A => n40609, Z => n40612);
   U28154 : BUF_X1 port map( A => n40615, Z => n40618);
   U28155 : BUF_X1 port map( A => n40621, Z => n40624);
   U28156 : BUF_X1 port map( A => n40627, Z => n40630);
   U28157 : BUF_X1 port map( A => n40633, Z => n40636);
   U28158 : BUF_X1 port map( A => n40639, Z => n40642);
   U28159 : BUF_X1 port map( A => n40645, Z => n40648);
   U28160 : BUF_X1 port map( A => n40651, Z => n40654);
   U28161 : BUF_X1 port map( A => n40657, Z => n40660);
   U28162 : BUF_X1 port map( A => n40663, Z => n40666);
   U28163 : BUF_X1 port map( A => n40669, Z => n40672);
   U28164 : BUF_X1 port map( A => n40675, Z => n40678);
   U28165 : BUF_X1 port map( A => n40681, Z => n40684);
   U28166 : BUF_X1 port map( A => n40687, Z => n40690);
   U28167 : BUF_X1 port map( A => n40693, Z => n40696);
   U28168 : BUF_X1 port map( A => n40699, Z => n40702);
   U28169 : BUF_X1 port map( A => n40705, Z => n40708);
   U28170 : BUF_X1 port map( A => n40711, Z => n40714);
   U28171 : BUF_X1 port map( A => n40717, Z => n40720);
   U28172 : BUF_X1 port map( A => n40723, Z => n40726);
   U28173 : BUF_X1 port map( A => n40729, Z => n40732);
   U28174 : BUF_X1 port map( A => n40735, Z => n40738);
   U28175 : BUF_X1 port map( A => n40741, Z => n40744);
   U28176 : BUF_X1 port map( A => n40747, Z => n40750);
   U28177 : BUF_X1 port map( A => n40753, Z => n40756);
   U28178 : BUF_X1 port map( A => n40759, Z => n40762);
   U28179 : BUF_X1 port map( A => n40765, Z => n40768);
   U28180 : BUF_X1 port map( A => n40771, Z => n40774);
   U28181 : BUF_X1 port map( A => n40777, Z => n40780);
   U28182 : BUF_X1 port map( A => n40783, Z => n40786);
   U28183 : BUF_X1 port map( A => n40789, Z => n40792);
   U28184 : BUF_X1 port map( A => n40795, Z => n40798);
   U28185 : BUF_X1 port map( A => n40801, Z => n40804);
   U28186 : BUF_X1 port map( A => n40807, Z => n40810);
   U28187 : BUF_X1 port map( A => n40813, Z => n40816);
   U28188 : BUF_X1 port map( A => n40819, Z => n40822);
   U28189 : BUF_X1 port map( A => n40825, Z => n40828);
   U28190 : BUF_X1 port map( A => n40831, Z => n40834);
   U28191 : BUF_X1 port map( A => n40837, Z => n40840);
   U28192 : BUF_X1 port map( A => n40843, Z => n40846);
   U28193 : BUF_X1 port map( A => n40849, Z => n40852);
   U28194 : BUF_X1 port map( A => n40855, Z => n40858);
   U28195 : BUF_X1 port map( A => n40861, Z => n40864);
   U28196 : BUF_X1 port map( A => n40867, Z => n40870);
   U28197 : BUF_X1 port map( A => n40873, Z => n40876);
   U28198 : BUF_X1 port map( A => n40879, Z => n40882);
   U28199 : BUF_X1 port map( A => n40885, Z => n40888);
   U28200 : BUF_X1 port map( A => n40891, Z => n40894);
   U28201 : BUF_X1 port map( A => n40897, Z => n40900);
   U28202 : BUF_X1 port map( A => n40903, Z => n40906);
   U28203 : BUF_X1 port map( A => n40909, Z => n40912);
   U28204 : BUF_X1 port map( A => n40915, Z => n40918);
   U28205 : BUF_X1 port map( A => n40921, Z => n40924);
   U28206 : BUF_X1 port map( A => n40927, Z => n40930);
   U28207 : BUF_X1 port map( A => n40933, Z => n40936);
   U28208 : BUF_X1 port map( A => n40939, Z => n40942);
   U28209 : BUF_X1 port map( A => n40945, Z => n40948);
   U28210 : BUF_X1 port map( A => n40951, Z => n40954);
   U28211 : BUF_X1 port map( A => n40957, Z => n40960);
   U28212 : BUF_X1 port map( A => n40963, Z => n40966);
   U28213 : BUF_X1 port map( A => n40969, Z => n40972);
   U28214 : BUF_X1 port map( A => n40975, Z => n40978);
   U28215 : BUF_X1 port map( A => n40596, Z => n40599);
   U28216 : BUF_X1 port map( A => n40602, Z => n40605);
   U28217 : BUF_X1 port map( A => n40608, Z => n40611);
   U28218 : BUF_X1 port map( A => n40614, Z => n40617);
   U28219 : BUF_X1 port map( A => n40620, Z => n40623);
   U28220 : BUF_X1 port map( A => n40626, Z => n40629);
   U28221 : BUF_X1 port map( A => n40632, Z => n40635);
   U28222 : BUF_X1 port map( A => n40638, Z => n40641);
   U28223 : BUF_X1 port map( A => n40644, Z => n40647);
   U28224 : BUF_X1 port map( A => n40650, Z => n40653);
   U28225 : BUF_X1 port map( A => n40656, Z => n40659);
   U28226 : BUF_X1 port map( A => n40662, Z => n40665);
   U28227 : BUF_X1 port map( A => n40668, Z => n40671);
   U28228 : BUF_X1 port map( A => n40674, Z => n40677);
   U28229 : BUF_X1 port map( A => n40680, Z => n40683);
   U28230 : BUF_X1 port map( A => n40686, Z => n40689);
   U28231 : BUF_X1 port map( A => n40692, Z => n40695);
   U28232 : BUF_X1 port map( A => n40698, Z => n40701);
   U28233 : BUF_X1 port map( A => n40704, Z => n40707);
   U28234 : BUF_X1 port map( A => n40710, Z => n40713);
   U28235 : BUF_X1 port map( A => n40716, Z => n40719);
   U28236 : BUF_X1 port map( A => n40722, Z => n40725);
   U28237 : BUF_X1 port map( A => n40728, Z => n40731);
   U28238 : BUF_X1 port map( A => n40734, Z => n40737);
   U28239 : BUF_X1 port map( A => n40740, Z => n40743);
   U28240 : BUF_X1 port map( A => n40746, Z => n40749);
   U28241 : BUF_X1 port map( A => n40752, Z => n40755);
   U28242 : BUF_X1 port map( A => n40758, Z => n40761);
   U28243 : BUF_X1 port map( A => n40764, Z => n40767);
   U28244 : BUF_X1 port map( A => n40770, Z => n40773);
   U28245 : BUF_X1 port map( A => n40776, Z => n40779);
   U28246 : BUF_X1 port map( A => n40782, Z => n40785);
   U28247 : BUF_X1 port map( A => n40788, Z => n40791);
   U28248 : BUF_X1 port map( A => n40794, Z => n40797);
   U28249 : BUF_X1 port map( A => n40800, Z => n40803);
   U28250 : BUF_X1 port map( A => n40806, Z => n40809);
   U28251 : BUF_X1 port map( A => n40812, Z => n40815);
   U28252 : BUF_X1 port map( A => n40818, Z => n40821);
   U28253 : BUF_X1 port map( A => n40824, Z => n40827);
   U28254 : BUF_X1 port map( A => n40830, Z => n40833);
   U28255 : BUF_X1 port map( A => n40836, Z => n40839);
   U28256 : BUF_X1 port map( A => n40842, Z => n40845);
   U28257 : BUF_X1 port map( A => n40848, Z => n40851);
   U28258 : BUF_X1 port map( A => n40854, Z => n40857);
   U28259 : BUF_X1 port map( A => n40860, Z => n40863);
   U28260 : BUF_X1 port map( A => n40866, Z => n40869);
   U28261 : BUF_X1 port map( A => n40872, Z => n40875);
   U28262 : BUF_X1 port map( A => n40878, Z => n40881);
   U28263 : BUF_X1 port map( A => n40884, Z => n40887);
   U28264 : BUF_X1 port map( A => n40890, Z => n40893);
   U28265 : BUF_X1 port map( A => n40896, Z => n40899);
   U28266 : BUF_X1 port map( A => n40902, Z => n40905);
   U28267 : BUF_X1 port map( A => n40908, Z => n40911);
   U28268 : BUF_X1 port map( A => n40914, Z => n40917);
   U28269 : BUF_X1 port map( A => n40920, Z => n40923);
   U28270 : BUF_X1 port map( A => n40926, Z => n40929);
   U28271 : BUF_X1 port map( A => n40932, Z => n40935);
   U28272 : BUF_X1 port map( A => n40938, Z => n40941);
   U28273 : BUF_X1 port map( A => n40944, Z => n40947);
   U28274 : BUF_X1 port map( A => n40950, Z => n40953);
   U28275 : BUF_X1 port map( A => n40956, Z => n40959);
   U28276 : BUF_X1 port map( A => n40962, Z => n40965);
   U28277 : BUF_X1 port map( A => n40968, Z => n40971);
   U28278 : BUF_X1 port map( A => n40974, Z => n40977);
   U28279 : BUF_X1 port map( A => n40734, Z => n40736);
   U28280 : BUF_X1 port map( A => n40740, Z => n40742);
   U28281 : BUF_X1 port map( A => n40746, Z => n40748);
   U28282 : BUF_X1 port map( A => n40752, Z => n40754);
   U28283 : BUF_X1 port map( A => n40758, Z => n40760);
   U28284 : BUF_X1 port map( A => n40764, Z => n40766);
   U28285 : BUF_X1 port map( A => n40770, Z => n40772);
   U28286 : BUF_X1 port map( A => n40776, Z => n40778);
   U28287 : BUF_X1 port map( A => n40782, Z => n40784);
   U28288 : BUF_X1 port map( A => n40788, Z => n40790);
   U28289 : BUF_X1 port map( A => n40794, Z => n40796);
   U28290 : BUF_X1 port map( A => n40800, Z => n40802);
   U28291 : BUF_X1 port map( A => n40806, Z => n40808);
   U28292 : BUF_X1 port map( A => n40812, Z => n40814);
   U28293 : BUF_X1 port map( A => n40818, Z => n40820);
   U28294 : BUF_X1 port map( A => n40824, Z => n40826);
   U28295 : BUF_X1 port map( A => n40830, Z => n40832);
   U28296 : BUF_X1 port map( A => n40836, Z => n40838);
   U28297 : BUF_X1 port map( A => n40842, Z => n40844);
   U28298 : BUF_X1 port map( A => n40848, Z => n40850);
   U28299 : BUF_X1 port map( A => n40854, Z => n40856);
   U28300 : BUF_X1 port map( A => n40860, Z => n40862);
   U28301 : BUF_X1 port map( A => n40866, Z => n40868);
   U28302 : BUF_X1 port map( A => n40872, Z => n40874);
   U28303 : BUF_X1 port map( A => n40878, Z => n40880);
   U28304 : BUF_X1 port map( A => n40884, Z => n40886);
   U28305 : BUF_X1 port map( A => n40890, Z => n40892);
   U28306 : BUF_X1 port map( A => n40896, Z => n40898);
   U28307 : BUF_X1 port map( A => n40902, Z => n40904);
   U28308 : BUF_X1 port map( A => n40908, Z => n40910);
   U28309 : BUF_X1 port map( A => n40914, Z => n40916);
   U28310 : BUF_X1 port map( A => n40920, Z => n40922);
   U28311 : BUF_X1 port map( A => n40926, Z => n40928);
   U28312 : BUF_X1 port map( A => n40932, Z => n40934);
   U28313 : BUF_X1 port map( A => n40938, Z => n40940);
   U28314 : BUF_X1 port map( A => n40944, Z => n40946);
   U28315 : BUF_X1 port map( A => n40950, Z => n40952);
   U28316 : BUF_X1 port map( A => n40956, Z => n40958);
   U28317 : BUF_X1 port map( A => n40962, Z => n40964);
   U28318 : BUF_X1 port map( A => n40968, Z => n40970);
   U28319 : BUF_X1 port map( A => n40974, Z => n40976);
   U28320 : BUF_X1 port map( A => n40596, Z => n40598);
   U28321 : BUF_X1 port map( A => n40602, Z => n40604);
   U28322 : BUF_X1 port map( A => n40608, Z => n40610);
   U28323 : BUF_X1 port map( A => n40614, Z => n40616);
   U28324 : BUF_X1 port map( A => n40620, Z => n40622);
   U28325 : BUF_X1 port map( A => n40626, Z => n40628);
   U28326 : BUF_X1 port map( A => n40632, Z => n40634);
   U28327 : BUF_X1 port map( A => n40638, Z => n40640);
   U28328 : BUF_X1 port map( A => n40644, Z => n40646);
   U28329 : BUF_X1 port map( A => n40650, Z => n40652);
   U28330 : BUF_X1 port map( A => n40656, Z => n40658);
   U28331 : BUF_X1 port map( A => n40662, Z => n40664);
   U28332 : BUF_X1 port map( A => n40668, Z => n40670);
   U28333 : BUF_X1 port map( A => n40674, Z => n40676);
   U28334 : BUF_X1 port map( A => n40680, Z => n40682);
   U28335 : BUF_X1 port map( A => n40686, Z => n40688);
   U28336 : BUF_X1 port map( A => n40692, Z => n40694);
   U28337 : BUF_X1 port map( A => n40698, Z => n40700);
   U28338 : BUF_X1 port map( A => n40704, Z => n40706);
   U28339 : BUF_X1 port map( A => n40710, Z => n40712);
   U28340 : BUF_X1 port map( A => n40716, Z => n40718);
   U28341 : BUF_X1 port map( A => n40722, Z => n40724);
   U28342 : BUF_X1 port map( A => n40728, Z => n40730);
   U28343 : BUF_X1 port map( A => n40981, Z => n40985);
   U28344 : BUF_X1 port map( A => n40987, Z => n40991);
   U28345 : BUF_X1 port map( A => n40993, Z => n40997);
   U28346 : BUF_X1 port map( A => n40999, Z => n41003);
   U28347 : BUF_X1 port map( A => n41005, Z => n41009);
   U28348 : BUF_X1 port map( A => n41011, Z => n41015);
   U28349 : BUF_X1 port map( A => n41017, Z => n41021);
   U28350 : BUF_X1 port map( A => n41023, Z => n41027);
   U28351 : BUF_X1 port map( A => n41029, Z => n41033);
   U28352 : BUF_X1 port map( A => n41035, Z => n41039);
   U28353 : BUF_X1 port map( A => n41041, Z => n41045);
   U28354 : BUF_X1 port map( A => n41047, Z => n41051);
   U28355 : BUF_X1 port map( A => n41053, Z => n41057);
   U28356 : BUF_X1 port map( A => n41059, Z => n41063);
   U28357 : BUF_X1 port map( A => n41065, Z => n41069);
   U28358 : BUF_X1 port map( A => n41071, Z => n41075);
   U28359 : BUF_X1 port map( A => n41077, Z => n41081);
   U28360 : BUF_X1 port map( A => n41083, Z => n41087);
   U28361 : BUF_X1 port map( A => n41089, Z => n41093);
   U28362 : BUF_X1 port map( A => n41095, Z => n41099);
   U28363 : BUF_X1 port map( A => n41101, Z => n41105);
   U28364 : BUF_X1 port map( A => n41107, Z => n41111);
   U28365 : BUF_X1 port map( A => n41113, Z => n41117);
   U28366 : BUF_X1 port map( A => n41119, Z => n41123);
   U28367 : BUF_X1 port map( A => n41125, Z => n41129);
   U28368 : BUF_X1 port map( A => n41131, Z => n41135);
   U28369 : BUF_X1 port map( A => n41137, Z => n41141);
   U28370 : BUF_X1 port map( A => n41143, Z => n41147);
   U28371 : BUF_X1 port map( A => n41149, Z => n41153);
   U28372 : BUF_X1 port map( A => n41155, Z => n41159);
   U28373 : BUF_X1 port map( A => n41161, Z => n41165);
   U28374 : BUF_X1 port map( A => n41167, Z => n41171);
   U28375 : BUF_X1 port map( A => n41173, Z => n41177);
   U28376 : BUF_X1 port map( A => n41179, Z => n41183);
   U28377 : BUF_X1 port map( A => n41185, Z => n41189);
   U28378 : BUF_X1 port map( A => n41191, Z => n41195);
   U28379 : BUF_X1 port map( A => n41197, Z => n41201);
   U28380 : BUF_X1 port map( A => n41203, Z => n41207);
   U28381 : BUF_X1 port map( A => n41209, Z => n41213);
   U28382 : BUF_X1 port map( A => n41215, Z => n41219);
   U28383 : BUF_X1 port map( A => n41221, Z => n41225);
   U28384 : BUF_X1 port map( A => n41227, Z => n41231);
   U28385 : BUF_X1 port map( A => n41233, Z => n41237);
   U28386 : BUF_X1 port map( A => n41239, Z => n41243);
   U28387 : BUF_X1 port map( A => n41245, Z => n41249);
   U28388 : BUF_X1 port map( A => n41251, Z => n41255);
   U28389 : BUF_X1 port map( A => n41257, Z => n41261);
   U28390 : BUF_X1 port map( A => n41263, Z => n41267);
   U28391 : BUF_X1 port map( A => n41269, Z => n41273);
   U28392 : BUF_X1 port map( A => n41275, Z => n41279);
   U28393 : BUF_X1 port map( A => n41281, Z => n41285);
   U28394 : BUF_X1 port map( A => n41287, Z => n41291);
   U28395 : BUF_X1 port map( A => n41293, Z => n41297);
   U28396 : BUF_X1 port map( A => n41299, Z => n41303);
   U28397 : BUF_X1 port map( A => n41305, Z => n41309);
   U28398 : BUF_X1 port map( A => n41311, Z => n41315);
   U28399 : BUF_X1 port map( A => n41317, Z => n41321);
   U28400 : BUF_X1 port map( A => n41323, Z => n41327);
   U28401 : BUF_X1 port map( A => n41329, Z => n41333);
   U28402 : BUF_X1 port map( A => n41335, Z => n41339);
   U28403 : BUF_X1 port map( A => n41341, Z => n41345);
   U28404 : BUF_X1 port map( A => n41347, Z => n41351);
   U28405 : BUF_X1 port map( A => n41353, Z => n41357);
   U28406 : BUF_X1 port map( A => n41359, Z => n41363);
   U28407 : BUF_X1 port map( A => n40597, Z => n40601);
   U28408 : BUF_X1 port map( A => n40603, Z => n40607);
   U28409 : BUF_X1 port map( A => n40609, Z => n40613);
   U28410 : BUF_X1 port map( A => n40615, Z => n40619);
   U28411 : BUF_X1 port map( A => n40621, Z => n40625);
   U28412 : BUF_X1 port map( A => n40627, Z => n40631);
   U28413 : BUF_X1 port map( A => n40633, Z => n40637);
   U28414 : BUF_X1 port map( A => n40639, Z => n40643);
   U28415 : BUF_X1 port map( A => n40645, Z => n40649);
   U28416 : BUF_X1 port map( A => n40651, Z => n40655);
   U28417 : BUF_X1 port map( A => n40657, Z => n40661);
   U28418 : BUF_X1 port map( A => n40663, Z => n40667);
   U28419 : BUF_X1 port map( A => n40669, Z => n40673);
   U28420 : BUF_X1 port map( A => n40675, Z => n40679);
   U28421 : BUF_X1 port map( A => n40681, Z => n40685);
   U28422 : BUF_X1 port map( A => n40687, Z => n40691);
   U28423 : BUF_X1 port map( A => n40693, Z => n40697);
   U28424 : BUF_X1 port map( A => n40699, Z => n40703);
   U28425 : BUF_X1 port map( A => n40705, Z => n40709);
   U28426 : BUF_X1 port map( A => n40711, Z => n40715);
   U28427 : BUF_X1 port map( A => n40717, Z => n40721);
   U28428 : BUF_X1 port map( A => n40723, Z => n40727);
   U28429 : BUF_X1 port map( A => n40729, Z => n40733);
   U28430 : BUF_X1 port map( A => n40735, Z => n40739);
   U28431 : BUF_X1 port map( A => n40741, Z => n40745);
   U28432 : BUF_X1 port map( A => n40747, Z => n40751);
   U28433 : BUF_X1 port map( A => n40753, Z => n40757);
   U28434 : BUF_X1 port map( A => n40759, Z => n40763);
   U28435 : BUF_X1 port map( A => n40765, Z => n40769);
   U28436 : BUF_X1 port map( A => n40771, Z => n40775);
   U28437 : BUF_X1 port map( A => n40777, Z => n40781);
   U28438 : BUF_X1 port map( A => n40783, Z => n40787);
   U28439 : BUF_X1 port map( A => n40789, Z => n40793);
   U28440 : BUF_X1 port map( A => n40795, Z => n40799);
   U28441 : BUF_X1 port map( A => n40801, Z => n40805);
   U28442 : BUF_X1 port map( A => n40807, Z => n40811);
   U28443 : BUF_X1 port map( A => n40813, Z => n40817);
   U28444 : BUF_X1 port map( A => n40819, Z => n40823);
   U28445 : BUF_X1 port map( A => n40825, Z => n40829);
   U28446 : BUF_X1 port map( A => n40831, Z => n40835);
   U28447 : BUF_X1 port map( A => n40837, Z => n40841);
   U28448 : BUF_X1 port map( A => n40843, Z => n40847);
   U28449 : BUF_X1 port map( A => n40849, Z => n40853);
   U28450 : BUF_X1 port map( A => n40855, Z => n40859);
   U28451 : BUF_X1 port map( A => n40861, Z => n40865);
   U28452 : BUF_X1 port map( A => n40867, Z => n40871);
   U28453 : BUF_X1 port map( A => n40873, Z => n40877);
   U28454 : BUF_X1 port map( A => n40879, Z => n40883);
   U28455 : BUF_X1 port map( A => n40885, Z => n40889);
   U28456 : BUF_X1 port map( A => n40891, Z => n40895);
   U28457 : BUF_X1 port map( A => n40897, Z => n40901);
   U28458 : BUF_X1 port map( A => n40903, Z => n40907);
   U28459 : BUF_X1 port map( A => n40909, Z => n40913);
   U28460 : BUF_X1 port map( A => n40915, Z => n40919);
   U28461 : BUF_X1 port map( A => n40921, Z => n40925);
   U28462 : BUF_X1 port map( A => n40927, Z => n40931);
   U28463 : BUF_X1 port map( A => n40933, Z => n40937);
   U28464 : BUF_X1 port map( A => n40939, Z => n40943);
   U28465 : BUF_X1 port map( A => n40945, Z => n40949);
   U28466 : BUF_X1 port map( A => n40951, Z => n40955);
   U28467 : BUF_X1 port map( A => n40957, Z => n40961);
   U28468 : BUF_X1 port map( A => n40963, Z => n40967);
   U28469 : BUF_X1 port map( A => n40969, Z => n40973);
   U28470 : BUF_X1 port map( A => n40975, Z => n40979);
   U28471 : NAND2_X1 port map( A1 => n32244, A2 => n33208, ZN => n34697);
   U28472 : NAND2_X1 port map( A1 => n32244, A2 => n33207, ZN => n35971);
   U28473 : OAI221_X1 port map( B1 => n33258, B2 => n33274, C1 => n33259, C2 =>
                           n33275, A => n41364, ZN => n33273);
   U28474 : OAI221_X1 port map( B1 => n33258, B2 => n33264, C1 => n33259, C2 =>
                           n33265, A => n41364, ZN => n33263);
   U28475 : OAI221_X1 port map( B1 => n33258, B2 => n33269, C1 => n33259, C2 =>
                           n33270, A => n41364, ZN => n33268);
   U28476 : OAI221_X1 port map( B1 => n33258, B2 => n32157, C1 => n33259, C2 =>
                           n33280, A => n41365, ZN => n33278);
   U28477 : OAI221_X1 port map( B1 => n33258, B2 => n33255, C1 => n33259, C2 =>
                           n33260, A => n41364, ZN => n33254);
   U28478 : OAI221_X1 port map( B1 => n33258, B2 => n32158, C1 => n33259, C2 =>
                           n33285, A => n41364, ZN => n33283);
   U28479 : OAI221_X1 port map( B1 => n33258, B2 => n32159, C1 => n33259, C2 =>
                           n33290, A => n41365, ZN => n33288);
   U28480 : OAI221_X1 port map( B1 => n33258, B2 => n32160, C1 => n33259, C2 =>
                           n33296, A => n41365, ZN => n33293);
   U28481 : NOR3_X1 port map( A1 => n32254, A2 => N689, A3 => n32251, ZN => 
                           n37231);
   U28482 : NOR3_X1 port map( A1 => n34694, A2 => N6271, A3 => n32166, ZN => 
                           n34676);
   U28483 : NOR3_X1 port map( A1 => n35968, A2 => N6396, A3 => n32171, ZN => 
                           n35950);
   U28484 : NOR3_X1 port map( A1 => n33398, A2 => N689, A3 => n32251, ZN => 
                           n37234);
   U28485 : NOR3_X1 port map( A1 => N688, A2 => N689, A3 => n32254, ZN => 
                           n37235);
   U28486 : NOR3_X1 port map( A1 => n33398, A2 => N688, A3 => n32248, ZN => 
                           n37230);
   U28487 : NOR3_X1 port map( A1 => N688, A2 => N689, A3 => n33398, ZN => 
                           n37233);
   U28488 : NOR3_X1 port map( A1 => n32254, A2 => N688, A3 => n32248, ZN => 
                           n37227);
   U28489 : NOR3_X1 port map( A1 => n32168, A2 => N6270, A3 => n32165, ZN => 
                           n34675);
   U28490 : NOR3_X1 port map( A1 => n32173, A2 => N6395, A3 => n32170, ZN => 
                           n35949);
   U28491 : NOR3_X1 port map( A1 => n33398, A2 => n32251, A3 => n32248, ZN => 
                           n37229);
   U28492 : NOR3_X1 port map( A1 => n32166, A2 => N6271, A3 => n32168, ZN => 
                           n34679);
   U28493 : NOR3_X1 port map( A1 => n32171, A2 => N6396, A3 => n32173, ZN => 
                           n35953);
   U28494 : NOR3_X1 port map( A1 => N6270, A2 => N6271, A3 => n34694, ZN => 
                           n34680);
   U28495 : NOR3_X1 port map( A1 => N6395, A2 => N6396, A3 => n35968, ZN => 
                           n35954);
   U28496 : NOR3_X1 port map( A1 => N6270, A2 => N6271, A3 => n32168, ZN => 
                           n34678);
   U28497 : NOR3_X1 port map( A1 => n34694, A2 => N6270, A3 => n32165, ZN => 
                           n34671);
   U28498 : NOR3_X1 port map( A1 => N6395, A2 => N6396, A3 => n32173, ZN => 
                           n35952);
   U28499 : NOR3_X1 port map( A1 => n35968, A2 => N6395, A3 => n32170, ZN => 
                           n35945);
   U28500 : NOR3_X1 port map( A1 => n32166, A2 => n34694, A3 => n32165, ZN => 
                           n34673);
   U28501 : NOR3_X1 port map( A1 => n32171, A2 => n35968, A3 => n32170, ZN => 
                           n35947);
   U28502 : NOR2_X1 port map( A1 => n37240, A2 => N690, ZN => n37239);
   U28503 : NOR2_X1 port map( A1 => n32164, A2 => N6273, ZN => n34690);
   U28504 : NOR2_X1 port map( A1 => n32169, A2 => N6398, ZN => n35964);
   U28505 : NOR3_X1 port map( A1 => N929, A2 => N930, A3 => n33402, ZN => 
                           n33289);
   U28506 : NOR3_X1 port map( A1 => n33402, A2 => N930, A3 => n32161, ZN => 
                           n33279);
   U28507 : NOR3_X1 port map( A1 => n32161, A2 => N930, A3 => n32163, ZN => 
                           n33284);
   U28508 : NOR3_X1 port map( A1 => N929, A2 => N930, A3 => n32163, ZN => 
                           n33295);
   U28509 : NOR2_X1 port map( A1 => n32246, A2 => n37240, ZN => n37236);
   U28510 : NAND2_X1 port map( A1 => n32244, A2 => n33209, ZN => n33422);
   U28511 : NAND3_X1 port map( A1 => N929, A2 => n32163, A3 => N930, ZN => 
                           n33255);
   U28512 : AOI221_X1 port map( B1 => n39638, B2 => n32822, C1 => n39632, C2 =>
                           n32774, A => n33558, ZN => n33555);
   U28513 : OAI222_X1 port map( A1 => n30988, A2 => n39626, B1 => n31052, B2 =>
                           n39620, C1 => n30924, C2 => n39614, ZN => n33558);
   U28514 : AOI221_X1 port map( B1 => n39386, B2 => n32822, C1 => n39380, C2 =>
                           n32774, A => n34832, ZN => n34829);
   U28515 : OAI222_X1 port map( A1 => n30988, A2 => n39374, B1 => n31052, B2 =>
                           n39368, C1 => n30924, C2 => n39362, ZN => n34832);
   U28516 : AOI221_X1 port map( B1 => n39638, B2 => n32821, C1 => n39632, C2 =>
                           n32773, A => n33577, ZN => n33574);
   U28517 : OAI222_X1 port map( A1 => n30987, A2 => n39626, B1 => n31051, B2 =>
                           n39620, C1 => n30923, C2 => n39614, ZN => n33577);
   U28518 : AOI221_X1 port map( B1 => n39386, B2 => n32821, C1 => n39380, C2 =>
                           n32773, A => n34851, ZN => n34848);
   U28519 : OAI222_X1 port map( A1 => n30987, A2 => n39374, B1 => n31051, B2 =>
                           n39368, C1 => n30923, C2 => n39362, ZN => n34851);
   U28520 : AOI221_X1 port map( B1 => n39638, B2 => n32820, C1 => n39632, C2 =>
                           n32772, A => n33596, ZN => n33593);
   U28521 : OAI222_X1 port map( A1 => n30986, A2 => n39626, B1 => n31050, B2 =>
                           n39620, C1 => n30922, C2 => n39614, ZN => n33596);
   U28522 : AOI221_X1 port map( B1 => n39386, B2 => n32820, C1 => n39380, C2 =>
                           n32772, A => n34870, ZN => n34867);
   U28523 : OAI222_X1 port map( A1 => n30986, A2 => n39374, B1 => n31050, B2 =>
                           n39368, C1 => n30922, C2 => n39362, ZN => n34870);
   U28524 : AOI221_X1 port map( B1 => n39638, B2 => n32819, C1 => n39632, C2 =>
                           n32771, A => n33615, ZN => n33612);
   U28525 : OAI222_X1 port map( A1 => n30985, A2 => n39626, B1 => n31049, B2 =>
                           n39620, C1 => n30921, C2 => n39614, ZN => n33615);
   U28526 : AOI221_X1 port map( B1 => n39386, B2 => n32819, C1 => n39380, C2 =>
                           n32771, A => n34889, ZN => n34886);
   U28527 : OAI222_X1 port map( A1 => n30985, A2 => n39374, B1 => n31049, B2 =>
                           n39368, C1 => n30921, C2 => n39362, ZN => n34889);
   U28528 : AOI221_X1 port map( B1 => n39638, B2 => n32818, C1 => n39632, C2 =>
                           n32770, A => n33634, ZN => n33631);
   U28529 : OAI222_X1 port map( A1 => n30984, A2 => n39626, B1 => n31048, B2 =>
                           n39620, C1 => n30920, C2 => n39614, ZN => n33634);
   U28530 : AOI221_X1 port map( B1 => n39386, B2 => n32818, C1 => n39380, C2 =>
                           n32770, A => n34908, ZN => n34905);
   U28531 : OAI222_X1 port map( A1 => n30984, A2 => n39374, B1 => n31048, B2 =>
                           n39368, C1 => n30920, C2 => n39362, ZN => n34908);
   U28532 : AOI221_X1 port map( B1 => n39638, B2 => n32817, C1 => n39632, C2 =>
                           n32769, A => n33653, ZN => n33650);
   U28533 : OAI222_X1 port map( A1 => n30983, A2 => n39626, B1 => n31047, B2 =>
                           n39620, C1 => n30919, C2 => n39614, ZN => n33653);
   U28534 : AOI221_X1 port map( B1 => n39386, B2 => n32817, C1 => n39380, C2 =>
                           n32769, A => n34927, ZN => n34924);
   U28535 : OAI222_X1 port map( A1 => n30983, A2 => n39374, B1 => n31047, B2 =>
                           n39368, C1 => n30919, C2 => n39362, ZN => n34927);
   U28536 : AOI221_X1 port map( B1 => n39638, B2 => n32816, C1 => n39632, C2 =>
                           n32768, A => n33672, ZN => n33669);
   U28537 : OAI222_X1 port map( A1 => n30982, A2 => n39626, B1 => n31046, B2 =>
                           n39620, C1 => n30918, C2 => n39614, ZN => n33672);
   U28538 : AOI221_X1 port map( B1 => n39386, B2 => n32816, C1 => n39380, C2 =>
                           n32768, A => n34946, ZN => n34943);
   U28539 : OAI222_X1 port map( A1 => n30982, A2 => n39374, B1 => n31046, B2 =>
                           n39368, C1 => n30918, C2 => n39362, ZN => n34946);
   U28540 : AOI221_X1 port map( B1 => n39638, B2 => n32815, C1 => n39632, C2 =>
                           n32767, A => n33691, ZN => n33688);
   U28541 : OAI222_X1 port map( A1 => n30981, A2 => n39626, B1 => n31045, B2 =>
                           n39620, C1 => n30917, C2 => n39614, ZN => n33691);
   U28542 : AOI221_X1 port map( B1 => n39386, B2 => n32815, C1 => n39380, C2 =>
                           n32767, A => n34965, ZN => n34962);
   U28543 : OAI222_X1 port map( A1 => n30981, A2 => n39374, B1 => n31045, B2 =>
                           n39368, C1 => n30917, C2 => n39362, ZN => n34965);
   U28544 : AOI221_X1 port map( B1 => n39638, B2 => n32814, C1 => n39632, C2 =>
                           n32766, A => n33710, ZN => n33707);
   U28545 : OAI222_X1 port map( A1 => n30980, A2 => n39626, B1 => n31044, B2 =>
                           n39620, C1 => n30916, C2 => n39614, ZN => n33710);
   U28546 : AOI221_X1 port map( B1 => n39386, B2 => n32814, C1 => n39380, C2 =>
                           n32766, A => n34984, ZN => n34981);
   U28547 : OAI222_X1 port map( A1 => n30980, A2 => n39374, B1 => n31044, B2 =>
                           n39368, C1 => n30916, C2 => n39362, ZN => n34984);
   U28548 : AOI221_X1 port map( B1 => n39638, B2 => n32813, C1 => n39632, C2 =>
                           n32765, A => n33729, ZN => n33726);
   U28549 : OAI222_X1 port map( A1 => n30979, A2 => n39626, B1 => n31043, B2 =>
                           n39620, C1 => n30915, C2 => n39614, ZN => n33729);
   U28550 : AOI221_X1 port map( B1 => n39386, B2 => n32813, C1 => n39380, C2 =>
                           n32765, A => n35003, ZN => n35000);
   U28551 : OAI222_X1 port map( A1 => n30979, A2 => n39374, B1 => n31043, B2 =>
                           n39368, C1 => n30915, C2 => n39362, ZN => n35003);
   U28552 : AOI221_X1 port map( B1 => n39638, B2 => n32812, C1 => n39632, C2 =>
                           n32764, A => n33748, ZN => n33745);
   U28553 : OAI222_X1 port map( A1 => n30978, A2 => n39626, B1 => n31042, B2 =>
                           n39620, C1 => n30914, C2 => n39614, ZN => n33748);
   U28554 : AOI221_X1 port map( B1 => n39386, B2 => n32812, C1 => n39380, C2 =>
                           n32764, A => n35022, ZN => n35019);
   U28555 : OAI222_X1 port map( A1 => n30978, A2 => n39374, B1 => n31042, B2 =>
                           n39368, C1 => n30914, C2 => n39362, ZN => n35022);
   U28556 : AOI221_X1 port map( B1 => n39638, B2 => n32811, C1 => n39632, C2 =>
                           n32763, A => n33767, ZN => n33764);
   U28557 : OAI222_X1 port map( A1 => n30977, A2 => n39626, B1 => n31041, B2 =>
                           n39620, C1 => n30913, C2 => n39614, ZN => n33767);
   U28558 : AOI221_X1 port map( B1 => n39386, B2 => n32811, C1 => n39380, C2 =>
                           n32763, A => n35041, ZN => n35038);
   U28559 : OAI222_X1 port map( A1 => n30977, A2 => n39374, B1 => n31041, B2 =>
                           n39368, C1 => n30913, C2 => n39362, ZN => n35041);
   U28560 : AOI221_X1 port map( B1 => n39637, B2 => n32810, C1 => n39631, C2 =>
                           n32762, A => n33786, ZN => n33783);
   U28561 : OAI222_X1 port map( A1 => n30976, A2 => n39625, B1 => n31040, B2 =>
                           n39619, C1 => n30912, C2 => n39613, ZN => n33786);
   U28562 : AOI221_X1 port map( B1 => n39385, B2 => n32810, C1 => n39379, C2 =>
                           n32762, A => n35060, ZN => n35057);
   U28563 : OAI222_X1 port map( A1 => n30976, A2 => n39373, B1 => n31040, B2 =>
                           n39367, C1 => n30912, C2 => n39361, ZN => n35060);
   U28564 : AOI221_X1 port map( B1 => n39637, B2 => n32809, C1 => n39631, C2 =>
                           n32761, A => n33805, ZN => n33802);
   U28565 : OAI222_X1 port map( A1 => n30975, A2 => n39625, B1 => n31039, B2 =>
                           n39619, C1 => n30911, C2 => n39613, ZN => n33805);
   U28566 : AOI221_X1 port map( B1 => n39385, B2 => n32809, C1 => n39379, C2 =>
                           n32761, A => n35079, ZN => n35076);
   U28567 : OAI222_X1 port map( A1 => n30975, A2 => n39373, B1 => n31039, B2 =>
                           n39367, C1 => n30911, C2 => n39361, ZN => n35079);
   U28568 : AOI221_X1 port map( B1 => n39637, B2 => n32808, C1 => n39631, C2 =>
                           n32760, A => n33824, ZN => n33821);
   U28569 : OAI222_X1 port map( A1 => n30974, A2 => n39625, B1 => n31038, B2 =>
                           n39619, C1 => n30910, C2 => n39613, ZN => n33824);
   U28570 : AOI221_X1 port map( B1 => n39385, B2 => n32808, C1 => n39379, C2 =>
                           n32760, A => n35098, ZN => n35095);
   U28571 : OAI222_X1 port map( A1 => n30974, A2 => n39373, B1 => n31038, B2 =>
                           n39367, C1 => n30910, C2 => n39361, ZN => n35098);
   U28572 : AOI221_X1 port map( B1 => n39637, B2 => n32807, C1 => n39631, C2 =>
                           n32759, A => n33843, ZN => n33840);
   U28573 : OAI222_X1 port map( A1 => n30973, A2 => n39625, B1 => n31037, B2 =>
                           n39619, C1 => n30909, C2 => n39613, ZN => n33843);
   U28574 : AOI221_X1 port map( B1 => n39385, B2 => n32807, C1 => n39379, C2 =>
                           n32759, A => n35117, ZN => n35114);
   U28575 : OAI222_X1 port map( A1 => n30973, A2 => n39373, B1 => n31037, B2 =>
                           n39367, C1 => n30909, C2 => n39361, ZN => n35117);
   U28576 : AOI221_X1 port map( B1 => n39637, B2 => n32806, C1 => n39631, C2 =>
                           n32758, A => n33862, ZN => n33859);
   U28577 : OAI222_X1 port map( A1 => n30972, A2 => n39625, B1 => n31036, B2 =>
                           n39619, C1 => n30908, C2 => n39613, ZN => n33862);
   U28578 : AOI221_X1 port map( B1 => n39385, B2 => n32806, C1 => n39379, C2 =>
                           n32758, A => n35136, ZN => n35133);
   U28579 : OAI222_X1 port map( A1 => n30972, A2 => n39373, B1 => n31036, B2 =>
                           n39367, C1 => n30908, C2 => n39361, ZN => n35136);
   U28580 : AOI221_X1 port map( B1 => n39637, B2 => n32805, C1 => n39631, C2 =>
                           n32757, A => n33881, ZN => n33878);
   U28581 : OAI222_X1 port map( A1 => n30971, A2 => n39625, B1 => n31035, B2 =>
                           n39619, C1 => n30907, C2 => n39613, ZN => n33881);
   U28582 : AOI221_X1 port map( B1 => n39385, B2 => n32805, C1 => n39379, C2 =>
                           n32757, A => n35155, ZN => n35152);
   U28583 : OAI222_X1 port map( A1 => n30971, A2 => n39373, B1 => n31035, B2 =>
                           n39367, C1 => n30907, C2 => n39361, ZN => n35155);
   U28584 : AOI221_X1 port map( B1 => n39637, B2 => n32804, C1 => n39631, C2 =>
                           n32756, A => n33900, ZN => n33897);
   U28585 : OAI222_X1 port map( A1 => n30970, A2 => n39625, B1 => n31034, B2 =>
                           n39619, C1 => n30906, C2 => n39613, ZN => n33900);
   U28586 : AOI221_X1 port map( B1 => n39385, B2 => n32804, C1 => n39379, C2 =>
                           n32756, A => n35174, ZN => n35171);
   U28587 : OAI222_X1 port map( A1 => n30970, A2 => n39373, B1 => n31034, B2 =>
                           n39367, C1 => n30906, C2 => n39361, ZN => n35174);
   U28588 : AOI221_X1 port map( B1 => n39637, B2 => n32803, C1 => n39631, C2 =>
                           n32755, A => n33919, ZN => n33916);
   U28589 : OAI222_X1 port map( A1 => n30969, A2 => n39625, B1 => n31033, B2 =>
                           n39619, C1 => n30905, C2 => n39613, ZN => n33919);
   U28590 : AOI221_X1 port map( B1 => n39385, B2 => n32803, C1 => n39379, C2 =>
                           n32755, A => n35193, ZN => n35190);
   U28591 : OAI222_X1 port map( A1 => n30969, A2 => n39373, B1 => n31033, B2 =>
                           n39367, C1 => n30905, C2 => n39361, ZN => n35193);
   U28592 : AOI221_X1 port map( B1 => n39637, B2 => n32802, C1 => n39631, C2 =>
                           n32754, A => n33938, ZN => n33935);
   U28593 : OAI222_X1 port map( A1 => n30968, A2 => n39625, B1 => n31032, B2 =>
                           n39619, C1 => n30904, C2 => n39613, ZN => n33938);
   U28594 : AOI221_X1 port map( B1 => n39385, B2 => n32802, C1 => n39379, C2 =>
                           n32754, A => n35212, ZN => n35209);
   U28595 : OAI222_X1 port map( A1 => n30968, A2 => n39373, B1 => n31032, B2 =>
                           n39367, C1 => n30904, C2 => n39361, ZN => n35212);
   U28596 : AOI221_X1 port map( B1 => n39637, B2 => n32801, C1 => n39631, C2 =>
                           n32753, A => n33957, ZN => n33954);
   U28597 : OAI222_X1 port map( A1 => n30967, A2 => n39625, B1 => n31031, B2 =>
                           n39619, C1 => n30903, C2 => n39613, ZN => n33957);
   U28598 : AOI221_X1 port map( B1 => n39385, B2 => n32801, C1 => n39379, C2 =>
                           n32753, A => n35231, ZN => n35228);
   U28599 : OAI222_X1 port map( A1 => n30967, A2 => n39373, B1 => n31031, B2 =>
                           n39367, C1 => n30903, C2 => n39361, ZN => n35231);
   U28600 : AOI221_X1 port map( B1 => n39637, B2 => n32800, C1 => n39631, C2 =>
                           n32752, A => n33976, ZN => n33973);
   U28601 : OAI222_X1 port map( A1 => n30966, A2 => n39625, B1 => n31030, B2 =>
                           n39619, C1 => n30902, C2 => n39613, ZN => n33976);
   U28602 : AOI221_X1 port map( B1 => n39385, B2 => n32800, C1 => n39379, C2 =>
                           n32752, A => n35250, ZN => n35247);
   U28603 : OAI222_X1 port map( A1 => n30966, A2 => n39373, B1 => n31030, B2 =>
                           n39367, C1 => n30902, C2 => n39361, ZN => n35250);
   U28604 : AOI221_X1 port map( B1 => n39637, B2 => n32799, C1 => n39631, C2 =>
                           n32751, A => n33995, ZN => n33992);
   U28605 : OAI222_X1 port map( A1 => n30965, A2 => n39625, B1 => n31029, B2 =>
                           n39619, C1 => n30901, C2 => n39613, ZN => n33995);
   U28606 : AOI221_X1 port map( B1 => n39385, B2 => n32799, C1 => n39379, C2 =>
                           n32751, A => n35269, ZN => n35266);
   U28607 : OAI222_X1 port map( A1 => n30965, A2 => n39373, B1 => n31029, B2 =>
                           n39367, C1 => n30901, C2 => n39361, ZN => n35269);
   U28608 : AOI221_X1 port map( B1 => n39636, B2 => n32798, C1 => n39630, C2 =>
                           n32750, A => n34014, ZN => n34011);
   U28609 : OAI222_X1 port map( A1 => n30964, A2 => n39624, B1 => n31028, B2 =>
                           n39618, C1 => n30900, C2 => n39612, ZN => n34014);
   U28610 : AOI221_X1 port map( B1 => n39384, B2 => n32798, C1 => n39378, C2 =>
                           n32750, A => n35288, ZN => n35285);
   U28611 : OAI222_X1 port map( A1 => n30964, A2 => n39372, B1 => n31028, B2 =>
                           n39366, C1 => n30900, C2 => n39360, ZN => n35288);
   U28612 : AOI221_X1 port map( B1 => n39636, B2 => n32797, C1 => n39630, C2 =>
                           n32749, A => n34033, ZN => n34030);
   U28613 : OAI222_X1 port map( A1 => n30963, A2 => n39624, B1 => n31027, B2 =>
                           n39618, C1 => n30899, C2 => n39612, ZN => n34033);
   U28614 : AOI221_X1 port map( B1 => n39384, B2 => n32797, C1 => n39378, C2 =>
                           n32749, A => n35307, ZN => n35304);
   U28615 : OAI222_X1 port map( A1 => n30963, A2 => n39372, B1 => n31027, B2 =>
                           n39366, C1 => n30899, C2 => n39360, ZN => n35307);
   U28616 : AOI221_X1 port map( B1 => n39636, B2 => n32796, C1 => n39630, C2 =>
                           n32748, A => n34052, ZN => n34049);
   U28617 : OAI222_X1 port map( A1 => n30962, A2 => n39624, B1 => n31026, B2 =>
                           n39618, C1 => n30898, C2 => n39612, ZN => n34052);
   U28618 : AOI221_X1 port map( B1 => n39384, B2 => n32796, C1 => n39378, C2 =>
                           n32748, A => n35326, ZN => n35323);
   U28619 : OAI222_X1 port map( A1 => n30962, A2 => n39372, B1 => n31026, B2 =>
                           n39366, C1 => n30898, C2 => n39360, ZN => n35326);
   U28620 : AOI221_X1 port map( B1 => n39636, B2 => n32795, C1 => n39630, C2 =>
                           n32747, A => n34071, ZN => n34068);
   U28621 : OAI222_X1 port map( A1 => n30961, A2 => n39624, B1 => n31025, B2 =>
                           n39618, C1 => n30897, C2 => n39612, ZN => n34071);
   U28622 : AOI221_X1 port map( B1 => n39384, B2 => n32795, C1 => n39378, C2 =>
                           n32747, A => n35345, ZN => n35342);
   U28623 : OAI222_X1 port map( A1 => n30961, A2 => n39372, B1 => n31025, B2 =>
                           n39366, C1 => n30897, C2 => n39360, ZN => n35345);
   U28624 : AOI221_X1 port map( B1 => n39636, B2 => n32794, C1 => n39630, C2 =>
                           n32746, A => n34090, ZN => n34087);
   U28625 : OAI222_X1 port map( A1 => n30960, A2 => n39624, B1 => n31024, B2 =>
                           n39618, C1 => n30896, C2 => n39612, ZN => n34090);
   U28626 : AOI221_X1 port map( B1 => n39384, B2 => n32794, C1 => n39378, C2 =>
                           n32746, A => n35364, ZN => n35361);
   U28627 : OAI222_X1 port map( A1 => n30960, A2 => n39372, B1 => n31024, B2 =>
                           n39366, C1 => n30896, C2 => n39360, ZN => n35364);
   U28628 : AOI221_X1 port map( B1 => n39636, B2 => n32793, C1 => n39630, C2 =>
                           n32745, A => n34109, ZN => n34106);
   U28629 : OAI222_X1 port map( A1 => n30959, A2 => n39624, B1 => n31023, B2 =>
                           n39618, C1 => n30895, C2 => n39612, ZN => n34109);
   U28630 : AOI221_X1 port map( B1 => n39384, B2 => n32793, C1 => n39378, C2 =>
                           n32745, A => n35383, ZN => n35380);
   U28631 : OAI222_X1 port map( A1 => n30959, A2 => n39372, B1 => n31023, B2 =>
                           n39366, C1 => n30895, C2 => n39360, ZN => n35383);
   U28632 : AOI221_X1 port map( B1 => n39636, B2 => n32792, C1 => n39630, C2 =>
                           n32744, A => n34128, ZN => n34125);
   U28633 : OAI222_X1 port map( A1 => n30958, A2 => n39624, B1 => n31022, B2 =>
                           n39618, C1 => n30894, C2 => n39612, ZN => n34128);
   U28634 : AOI221_X1 port map( B1 => n39384, B2 => n32792, C1 => n39378, C2 =>
                           n32744, A => n35402, ZN => n35399);
   U28635 : OAI222_X1 port map( A1 => n30958, A2 => n39372, B1 => n31022, B2 =>
                           n39366, C1 => n30894, C2 => n39360, ZN => n35402);
   U28636 : AOI221_X1 port map( B1 => n39636, B2 => n32791, C1 => n39630, C2 =>
                           n32743, A => n34147, ZN => n34144);
   U28637 : OAI222_X1 port map( A1 => n30957, A2 => n39624, B1 => n31021, B2 =>
                           n39618, C1 => n30893, C2 => n39612, ZN => n34147);
   U28638 : AOI221_X1 port map( B1 => n39384, B2 => n32791, C1 => n39378, C2 =>
                           n32743, A => n35421, ZN => n35418);
   U28639 : OAI222_X1 port map( A1 => n30957, A2 => n39372, B1 => n31021, B2 =>
                           n39366, C1 => n30893, C2 => n39360, ZN => n35421);
   U28640 : AOI221_X1 port map( B1 => n39636, B2 => n32790, C1 => n39630, C2 =>
                           n32742, A => n34166, ZN => n34163);
   U28641 : OAI222_X1 port map( A1 => n30956, A2 => n39624, B1 => n31020, B2 =>
                           n39618, C1 => n30892, C2 => n39612, ZN => n34166);
   U28642 : AOI221_X1 port map( B1 => n39384, B2 => n32790, C1 => n39378, C2 =>
                           n32742, A => n35440, ZN => n35437);
   U28643 : OAI222_X1 port map( A1 => n30956, A2 => n39372, B1 => n31020, B2 =>
                           n39366, C1 => n30892, C2 => n39360, ZN => n35440);
   U28644 : AOI221_X1 port map( B1 => n39636, B2 => n32789, C1 => n39630, C2 =>
                           n32741, A => n34185, ZN => n34182);
   U28645 : OAI222_X1 port map( A1 => n30955, A2 => n39624, B1 => n31019, B2 =>
                           n39618, C1 => n30891, C2 => n39612, ZN => n34185);
   U28646 : AOI221_X1 port map( B1 => n39384, B2 => n32789, C1 => n39378, C2 =>
                           n32741, A => n35459, ZN => n35456);
   U28647 : OAI222_X1 port map( A1 => n30955, A2 => n39372, B1 => n31019, B2 =>
                           n39366, C1 => n30891, C2 => n39360, ZN => n35459);
   U28648 : AOI221_X1 port map( B1 => n39636, B2 => n32788, C1 => n39630, C2 =>
                           n32740, A => n34204, ZN => n34201);
   U28649 : OAI222_X1 port map( A1 => n30954, A2 => n39624, B1 => n31018, B2 =>
                           n39618, C1 => n30890, C2 => n39612, ZN => n34204);
   U28650 : AOI221_X1 port map( B1 => n39384, B2 => n32788, C1 => n39378, C2 =>
                           n32740, A => n35478, ZN => n35475);
   U28651 : OAI222_X1 port map( A1 => n30954, A2 => n39372, B1 => n31018, B2 =>
                           n39366, C1 => n30890, C2 => n39360, ZN => n35478);
   U28652 : AOI221_X1 port map( B1 => n39636, B2 => n32787, C1 => n39630, C2 =>
                           n32739, A => n34223, ZN => n34220);
   U28653 : OAI222_X1 port map( A1 => n30953, A2 => n39624, B1 => n31017, B2 =>
                           n39618, C1 => n30889, C2 => n39612, ZN => n34223);
   U28654 : AOI221_X1 port map( B1 => n39384, B2 => n32787, C1 => n39378, C2 =>
                           n32739, A => n35497, ZN => n35494);
   U28655 : OAI222_X1 port map( A1 => n30953, A2 => n39372, B1 => n31017, B2 =>
                           n39366, C1 => n30889, C2 => n39360, ZN => n35497);
   U28656 : AOI221_X1 port map( B1 => n39635, B2 => n32786, C1 => n39629, C2 =>
                           n32738, A => n34242, ZN => n34239);
   U28657 : OAI222_X1 port map( A1 => n30952, A2 => n39623, B1 => n31016, B2 =>
                           n39617, C1 => n30888, C2 => n39611, ZN => n34242);
   U28658 : AOI221_X1 port map( B1 => n39383, B2 => n32786, C1 => n39377, C2 =>
                           n32738, A => n35516, ZN => n35513);
   U28659 : OAI222_X1 port map( A1 => n30952, A2 => n39371, B1 => n31016, B2 =>
                           n39365, C1 => n30888, C2 => n39359, ZN => n35516);
   U28660 : AOI221_X1 port map( B1 => n39635, B2 => n32785, C1 => n39629, C2 =>
                           n32737, A => n34261, ZN => n34258);
   U28661 : OAI222_X1 port map( A1 => n30951, A2 => n39623, B1 => n31015, B2 =>
                           n39617, C1 => n30887, C2 => n39611, ZN => n34261);
   U28662 : AOI221_X1 port map( B1 => n39383, B2 => n32785, C1 => n39377, C2 =>
                           n32737, A => n35535, ZN => n35532);
   U28663 : OAI222_X1 port map( A1 => n30951, A2 => n39371, B1 => n31015, B2 =>
                           n39365, C1 => n30887, C2 => n39359, ZN => n35535);
   U28664 : AOI221_X1 port map( B1 => n39635, B2 => n32784, C1 => n39629, C2 =>
                           n32736, A => n34280, ZN => n34277);
   U28665 : OAI222_X1 port map( A1 => n30950, A2 => n39623, B1 => n31014, B2 =>
                           n39617, C1 => n30886, C2 => n39611, ZN => n34280);
   U28666 : AOI221_X1 port map( B1 => n39383, B2 => n32784, C1 => n39377, C2 =>
                           n32736, A => n35554, ZN => n35551);
   U28667 : OAI222_X1 port map( A1 => n30950, A2 => n39371, B1 => n31014, B2 =>
                           n39365, C1 => n30886, C2 => n39359, ZN => n35554);
   U28668 : AOI221_X1 port map( B1 => n39635, B2 => n32783, C1 => n39629, C2 =>
                           n32735, A => n34299, ZN => n34296);
   U28669 : OAI222_X1 port map( A1 => n30949, A2 => n39623, B1 => n31013, B2 =>
                           n39617, C1 => n30885, C2 => n39611, ZN => n34299);
   U28670 : AOI221_X1 port map( B1 => n39383, B2 => n32783, C1 => n39377, C2 =>
                           n32735, A => n35573, ZN => n35570);
   U28671 : OAI222_X1 port map( A1 => n30949, A2 => n39371, B1 => n31013, B2 =>
                           n39365, C1 => n30885, C2 => n39359, ZN => n35573);
   U28672 : AOI221_X1 port map( B1 => n39635, B2 => n32782, C1 => n39629, C2 =>
                           n32734, A => n34318, ZN => n34315);
   U28673 : OAI222_X1 port map( A1 => n30948, A2 => n39623, B1 => n31012, B2 =>
                           n39617, C1 => n30884, C2 => n39611, ZN => n34318);
   U28674 : AOI221_X1 port map( B1 => n39383, B2 => n32782, C1 => n39377, C2 =>
                           n32734, A => n35592, ZN => n35589);
   U28675 : OAI222_X1 port map( A1 => n30948, A2 => n39371, B1 => n31012, B2 =>
                           n39365, C1 => n30884, C2 => n39359, ZN => n35592);
   U28676 : AOI221_X1 port map( B1 => n39635, B2 => n32781, C1 => n39629, C2 =>
                           n32733, A => n34337, ZN => n34334);
   U28677 : OAI222_X1 port map( A1 => n30947, A2 => n39623, B1 => n31011, B2 =>
                           n39617, C1 => n30883, C2 => n39611, ZN => n34337);
   U28678 : AOI221_X1 port map( B1 => n39383, B2 => n32781, C1 => n39377, C2 =>
                           n32733, A => n35611, ZN => n35608);
   U28679 : OAI222_X1 port map( A1 => n30947, A2 => n39371, B1 => n31011, B2 =>
                           n39365, C1 => n30883, C2 => n39359, ZN => n35611);
   U28680 : AOI221_X1 port map( B1 => n39635, B2 => n32780, C1 => n39629, C2 =>
                           n32732, A => n34356, ZN => n34353);
   U28681 : OAI222_X1 port map( A1 => n30946, A2 => n39623, B1 => n31010, B2 =>
                           n39617, C1 => n30882, C2 => n39611, ZN => n34356);
   U28682 : AOI221_X1 port map( B1 => n39383, B2 => n32780, C1 => n39377, C2 =>
                           n32732, A => n35630, ZN => n35627);
   U28683 : OAI222_X1 port map( A1 => n30946, A2 => n39371, B1 => n31010, B2 =>
                           n39365, C1 => n30882, C2 => n39359, ZN => n35630);
   U28684 : AOI221_X1 port map( B1 => n39635, B2 => n32779, C1 => n39629, C2 =>
                           n32731, A => n34375, ZN => n34372);
   U28685 : OAI222_X1 port map( A1 => n30945, A2 => n39623, B1 => n31009, B2 =>
                           n39617, C1 => n30881, C2 => n39611, ZN => n34375);
   U28686 : AOI221_X1 port map( B1 => n39383, B2 => n32779, C1 => n39377, C2 =>
                           n32731, A => n35649, ZN => n35646);
   U28687 : OAI222_X1 port map( A1 => n30945, A2 => n39371, B1 => n31009, B2 =>
                           n39365, C1 => n30881, C2 => n39359, ZN => n35649);
   U28688 : AOI221_X1 port map( B1 => n39635, B2 => n32778, C1 => n39629, C2 =>
                           n32730, A => n34394, ZN => n34391);
   U28689 : OAI222_X1 port map( A1 => n30944, A2 => n39623, B1 => n31008, B2 =>
                           n39617, C1 => n30880, C2 => n39611, ZN => n34394);
   U28690 : AOI221_X1 port map( B1 => n39383, B2 => n32778, C1 => n39377, C2 =>
                           n32730, A => n35668, ZN => n35665);
   U28691 : OAI222_X1 port map( A1 => n30944, A2 => n39371, B1 => n31008, B2 =>
                           n39365, C1 => n30880, C2 => n39359, ZN => n35668);
   U28692 : AOI221_X1 port map( B1 => n39635, B2 => n32777, C1 => n39629, C2 =>
                           n32729, A => n34413, ZN => n34410);
   U28693 : OAI222_X1 port map( A1 => n30943, A2 => n39623, B1 => n31007, B2 =>
                           n39617, C1 => n30879, C2 => n39611, ZN => n34413);
   U28694 : AOI221_X1 port map( B1 => n39383, B2 => n32777, C1 => n39377, C2 =>
                           n32729, A => n35687, ZN => n35684);
   U28695 : OAI222_X1 port map( A1 => n30943, A2 => n39371, B1 => n31007, B2 =>
                           n39365, C1 => n30879, C2 => n39359, ZN => n35687);
   U28696 : AOI221_X1 port map( B1 => n39635, B2 => n32776, C1 => n39629, C2 =>
                           n32728, A => n34432, ZN => n34429);
   U28697 : OAI222_X1 port map( A1 => n30942, A2 => n39623, B1 => n31006, B2 =>
                           n39617, C1 => n30878, C2 => n39611, ZN => n34432);
   U28698 : AOI221_X1 port map( B1 => n39383, B2 => n32776, C1 => n39377, C2 =>
                           n32728, A => n35706, ZN => n35703);
   U28699 : OAI222_X1 port map( A1 => n30942, A2 => n39371, B1 => n31006, B2 =>
                           n39365, C1 => n30878, C2 => n39359, ZN => n35706);
   U28700 : AOI221_X1 port map( B1 => n39635, B2 => n32775, C1 => n39629, C2 =>
                           n32727, A => n34451, ZN => n34448);
   U28701 : OAI222_X1 port map( A1 => n30941, A2 => n39623, B1 => n31005, B2 =>
                           n39617, C1 => n30877, C2 => n39611, ZN => n34451);
   U28702 : AOI221_X1 port map( B1 => n39383, B2 => n32775, C1 => n39377, C2 =>
                           n32727, A => n35725, ZN => n35722);
   U28703 : OAI222_X1 port map( A1 => n30941, A2 => n39371, B1 => n31005, B2 =>
                           n39365, C1 => n30877, C2 => n39359, ZN => n35725);
   U28704 : AOI221_X1 port map( B1 => n39634, B2 => n32846, C1 => n39628, C2 =>
                           n32834, A => n34470, ZN => n34467);
   U28705 : OAI222_X1 port map( A1 => n30940, A2 => n39622, B1 => n31004, B2 =>
                           n39616, C1 => n30876, C2 => n39610, ZN => n34470);
   U28706 : AOI221_X1 port map( B1 => n39382, B2 => n32846, C1 => n39376, C2 =>
                           n32834, A => n35744, ZN => n35741);
   U28707 : OAI222_X1 port map( A1 => n30940, A2 => n39370, B1 => n31004, B2 =>
                           n39364, C1 => n30876, C2 => n39358, ZN => n35744);
   U28708 : AOI221_X1 port map( B1 => n39634, B2 => n32845, C1 => n39628, C2 =>
                           n32833, A => n34489, ZN => n34486);
   U28709 : OAI222_X1 port map( A1 => n30939, A2 => n39622, B1 => n31003, B2 =>
                           n39616, C1 => n30875, C2 => n39610, ZN => n34489);
   U28710 : AOI221_X1 port map( B1 => n39382, B2 => n32845, C1 => n39376, C2 =>
                           n32833, A => n35763, ZN => n35760);
   U28711 : OAI222_X1 port map( A1 => n30939, A2 => n39370, B1 => n31003, B2 =>
                           n39364, C1 => n30875, C2 => n39358, ZN => n35763);
   U28712 : AOI221_X1 port map( B1 => n39634, B2 => n32844, C1 => n39628, C2 =>
                           n32832, A => n34508, ZN => n34505);
   U28713 : OAI222_X1 port map( A1 => n30938, A2 => n39622, B1 => n31002, B2 =>
                           n39616, C1 => n30874, C2 => n39610, ZN => n34508);
   U28714 : AOI221_X1 port map( B1 => n39382, B2 => n32844, C1 => n39376, C2 =>
                           n32832, A => n35782, ZN => n35779);
   U28715 : OAI222_X1 port map( A1 => n30938, A2 => n39370, B1 => n31002, B2 =>
                           n39364, C1 => n30874, C2 => n39358, ZN => n35782);
   U28716 : AOI221_X1 port map( B1 => n39634, B2 => n32843, C1 => n39628, C2 =>
                           n32831, A => n34527, ZN => n34524);
   U28717 : OAI222_X1 port map( A1 => n30937, A2 => n39622, B1 => n31001, B2 =>
                           n39616, C1 => n30873, C2 => n39610, ZN => n34527);
   U28718 : AOI221_X1 port map( B1 => n39382, B2 => n32843, C1 => n39376, C2 =>
                           n32831, A => n35801, ZN => n35798);
   U28719 : OAI222_X1 port map( A1 => n30937, A2 => n39370, B1 => n31001, B2 =>
                           n39364, C1 => n30873, C2 => n39358, ZN => n35801);
   U28720 : AOI221_X1 port map( B1 => n39634, B2 => n32842, C1 => n39628, C2 =>
                           n32830, A => n34546, ZN => n34543);
   U28721 : OAI222_X1 port map( A1 => n30936, A2 => n39622, B1 => n31000, B2 =>
                           n39616, C1 => n30872, C2 => n39610, ZN => n34546);
   U28722 : AOI221_X1 port map( B1 => n39382, B2 => n32842, C1 => n39376, C2 =>
                           n32830, A => n35820, ZN => n35817);
   U28723 : OAI222_X1 port map( A1 => n30936, A2 => n39370, B1 => n31000, B2 =>
                           n39364, C1 => n30872, C2 => n39358, ZN => n35820);
   U28724 : AOI221_X1 port map( B1 => n39634, B2 => n32841, C1 => n39628, C2 =>
                           n32829, A => n34565, ZN => n34562);
   U28725 : OAI222_X1 port map( A1 => n30935, A2 => n39622, B1 => n30999, B2 =>
                           n39616, C1 => n30871, C2 => n39610, ZN => n34565);
   U28726 : AOI221_X1 port map( B1 => n39382, B2 => n32841, C1 => n39376, C2 =>
                           n32829, A => n35839, ZN => n35836);
   U28727 : OAI222_X1 port map( A1 => n30935, A2 => n39370, B1 => n30999, B2 =>
                           n39364, C1 => n30871, C2 => n39358, ZN => n35839);
   U28728 : AOI221_X1 port map( B1 => n39634, B2 => n32840, C1 => n39628, C2 =>
                           n32828, A => n34584, ZN => n34581);
   U28729 : OAI222_X1 port map( A1 => n30934, A2 => n39622, B1 => n30998, B2 =>
                           n39616, C1 => n30870, C2 => n39610, ZN => n34584);
   U28730 : AOI221_X1 port map( B1 => n39382, B2 => n32840, C1 => n39376, C2 =>
                           n32828, A => n35858, ZN => n35855);
   U28731 : OAI222_X1 port map( A1 => n30934, A2 => n39370, B1 => n30998, B2 =>
                           n39364, C1 => n30870, C2 => n39358, ZN => n35858);
   U28732 : AOI221_X1 port map( B1 => n39634, B2 => n32839, C1 => n39628, C2 =>
                           n32827, A => n34603, ZN => n34600);
   U28733 : OAI222_X1 port map( A1 => n30933, A2 => n39622, B1 => n30997, B2 =>
                           n39616, C1 => n30869, C2 => n39610, ZN => n34603);
   U28734 : AOI221_X1 port map( B1 => n39382, B2 => n32839, C1 => n39376, C2 =>
                           n32827, A => n35877, ZN => n35874);
   U28735 : OAI222_X1 port map( A1 => n30933, A2 => n39370, B1 => n30997, B2 =>
                           n39364, C1 => n30869, C2 => n39358, ZN => n35877);
   U28736 : AOI221_X1 port map( B1 => n39634, B2 => n32838, C1 => n39628, C2 =>
                           n32826, A => n34622, ZN => n34619);
   U28737 : OAI222_X1 port map( A1 => n30932, A2 => n39622, B1 => n30996, B2 =>
                           n39616, C1 => n30868, C2 => n39610, ZN => n34622);
   U28738 : AOI221_X1 port map( B1 => n39382, B2 => n32838, C1 => n39376, C2 =>
                           n32826, A => n35896, ZN => n35893);
   U28739 : OAI222_X1 port map( A1 => n30932, A2 => n39370, B1 => n30996, B2 =>
                           n39364, C1 => n30868, C2 => n39358, ZN => n35896);
   U28740 : AOI221_X1 port map( B1 => n39634, B2 => n32837, C1 => n39628, C2 =>
                           n32825, A => n34641, ZN => n34638);
   U28741 : OAI222_X1 port map( A1 => n30931, A2 => n39622, B1 => n30995, B2 =>
                           n39616, C1 => n30867, C2 => n39610, ZN => n34641);
   U28742 : AOI221_X1 port map( B1 => n39382, B2 => n32837, C1 => n39376, C2 =>
                           n32825, A => n35915, ZN => n35912);
   U28743 : OAI222_X1 port map( A1 => n30931, A2 => n39370, B1 => n30995, B2 =>
                           n39364, C1 => n30867, C2 => n39358, ZN => n35915);
   U28744 : AOI221_X1 port map( B1 => n39634, B2 => n32836, C1 => n39628, C2 =>
                           n32824, A => n34660, ZN => n34657);
   U28745 : OAI222_X1 port map( A1 => n30930, A2 => n39622, B1 => n30994, B2 =>
                           n39616, C1 => n30866, C2 => n39610, ZN => n34660);
   U28746 : AOI221_X1 port map( B1 => n39382, B2 => n32836, C1 => n39376, C2 =>
                           n32824, A => n35934, ZN => n35931);
   U28747 : OAI222_X1 port map( A1 => n30930, A2 => n39370, B1 => n30994, B2 =>
                           n39364, C1 => n30866, C2 => n39358, ZN => n35934);
   U28748 : AOI221_X1 port map( B1 => n39634, B2 => n32835, C1 => n39628, C2 =>
                           n32823, A => n34691, ZN => n34687);
   U28749 : OAI222_X1 port map( A1 => n30929, A2 => n39622, B1 => n30993, B2 =>
                           n39616, C1 => n30865, C2 => n39610, ZN => n34691);
   U28750 : AOI221_X1 port map( B1 => n39382, B2 => n32835, C1 => n39376, C2 =>
                           n32823, A => n35965, ZN => n35961);
   U28751 : OAI222_X1 port map( A1 => n30929, A2 => n39370, B1 => n30993, B2 =>
                           n39364, C1 => n30865, C2 => n39358, ZN => n35965);
   U28752 : NOR2_X1 port map( A1 => N932, A2 => N931, ZN => n33294);
   U28753 : OAI222_X1 port map( A1 => n40952, A2 => n39895, B1 => n41336, B2 =>
                           n39888, C1 => n39886, C2 => n30613, ZN => n7591);
   U28754 : OAI222_X1 port map( A1 => n40964, A2 => n39895, B1 => n41348, B2 =>
                           n39888, C1 => n39886, C2 => n30611, ZN => n7589);
   U28755 : OAI222_X1 port map( A1 => n40970, A2 => n39895, B1 => n41354, B2 =>
                           n39888, C1 => n39886, C2 => n30610, ZN => n7588);
   U28756 : OAI222_X1 port map( A1 => n40976, A2 => n39895, B1 => n41360, B2 =>
                           n39888, C1 => n39886, C2 => n30609, ZN => n7587);
   U28757 : OAI222_X1 port map( A1 => n40954, A2 => n40390, B1 => n41338, B2 =>
                           n40383, C1 => n40381, C2 => n31691, ZN => n9191);
   U28758 : OAI222_X1 port map( A1 => n40966, A2 => n40390, B1 => n41350, B2 =>
                           n40383, C1 => n40381, C2 => n31689, ZN => n9189);
   U28759 : OAI222_X1 port map( A1 => n40972, A2 => n40390, B1 => n41356, B2 =>
                           n40383, C1 => n40381, C2 => n31688, ZN => n9188);
   U28760 : OAI222_X1 port map( A1 => n40978, A2 => n40390, B1 => n41362, B2 =>
                           n40383, C1 => n40381, C2 => n31687, ZN => n9187);
   U28761 : OAI222_X1 port map( A1 => n40954, A2 => n40370, B1 => n41338, B2 =>
                           n40363, C1 => n40361, C2 => n31627, ZN => n9127);
   U28762 : OAI222_X1 port map( A1 => n40966, A2 => n40370, B1 => n41350, B2 =>
                           n40363, C1 => n40361, C2 => n31625, ZN => n9125);
   U28763 : OAI222_X1 port map( A1 => n40972, A2 => n40370, B1 => n41356, B2 =>
                           n40363, C1 => n40361, C2 => n31624, ZN => n9124);
   U28764 : OAI222_X1 port map( A1 => n40978, A2 => n40370, B1 => n41362, B2 =>
                           n40363, C1 => n40361, C2 => n31623, ZN => n9123);
   U28765 : OAI222_X1 port map( A1 => n40954, A2 => n40350, B1 => n41338, B2 =>
                           n40343, C1 => n40341, C2 => n31563, ZN => n9063);
   U28766 : OAI222_X1 port map( A1 => n40966, A2 => n40350, B1 => n41350, B2 =>
                           n40343, C1 => n40341, C2 => n31561, ZN => n9061);
   U28767 : OAI222_X1 port map( A1 => n40972, A2 => n40350, B1 => n41356, B2 =>
                           n40343, C1 => n40341, C2 => n31560, ZN => n9060);
   U28768 : OAI222_X1 port map( A1 => n40978, A2 => n40350, B1 => n41362, B2 =>
                           n40343, C1 => n40341, C2 => n31559, ZN => n9059);
   U28769 : OAI222_X1 port map( A1 => n40954, A2 => n40290, B1 => n41338, B2 =>
                           n40283, C1 => n40281, C2 => n31499, ZN => n8871);
   U28770 : OAI222_X1 port map( A1 => n40966, A2 => n40290, B1 => n41350, B2 =>
                           n40283, C1 => n40281, C2 => n31497, ZN => n8869);
   U28771 : OAI222_X1 port map( A1 => n40972, A2 => n40290, B1 => n41356, B2 =>
                           n40283, C1 => n40281, C2 => n31496, ZN => n8868);
   U28772 : OAI222_X1 port map( A1 => n40978, A2 => n40290, B1 => n41362, B2 =>
                           n40283, C1 => n40281, C2 => n31495, ZN => n8867);
   U28773 : OAI222_X1 port map( A1 => n40953, A2 => n40270, B1 => n41337, B2 =>
                           n40263, C1 => n40261, C2 => n31435, ZN => n8807);
   U28774 : OAI222_X1 port map( A1 => n40965, A2 => n40270, B1 => n41349, B2 =>
                           n40263, C1 => n40261, C2 => n31433, ZN => n8805);
   U28775 : OAI222_X1 port map( A1 => n40971, A2 => n40270, B1 => n41355, B2 =>
                           n40263, C1 => n40261, C2 => n31432, ZN => n8804);
   U28776 : OAI222_X1 port map( A1 => n40977, A2 => n40270, B1 => n41361, B2 =>
                           n40263, C1 => n40261, C2 => n31431, ZN => n8803);
   U28777 : OAI222_X1 port map( A1 => n40953, A2 => n40250, B1 => n41337, B2 =>
                           n40243, C1 => n40241, C2 => n31371, ZN => n8743);
   U28778 : OAI222_X1 port map( A1 => n40965, A2 => n40250, B1 => n41349, B2 =>
                           n40243, C1 => n40241, C2 => n31369, ZN => n8741);
   U28779 : OAI222_X1 port map( A1 => n40971, A2 => n40250, B1 => n41355, B2 =>
                           n40243, C1 => n40241, C2 => n31368, ZN => n8740);
   U28780 : OAI222_X1 port map( A1 => n40977, A2 => n40250, B1 => n41361, B2 =>
                           n40243, C1 => n40241, C2 => n31367, ZN => n8739);
   U28781 : OAI222_X1 port map( A1 => n40953, A2 => n40190, B1 => n41337, B2 =>
                           n40183, C1 => n40181, C2 => n31307, ZN => n8551);
   U28782 : OAI222_X1 port map( A1 => n40965, A2 => n40190, B1 => n41349, B2 =>
                           n40183, C1 => n40181, C2 => n31305, ZN => n8549);
   U28783 : OAI222_X1 port map( A1 => n40971, A2 => n40190, B1 => n41355, B2 =>
                           n40183, C1 => n40181, C2 => n31304, ZN => n8548);
   U28784 : OAI222_X1 port map( A1 => n40977, A2 => n40190, B1 => n41361, B2 =>
                           n40183, C1 => n40181, C2 => n31303, ZN => n8547);
   U28785 : OAI222_X1 port map( A1 => n40953, A2 => n40170, B1 => n41337, B2 =>
                           n40163, C1 => n40161, C2 => n31243, ZN => n8487);
   U28786 : OAI222_X1 port map( A1 => n40965, A2 => n40170, B1 => n41349, B2 =>
                           n40163, C1 => n40161, C2 => n31241, ZN => n8485);
   U28787 : OAI222_X1 port map( A1 => n40971, A2 => n40170, B1 => n41355, B2 =>
                           n40163, C1 => n40161, C2 => n31240, ZN => n8484);
   U28788 : OAI222_X1 port map( A1 => n40977, A2 => n40170, B1 => n41361, B2 =>
                           n40163, C1 => n40161, C2 => n31239, ZN => n8483);
   U28789 : OAI222_X1 port map( A1 => n40953, A2 => n40150, B1 => n41337, B2 =>
                           n40143, C1 => n40141, C2 => n31179, ZN => n8423);
   U28790 : OAI222_X1 port map( A1 => n40965, A2 => n40150, B1 => n41349, B2 =>
                           n40143, C1 => n40141, C2 => n31177, ZN => n8421);
   U28791 : OAI222_X1 port map( A1 => n40971, A2 => n40150, B1 => n41355, B2 =>
                           n40143, C1 => n40141, C2 => n31176, ZN => n8420);
   U28792 : OAI222_X1 port map( A1 => n40977, A2 => n40150, B1 => n41361, B2 =>
                           n40143, C1 => n40141, C2 => n31175, ZN => n8419);
   U28793 : OAI222_X1 port map( A1 => n40953, A2 => n40091, B1 => n41337, B2 =>
                           n40084, C1 => n40082, C2 => n30997, ZN => n8231);
   U28794 : OAI222_X1 port map( A1 => n40965, A2 => n40091, B1 => n41349, B2 =>
                           n40084, C1 => n40082, C2 => n30995, ZN => n8229);
   U28795 : OAI222_X1 port map( A1 => n40971, A2 => n40091, B1 => n41355, B2 =>
                           n40084, C1 => n40082, C2 => n30994, ZN => n8228);
   U28796 : OAI222_X1 port map( A1 => n40977, A2 => n40091, B1 => n41361, B2 =>
                           n40084, C1 => n40082, C2 => n30993, ZN => n8227);
   U28797 : OAI222_X1 port map( A1 => n40953, A2 => n40071, B1 => n41337, B2 =>
                           n40064, C1 => n40062, C2 => n30933, ZN => n8167);
   U28798 : OAI222_X1 port map( A1 => n40965, A2 => n40071, B1 => n41349, B2 =>
                           n40064, C1 => n40062, C2 => n30931, ZN => n8165);
   U28799 : OAI222_X1 port map( A1 => n40971, A2 => n40071, B1 => n41355, B2 =>
                           n40064, C1 => n40062, C2 => n30930, ZN => n8164);
   U28800 : OAI222_X1 port map( A1 => n40977, A2 => n40071, B1 => n41361, B2 =>
                           n40064, C1 => n40062, C2 => n30929, ZN => n8163);
   U28801 : OAI222_X1 port map( A1 => n40953, A2 => n40051, B1 => n41337, B2 =>
                           n40044, C1 => n40042, C2 => n30869, ZN => n8103);
   U28802 : OAI222_X1 port map( A1 => n40965, A2 => n40051, B1 => n41349, B2 =>
                           n40044, C1 => n40042, C2 => n30867, ZN => n8101);
   U28803 : OAI222_X1 port map( A1 => n40971, A2 => n40051, B1 => n41355, B2 =>
                           n40044, C1 => n40042, C2 => n30866, ZN => n8100);
   U28804 : OAI222_X1 port map( A1 => n40977, A2 => n40051, B1 => n41361, B2 =>
                           n40044, C1 => n40042, C2 => n30865, ZN => n8099);
   U28805 : OAI222_X1 port map( A1 => n40952, A2 => n39993, B1 => n41336, B2 =>
                           n39986, C1 => n39984, C2 => n30805, ZN => n7911);
   U28806 : OAI222_X1 port map( A1 => n40964, A2 => n39993, B1 => n41348, B2 =>
                           n39986, C1 => n39984, C2 => n30803, ZN => n7909);
   U28807 : OAI222_X1 port map( A1 => n40970, A2 => n39993, B1 => n41354, B2 =>
                           n39986, C1 => n39984, C2 => n30802, ZN => n7908);
   U28808 : OAI222_X1 port map( A1 => n40976, A2 => n39993, B1 => n41360, B2 =>
                           n39986, C1 => n39984, C2 => n30801, ZN => n7907);
   U28809 : OAI222_X1 port map( A1 => n40952, A2 => n39973, B1 => n41336, B2 =>
                           n39966, C1 => n39964, C2 => n30741, ZN => n7847);
   U28810 : OAI222_X1 port map( A1 => n40964, A2 => n39973, B1 => n41348, B2 =>
                           n39966, C1 => n39964, C2 => n30739, ZN => n7845);
   U28811 : OAI222_X1 port map( A1 => n40970, A2 => n39973, B1 => n41354, B2 =>
                           n39966, C1 => n39964, C2 => n30738, ZN => n7844);
   U28812 : OAI222_X1 port map( A1 => n40976, A2 => n39973, B1 => n41360, B2 =>
                           n39966, C1 => n39964, C2 => n30737, ZN => n7843);
   U28813 : OAI222_X1 port map( A1 => n40590, A2 => n40955, B1 => n40583, B2 =>
                           n41339, C1 => n40581, C2 => n32054, ZN => n9831);
   U28814 : OAI222_X1 port map( A1 => n40590, A2 => n40967, B1 => n40583, B2 =>
                           n41351, C1 => n40581, C2 => n32053, ZN => n9829);
   U28815 : OAI222_X1 port map( A1 => n40590, A2 => n40973, B1 => n40583, B2 =>
                           n41357, C1 => n40581, C2 => n32052, ZN => n9828);
   U28816 : OAI222_X1 port map( A1 => n40590, A2 => n40979, B1 => n40583, B2 =>
                           n41363, C1 => n40581, C2 => n32051, ZN => n9827);
   U28817 : OAI222_X1 port map( A1 => n40955, A2 => n40570, B1 => n41339, B2 =>
                           n40563, C1 => n40561, C2 => n31995, ZN => n9767);
   U28818 : OAI222_X1 port map( A1 => n40967, A2 => n40570, B1 => n41351, B2 =>
                           n40563, C1 => n40561, C2 => n31993, ZN => n9765);
   U28819 : OAI222_X1 port map( A1 => n40973, A2 => n40570, B1 => n41357, B2 =>
                           n40563, C1 => n40561, C2 => n31992, ZN => n9764);
   U28820 : OAI222_X1 port map( A1 => n40979, A2 => n40570, B1 => n41363, B2 =>
                           n40563, C1 => n40561, C2 => n31991, ZN => n9763);
   U28821 : OAI222_X1 port map( A1 => n40955, A2 => n40550, B1 => n41339, B2 =>
                           n40543, C1 => n40541, C2 => n31935, ZN => n9703);
   U28822 : OAI222_X1 port map( A1 => n40967, A2 => n40550, B1 => n41351, B2 =>
                           n40543, C1 => n40541, C2 => n31933, ZN => n9701);
   U28823 : OAI222_X1 port map( A1 => n40973, A2 => n40550, B1 => n41357, B2 =>
                           n40543, C1 => n40541, C2 => n31932, ZN => n9700);
   U28824 : OAI222_X1 port map( A1 => n40979, A2 => n40550, B1 => n41363, B2 =>
                           n40543, C1 => n40541, C2 => n31931, ZN => n9699);
   U28825 : OAI222_X1 port map( A1 => n40954, A2 => n40490, B1 => n41338, B2 =>
                           n40483, C1 => n40481, C2 => n31875, ZN => n9511);
   U28826 : OAI222_X1 port map( A1 => n40966, A2 => n40490, B1 => n41350, B2 =>
                           n40483, C1 => n40481, C2 => n31873, ZN => n9509);
   U28827 : OAI222_X1 port map( A1 => n40972, A2 => n40490, B1 => n41356, B2 =>
                           n40483, C1 => n40481, C2 => n31872, ZN => n9508);
   U28828 : OAI222_X1 port map( A1 => n40978, A2 => n40490, B1 => n41362, B2 =>
                           n40483, C1 => n40481, C2 => n31871, ZN => n9507);
   U28829 : OAI222_X1 port map( A1 => n40954, A2 => n40470, B1 => n41338, B2 =>
                           n40463, C1 => n40461, C2 => n31815, ZN => n9447);
   U28830 : OAI222_X1 port map( A1 => n40966, A2 => n40470, B1 => n41350, B2 =>
                           n40463, C1 => n40461, C2 => n31813, ZN => n9445);
   U28831 : OAI222_X1 port map( A1 => n40972, A2 => n40470, B1 => n41356, B2 =>
                           n40463, C1 => n40461, C2 => n31812, ZN => n9444);
   U28832 : OAI222_X1 port map( A1 => n40978, A2 => n40470, B1 => n41362, B2 =>
                           n40463, C1 => n40461, C2 => n31811, ZN => n9443);
   U28833 : OAI222_X1 port map( A1 => n40954, A2 => n40450, B1 => n41338, B2 =>
                           n40443, C1 => n40441, C2 => n31755, ZN => n9383);
   U28834 : OAI222_X1 port map( A1 => n40966, A2 => n40450, B1 => n41350, B2 =>
                           n40443, C1 => n40441, C2 => n31753, ZN => n9381);
   U28835 : OAI222_X1 port map( A1 => n40972, A2 => n40450, B1 => n41356, B2 =>
                           n40443, C1 => n40441, C2 => n31752, ZN => n9380);
   U28836 : OAI222_X1 port map( A1 => n40978, A2 => n40450, B1 => n41362, B2 =>
                           n40443, C1 => n40441, C2 => n31751, ZN => n9379);
   U28837 : OAI222_X1 port map( A1 => n40952, A2 => n39953, B1 => n41336, B2 =>
                           n39946, C1 => n39944, C2 => n30677, ZN => n7783);
   U28838 : OAI222_X1 port map( A1 => n40964, A2 => n39953, B1 => n41348, B2 =>
                           n39946, C1 => n39944, C2 => n30675, ZN => n7781);
   U28839 : OAI222_X1 port map( A1 => n40970, A2 => n39953, B1 => n41354, B2 =>
                           n39946, C1 => n39944, C2 => n30674, ZN => n7780);
   U28840 : OAI222_X1 port map( A1 => n40976, A2 => n39953, B1 => n41360, B2 =>
                           n39946, C1 => n39944, C2 => n30673, ZN => n7779);
   U28841 : OAI222_X1 port map( A1 => n40952, A2 => n39875, B1 => n41336, B2 =>
                           n39868, C1 => n39866, C2 => n30549, ZN => n7527);
   U28842 : OAI222_X1 port map( A1 => n40964, A2 => n39875, B1 => n41348, B2 =>
                           n39868, C1 => n39866, C2 => n30547, ZN => n7525);
   U28843 : OAI222_X1 port map( A1 => n40970, A2 => n39875, B1 => n41354, B2 =>
                           n39868, C1 => n39866, C2 => n30546, ZN => n7524);
   U28844 : OAI222_X1 port map( A1 => n40976, A2 => n39875, B1 => n41360, B2 =>
                           n39868, C1 => n39866, C2 => n30545, ZN => n7523);
   U28845 : OAI222_X1 port map( A1 => n40952, A2 => n39855, B1 => n41336, B2 =>
                           n39848, C1 => n39846, C2 => n30485, ZN => n7463);
   U28846 : OAI222_X1 port map( A1 => n40964, A2 => n39855, B1 => n41348, B2 =>
                           n39848, C1 => n39846, C2 => n30483, ZN => n7461);
   U28847 : OAI222_X1 port map( A1 => n40970, A2 => n39855, B1 => n41354, B2 =>
                           n39848, C1 => n39846, C2 => n30482, ZN => n7460);
   U28848 : OAI222_X1 port map( A1 => n40976, A2 => n39855, B1 => n41360, B2 =>
                           n39848, C1 => n39846, C2 => n30481, ZN => n7459);
   U28849 : AOI221_X1 port map( B1 => n39162, B2 => n31109, C1 => n39156, C2 =>
                           n31173, A => n37024, ZN => n37023);
   U28850 : OAI222_X1 port map( A1 => n31291, A2 => n39150, B1 => n31355, B2 =>
                           n39144, C1 => n31227, C2 => n39138, ZN => n37024);
   U28851 : AOI221_X1 port map( B1 => n39163, B2 => n31108, C1 => n39157, C2 =>
                           n31172, A => n37005, ZN => n37004);
   U28852 : OAI222_X1 port map( A1 => n31290, A2 => n39151, B1 => n31354, B2 =>
                           n39145, C1 => n31226, C2 => n39139, ZN => n37005);
   U28853 : AOI221_X1 port map( B1 => n39163, B2 => n31107, C1 => n39157, C2 =>
                           n31171, A => n36986, ZN => n36985);
   U28854 : OAI222_X1 port map( A1 => n31289, A2 => n39151, B1 => n31353, B2 =>
                           n39145, C1 => n31225, C2 => n39139, ZN => n36986);
   U28855 : AOI221_X1 port map( B1 => n39163, B2 => n31106, C1 => n39157, C2 =>
                           n31170, A => n36967, ZN => n36966);
   U28856 : OAI222_X1 port map( A1 => n31288, A2 => n39151, B1 => n31352, B2 =>
                           n39145, C1 => n31224, C2 => n39139, ZN => n36967);
   U28857 : AOI221_X1 port map( B1 => n39163, B2 => n31105, C1 => n39157, C2 =>
                           n31169, A => n36948, ZN => n36947);
   U28858 : OAI222_X1 port map( A1 => n31287, A2 => n39151, B1 => n31351, B2 =>
                           n39145, C1 => n31223, C2 => n39139, ZN => n36948);
   U28859 : AOI221_X1 port map( B1 => n39163, B2 => n31104, C1 => n39157, C2 =>
                           n31168, A => n36929, ZN => n36928);
   U28860 : OAI222_X1 port map( A1 => n31286, A2 => n39151, B1 => n31350, B2 =>
                           n39145, C1 => n31222, C2 => n39139, ZN => n36929);
   U28861 : AOI221_X1 port map( B1 => n39163, B2 => n31103, C1 => n39157, C2 =>
                           n31167, A => n36910, ZN => n36909);
   U28862 : OAI222_X1 port map( A1 => n31285, A2 => n39151, B1 => n31349, B2 =>
                           n39145, C1 => n31221, C2 => n39139, ZN => n36910);
   U28863 : AOI221_X1 port map( B1 => n39163, B2 => n31102, C1 => n39157, C2 =>
                           n31166, A => n36891, ZN => n36890);
   U28864 : OAI222_X1 port map( A1 => n31284, A2 => n39151, B1 => n31348, B2 =>
                           n39145, C1 => n31220, C2 => n39139, ZN => n36891);
   U28865 : AOI221_X1 port map( B1 => n39163, B2 => n31101, C1 => n39157, C2 =>
                           n31165, A => n36872, ZN => n36871);
   U28866 : OAI222_X1 port map( A1 => n31283, A2 => n39151, B1 => n31347, B2 =>
                           n39145, C1 => n31219, C2 => n39139, ZN => n36872);
   U28867 : AOI221_X1 port map( B1 => n39163, B2 => n31100, C1 => n39157, C2 =>
                           n31164, A => n36853, ZN => n36852);
   U28868 : OAI222_X1 port map( A1 => n31282, A2 => n39151, B1 => n31346, B2 =>
                           n39145, C1 => n31218, C2 => n39139, ZN => n36853);
   U28869 : AOI221_X1 port map( B1 => n39163, B2 => n31099, C1 => n39157, C2 =>
                           n31163, A => n36834, ZN => n36833);
   U28870 : OAI222_X1 port map( A1 => n31281, A2 => n39151, B1 => n31345, B2 =>
                           n39145, C1 => n31217, C2 => n39139, ZN => n36834);
   U28871 : AOI221_X1 port map( B1 => n39163, B2 => n31098, C1 => n39157, C2 =>
                           n31162, A => n36815, ZN => n36814);
   U28872 : OAI222_X1 port map( A1 => n31280, A2 => n39151, B1 => n31344, B2 =>
                           n39145, C1 => n31216, C2 => n39139, ZN => n36815);
   U28873 : AOI221_X1 port map( B1 => n39163, B2 => n31097, C1 => n39157, C2 =>
                           n31161, A => n36796, ZN => n36795);
   U28874 : OAI222_X1 port map( A1 => n31279, A2 => n39151, B1 => n31343, B2 =>
                           n39145, C1 => n31215, C2 => n39139, ZN => n36796);
   U28875 : AOI221_X1 port map( B1 => n39164, B2 => n31096, C1 => n39158, C2 =>
                           n31160, A => n36777, ZN => n36776);
   U28876 : OAI222_X1 port map( A1 => n31278, A2 => n39152, B1 => n31342, B2 =>
                           n39146, C1 => n31214, C2 => n39140, ZN => n36777);
   U28877 : AOI221_X1 port map( B1 => n39164, B2 => n31095, C1 => n39158, C2 =>
                           n31159, A => n36758, ZN => n36757);
   U28878 : OAI222_X1 port map( A1 => n31277, A2 => n39152, B1 => n31341, B2 =>
                           n39146, C1 => n31213, C2 => n39140, ZN => n36758);
   U28879 : AOI221_X1 port map( B1 => n39164, B2 => n31094, C1 => n39158, C2 =>
                           n31158, A => n36739, ZN => n36738);
   U28880 : OAI222_X1 port map( A1 => n31276, A2 => n39152, B1 => n31340, B2 =>
                           n39146, C1 => n31212, C2 => n39140, ZN => n36739);
   U28881 : AOI221_X1 port map( B1 => n39164, B2 => n31093, C1 => n39158, C2 =>
                           n31157, A => n36720, ZN => n36719);
   U28882 : OAI222_X1 port map( A1 => n31275, A2 => n39152, B1 => n31339, B2 =>
                           n39146, C1 => n31211, C2 => n39140, ZN => n36720);
   U28883 : AOI221_X1 port map( B1 => n39164, B2 => n31092, C1 => n39158, C2 =>
                           n31156, A => n36701, ZN => n36700);
   U28884 : OAI222_X1 port map( A1 => n31274, A2 => n39152, B1 => n31338, B2 =>
                           n39146, C1 => n31210, C2 => n39140, ZN => n36701);
   U28885 : AOI221_X1 port map( B1 => n39164, B2 => n31091, C1 => n39158, C2 =>
                           n31155, A => n36682, ZN => n36681);
   U28886 : OAI222_X1 port map( A1 => n31273, A2 => n39152, B1 => n31337, B2 =>
                           n39146, C1 => n31209, C2 => n39140, ZN => n36682);
   U28887 : AOI221_X1 port map( B1 => n39164, B2 => n31090, C1 => n39158, C2 =>
                           n31154, A => n36663, ZN => n36662);
   U28888 : OAI222_X1 port map( A1 => n31272, A2 => n39152, B1 => n31336, B2 =>
                           n39146, C1 => n31208, C2 => n39140, ZN => n36663);
   U28889 : AOI221_X1 port map( B1 => n39164, B2 => n31089, C1 => n39158, C2 =>
                           n31153, A => n36644, ZN => n36643);
   U28890 : OAI222_X1 port map( A1 => n31271, A2 => n39152, B1 => n31335, B2 =>
                           n39146, C1 => n31207, C2 => n39140, ZN => n36644);
   U28891 : AOI221_X1 port map( B1 => n39164, B2 => n31088, C1 => n39158, C2 =>
                           n31152, A => n36625, ZN => n36624);
   U28892 : OAI222_X1 port map( A1 => n31270, A2 => n39152, B1 => n31334, B2 =>
                           n39146, C1 => n31206, C2 => n39140, ZN => n36625);
   U28893 : AOI221_X1 port map( B1 => n39164, B2 => n31087, C1 => n39158, C2 =>
                           n31151, A => n36606, ZN => n36605);
   U28894 : OAI222_X1 port map( A1 => n31269, A2 => n39152, B1 => n31333, B2 =>
                           n39146, C1 => n31205, C2 => n39140, ZN => n36606);
   U28895 : AOI221_X1 port map( B1 => n39164, B2 => n31086, C1 => n39158, C2 =>
                           n31150, A => n36587, ZN => n36586);
   U28896 : OAI222_X1 port map( A1 => n31268, A2 => n39152, B1 => n31332, B2 =>
                           n39146, C1 => n31204, C2 => n39140, ZN => n36587);
   U28897 : AOI221_X1 port map( B1 => n39164, B2 => n31085, C1 => n39158, C2 =>
                           n31149, A => n36568, ZN => n36567);
   U28898 : OAI222_X1 port map( A1 => n31267, A2 => n39152, B1 => n31331, B2 =>
                           n39146, C1 => n31203, C2 => n39140, ZN => n36568);
   U28899 : AOI221_X1 port map( B1 => n39165, B2 => n31084, C1 => n39159, C2 =>
                           n31148, A => n36549, ZN => n36548);
   U28900 : OAI222_X1 port map( A1 => n31266, A2 => n39153, B1 => n31330, B2 =>
                           n39147, C1 => n31202, C2 => n39141, ZN => n36549);
   U28901 : AOI221_X1 port map( B1 => n39165, B2 => n31083, C1 => n39159, C2 =>
                           n31147, A => n36530, ZN => n36529);
   U28902 : OAI222_X1 port map( A1 => n31265, A2 => n39153, B1 => n31329, B2 =>
                           n39147, C1 => n31201, C2 => n39141, ZN => n36530);
   U28903 : AOI221_X1 port map( B1 => n39165, B2 => n31082, C1 => n39159, C2 =>
                           n31146, A => n36511, ZN => n36510);
   U28904 : OAI222_X1 port map( A1 => n31264, A2 => n39153, B1 => n31328, B2 =>
                           n39147, C1 => n31200, C2 => n39141, ZN => n36511);
   U28905 : AOI221_X1 port map( B1 => n39165, B2 => n31081, C1 => n39159, C2 =>
                           n31145, A => n36492, ZN => n36491);
   U28906 : OAI222_X1 port map( A1 => n31263, A2 => n39153, B1 => n31327, B2 =>
                           n39147, C1 => n31199, C2 => n39141, ZN => n36492);
   U28907 : AOI221_X1 port map( B1 => n39165, B2 => n31080, C1 => n39159, C2 =>
                           n31144, A => n36473, ZN => n36472);
   U28908 : OAI222_X1 port map( A1 => n31262, A2 => n39153, B1 => n31326, B2 =>
                           n39147, C1 => n31198, C2 => n39141, ZN => n36473);
   U28909 : AOI221_X1 port map( B1 => n39165, B2 => n31079, C1 => n39159, C2 =>
                           n31143, A => n36454, ZN => n36453);
   U28910 : OAI222_X1 port map( A1 => n31261, A2 => n39153, B1 => n31325, B2 =>
                           n39147, C1 => n31197, C2 => n39141, ZN => n36454);
   U28911 : AOI221_X1 port map( B1 => n39165, B2 => n31078, C1 => n39159, C2 =>
                           n31142, A => n36435, ZN => n36434);
   U28912 : OAI222_X1 port map( A1 => n31260, A2 => n39153, B1 => n31324, B2 =>
                           n39147, C1 => n31196, C2 => n39141, ZN => n36435);
   U28913 : AOI221_X1 port map( B1 => n39165, B2 => n31077, C1 => n39159, C2 =>
                           n31141, A => n36416, ZN => n36415);
   U28914 : OAI222_X1 port map( A1 => n31259, A2 => n39153, B1 => n31323, B2 =>
                           n39147, C1 => n31195, C2 => n39141, ZN => n36416);
   U28915 : AOI221_X1 port map( B1 => n39165, B2 => n31076, C1 => n39159, C2 =>
                           n31140, A => n36397, ZN => n36396);
   U28916 : OAI222_X1 port map( A1 => n31258, A2 => n39153, B1 => n31322, B2 =>
                           n39147, C1 => n31194, C2 => n39141, ZN => n36397);
   U28917 : AOI221_X1 port map( B1 => n39165, B2 => n31075, C1 => n39159, C2 =>
                           n31139, A => n36378, ZN => n36377);
   U28918 : OAI222_X1 port map( A1 => n31257, A2 => n39153, B1 => n31321, B2 =>
                           n39147, C1 => n31193, C2 => n39141, ZN => n36378);
   U28919 : AOI221_X1 port map( B1 => n39165, B2 => n31074, C1 => n39159, C2 =>
                           n31138, A => n36359, ZN => n36358);
   U28920 : OAI222_X1 port map( A1 => n31256, A2 => n39153, B1 => n31320, B2 =>
                           n39147, C1 => n31192, C2 => n39141, ZN => n36359);
   U28921 : AOI221_X1 port map( B1 => n39165, B2 => n31073, C1 => n39159, C2 =>
                           n31137, A => n36340, ZN => n36339);
   U28922 : OAI222_X1 port map( A1 => n31255, A2 => n39153, B1 => n31319, B2 =>
                           n39147, C1 => n31191, C2 => n39141, ZN => n36340);
   U28923 : AOI221_X1 port map( B1 => n39166, B2 => n31072, C1 => n39160, C2 =>
                           n31136, A => n36321, ZN => n36320);
   U28924 : OAI222_X1 port map( A1 => n31254, A2 => n39154, B1 => n31318, B2 =>
                           n39148, C1 => n31190, C2 => n39142, ZN => n36321);
   U28925 : AOI221_X1 port map( B1 => n39166, B2 => n31071, C1 => n39160, C2 =>
                           n31135, A => n36302, ZN => n36301);
   U28926 : OAI222_X1 port map( A1 => n31253, A2 => n39154, B1 => n31317, B2 =>
                           n39148, C1 => n31189, C2 => n39142, ZN => n36302);
   U28927 : AOI221_X1 port map( B1 => n39166, B2 => n31070, C1 => n39160, C2 =>
                           n31134, A => n36283, ZN => n36282);
   U28928 : OAI222_X1 port map( A1 => n31252, A2 => n39154, B1 => n31316, B2 =>
                           n39148, C1 => n31188, C2 => n39142, ZN => n36283);
   U28929 : AOI221_X1 port map( B1 => n39166, B2 => n31069, C1 => n39160, C2 =>
                           n31133, A => n36264, ZN => n36263);
   U28930 : OAI222_X1 port map( A1 => n31251, A2 => n39154, B1 => n31315, B2 =>
                           n39148, C1 => n31187, C2 => n39142, ZN => n36264);
   U28931 : AOI221_X1 port map( B1 => n39166, B2 => n31068, C1 => n39160, C2 =>
                           n31132, A => n36245, ZN => n36244);
   U28932 : OAI222_X1 port map( A1 => n31250, A2 => n39154, B1 => n31314, B2 =>
                           n39148, C1 => n31186, C2 => n39142, ZN => n36245);
   U28933 : AOI221_X1 port map( B1 => n39166, B2 => n31067, C1 => n39160, C2 =>
                           n31131, A => n36226, ZN => n36225);
   U28934 : OAI222_X1 port map( A1 => n31249, A2 => n39154, B1 => n31313, B2 =>
                           n39148, C1 => n31185, C2 => n39142, ZN => n36226);
   U28935 : AOI221_X1 port map( B1 => n39167, B2 => n31060, C1 => n39161, C2 =>
                           n31124, A => n36093, ZN => n36092);
   U28936 : OAI222_X1 port map( A1 => n31242, A2 => n39155, B1 => n31306, B2 =>
                           n39149, C1 => n31178, C2 => n39143, ZN => n36093);
   U28937 : AOI221_X1 port map( B1 => n39167, B2 => n31059, C1 => n39161, C2 =>
                           n31123, A => n36074, ZN => n36073);
   U28938 : OAI222_X1 port map( A1 => n31241, A2 => n39155, B1 => n31305, B2 =>
                           n39149, C1 => n31177, C2 => n39143, ZN => n36074);
   U28939 : AOI221_X1 port map( B1 => n39167, B2 => n31058, C1 => n39161, C2 =>
                           n31122, A => n36055, ZN => n36054);
   U28940 : OAI222_X1 port map( A1 => n31240, A2 => n39155, B1 => n31304, B2 =>
                           n39149, C1 => n31176, C2 => n39143, ZN => n36055);
   U28941 : AOI221_X1 port map( B1 => n39167, B2 => n31057, C1 => n39161, C2 =>
                           n31121, A => n36018, ZN => n36015);
   U28942 : OAI222_X1 port map( A1 => n31239, A2 => n39155, B1 => n31303, B2 =>
                           n39149, C1 => n31175, C2 => n39143, ZN => n36018);
   U28943 : AOI221_X1 port map( B1 => n39162, B2 => n31110, C1 => n39156, C2 =>
                           n31174, A => n37043, ZN => n37042);
   U28944 : OAI222_X1 port map( A1 => n31292, A2 => n39150, B1 => n31356, B2 =>
                           n39144, C1 => n31228, C2 => n39138, ZN => n37043);
   U28945 : AOI221_X1 port map( B1 => n39166, B2 => n31066, C1 => n39160, C2 =>
                           n31130, A => n36207, ZN => n36206);
   U28946 : OAI222_X1 port map( A1 => n31248, A2 => n39154, B1 => n31312, B2 =>
                           n39148, C1 => n31184, C2 => n39142, ZN => n36207);
   U28947 : AOI221_X1 port map( B1 => n39166, B2 => n31065, C1 => n39160, C2 =>
                           n31129, A => n36188, ZN => n36187);
   U28948 : OAI222_X1 port map( A1 => n31247, A2 => n39154, B1 => n31311, B2 =>
                           n39148, C1 => n31183, C2 => n39142, ZN => n36188);
   U28949 : AOI221_X1 port map( B1 => n39166, B2 => n31064, C1 => n39160, C2 =>
                           n31128, A => n36169, ZN => n36168);
   U28950 : OAI222_X1 port map( A1 => n31246, A2 => n39154, B1 => n31310, B2 =>
                           n39148, C1 => n31182, C2 => n39142, ZN => n36169);
   U28951 : AOI221_X1 port map( B1 => n39166, B2 => n31063, C1 => n39160, C2 =>
                           n31127, A => n36150, ZN => n36149);
   U28952 : OAI222_X1 port map( A1 => n31245, A2 => n39154, B1 => n31309, B2 =>
                           n39148, C1 => n31181, C2 => n39142, ZN => n36150);
   U28953 : AOI221_X1 port map( B1 => n39166, B2 => n31062, C1 => n39160, C2 =>
                           n31126, A => n36131, ZN => n36130);
   U28954 : OAI222_X1 port map( A1 => n31244, A2 => n39154, B1 => n31308, B2 =>
                           n39148, C1 => n31180, C2 => n39142, ZN => n36131);
   U28955 : AOI221_X1 port map( B1 => n39166, B2 => n31061, C1 => n39160, C2 =>
                           n31125, A => n36112, ZN => n36111);
   U28956 : OAI222_X1 port map( A1 => n31243, A2 => n39154, B1 => n31307, B2 =>
                           n39148, C1 => n31179, C2 => n39142, ZN => n36112);
   U28957 : AOI221_X1 port map( B1 => n39668, B2 => n31110, C1 => n39662, C2 =>
                           n31174, A => n33671, ZN => n33670);
   U28958 : OAI222_X1 port map( A1 => n31292, A2 => n39656, B1 => n31356, B2 =>
                           n39650, C1 => n31228, C2 => n39644, ZN => n33671);
   U28959 : AOI221_X1 port map( B1 => n39416, B2 => n31110, C1 => n39410, C2 =>
                           n31174, A => n34945, ZN => n34944);
   U28960 : OAI222_X1 port map( A1 => n31292, A2 => n39404, B1 => n31356, B2 =>
                           n39398, C1 => n31228, C2 => n39392, ZN => n34945);
   U28961 : AOI221_X1 port map( B1 => n39668, B2 => n31109, C1 => n39662, C2 =>
                           n31173, A => n33690, ZN => n33689);
   U28962 : OAI222_X1 port map( A1 => n31291, A2 => n39656, B1 => n31355, B2 =>
                           n39650, C1 => n31227, C2 => n39644, ZN => n33690);
   U28963 : AOI221_X1 port map( B1 => n39416, B2 => n31109, C1 => n39410, C2 =>
                           n31173, A => n34964, ZN => n34963);
   U28964 : OAI222_X1 port map( A1 => n31291, A2 => n39404, B1 => n31355, B2 =>
                           n39398, C1 => n31227, C2 => n39392, ZN => n34964);
   U28965 : AOI221_X1 port map( B1 => n39668, B2 => n31108, C1 => n39662, C2 =>
                           n31172, A => n33709, ZN => n33708);
   U28966 : OAI222_X1 port map( A1 => n31290, A2 => n39656, B1 => n31354, B2 =>
                           n39650, C1 => n31226, C2 => n39644, ZN => n33709);
   U28967 : AOI221_X1 port map( B1 => n39416, B2 => n31108, C1 => n39410, C2 =>
                           n31172, A => n34983, ZN => n34982);
   U28968 : OAI222_X1 port map( A1 => n31290, A2 => n39404, B1 => n31354, B2 =>
                           n39398, C1 => n31226, C2 => n39392, ZN => n34983);
   U28969 : AOI221_X1 port map( B1 => n39668, B2 => n31107, C1 => n39662, C2 =>
                           n31171, A => n33728, ZN => n33727);
   U28970 : OAI222_X1 port map( A1 => n31289, A2 => n39656, B1 => n31353, B2 =>
                           n39650, C1 => n31225, C2 => n39644, ZN => n33728);
   U28971 : AOI221_X1 port map( B1 => n39416, B2 => n31107, C1 => n39410, C2 =>
                           n31171, A => n35002, ZN => n35001);
   U28972 : OAI222_X1 port map( A1 => n31289, A2 => n39404, B1 => n31353, B2 =>
                           n39398, C1 => n31225, C2 => n39392, ZN => n35002);
   U28973 : AOI221_X1 port map( B1 => n39668, B2 => n31106, C1 => n39662, C2 =>
                           n31170, A => n33747, ZN => n33746);
   U28974 : OAI222_X1 port map( A1 => n31288, A2 => n39656, B1 => n31352, B2 =>
                           n39650, C1 => n31224, C2 => n39644, ZN => n33747);
   U28975 : AOI221_X1 port map( B1 => n39416, B2 => n31106, C1 => n39410, C2 =>
                           n31170, A => n35021, ZN => n35020);
   U28976 : OAI222_X1 port map( A1 => n31288, A2 => n39404, B1 => n31352, B2 =>
                           n39398, C1 => n31224, C2 => n39392, ZN => n35021);
   U28977 : AOI221_X1 port map( B1 => n39668, B2 => n31105, C1 => n39662, C2 =>
                           n31169, A => n33766, ZN => n33765);
   U28978 : OAI222_X1 port map( A1 => n31287, A2 => n39656, B1 => n31351, B2 =>
                           n39650, C1 => n31223, C2 => n39644, ZN => n33766);
   U28979 : AOI221_X1 port map( B1 => n39416, B2 => n31105, C1 => n39410, C2 =>
                           n31169, A => n35040, ZN => n35039);
   U28980 : OAI222_X1 port map( A1 => n31287, A2 => n39404, B1 => n31351, B2 =>
                           n39398, C1 => n31223, C2 => n39392, ZN => n35040);
   U28981 : AOI221_X1 port map( B1 => n39667, B2 => n31104, C1 => n39661, C2 =>
                           n31168, A => n33785, ZN => n33784);
   U28982 : OAI222_X1 port map( A1 => n31286, A2 => n39655, B1 => n31350, B2 =>
                           n39649, C1 => n31222, C2 => n39643, ZN => n33785);
   U28983 : AOI221_X1 port map( B1 => n39415, B2 => n31104, C1 => n39409, C2 =>
                           n31168, A => n35059, ZN => n35058);
   U28984 : OAI222_X1 port map( A1 => n31286, A2 => n39403, B1 => n31350, B2 =>
                           n39397, C1 => n31222, C2 => n39391, ZN => n35059);
   U28985 : AOI221_X1 port map( B1 => n39667, B2 => n31103, C1 => n39661, C2 =>
                           n31167, A => n33804, ZN => n33803);
   U28986 : OAI222_X1 port map( A1 => n31285, A2 => n39655, B1 => n31349, B2 =>
                           n39649, C1 => n31221, C2 => n39643, ZN => n33804);
   U28987 : AOI221_X1 port map( B1 => n39415, B2 => n31103, C1 => n39409, C2 =>
                           n31167, A => n35078, ZN => n35077);
   U28988 : OAI222_X1 port map( A1 => n31285, A2 => n39403, B1 => n31349, B2 =>
                           n39397, C1 => n31221, C2 => n39391, ZN => n35078);
   U28989 : AOI221_X1 port map( B1 => n39667, B2 => n31102, C1 => n39661, C2 =>
                           n31166, A => n33823, ZN => n33822);
   U28990 : OAI222_X1 port map( A1 => n31284, A2 => n39655, B1 => n31348, B2 =>
                           n39649, C1 => n31220, C2 => n39643, ZN => n33823);
   U28991 : AOI221_X1 port map( B1 => n39415, B2 => n31102, C1 => n39409, C2 =>
                           n31166, A => n35097, ZN => n35096);
   U28992 : OAI222_X1 port map( A1 => n31284, A2 => n39403, B1 => n31348, B2 =>
                           n39397, C1 => n31220, C2 => n39391, ZN => n35097);
   U28993 : AOI221_X1 port map( B1 => n39667, B2 => n31101, C1 => n39661, C2 =>
                           n31165, A => n33842, ZN => n33841);
   U28994 : OAI222_X1 port map( A1 => n31283, A2 => n39655, B1 => n31347, B2 =>
                           n39649, C1 => n31219, C2 => n39643, ZN => n33842);
   U28995 : AOI221_X1 port map( B1 => n39415, B2 => n31101, C1 => n39409, C2 =>
                           n31165, A => n35116, ZN => n35115);
   U28996 : OAI222_X1 port map( A1 => n31283, A2 => n39403, B1 => n31347, B2 =>
                           n39397, C1 => n31219, C2 => n39391, ZN => n35116);
   U28997 : AOI221_X1 port map( B1 => n39667, B2 => n31100, C1 => n39661, C2 =>
                           n31164, A => n33861, ZN => n33860);
   U28998 : OAI222_X1 port map( A1 => n31282, A2 => n39655, B1 => n31346, B2 =>
                           n39649, C1 => n31218, C2 => n39643, ZN => n33861);
   U28999 : AOI221_X1 port map( B1 => n39415, B2 => n31100, C1 => n39409, C2 =>
                           n31164, A => n35135, ZN => n35134);
   U29000 : OAI222_X1 port map( A1 => n31282, A2 => n39403, B1 => n31346, B2 =>
                           n39397, C1 => n31218, C2 => n39391, ZN => n35135);
   U29001 : AOI221_X1 port map( B1 => n39667, B2 => n31099, C1 => n39661, C2 =>
                           n31163, A => n33880, ZN => n33879);
   U29002 : OAI222_X1 port map( A1 => n31281, A2 => n39655, B1 => n31345, B2 =>
                           n39649, C1 => n31217, C2 => n39643, ZN => n33880);
   U29003 : AOI221_X1 port map( B1 => n39415, B2 => n31099, C1 => n39409, C2 =>
                           n31163, A => n35154, ZN => n35153);
   U29004 : OAI222_X1 port map( A1 => n31281, A2 => n39403, B1 => n31345, B2 =>
                           n39397, C1 => n31217, C2 => n39391, ZN => n35154);
   U29005 : AOI221_X1 port map( B1 => n39667, B2 => n31098, C1 => n39661, C2 =>
                           n31162, A => n33899, ZN => n33898);
   U29006 : OAI222_X1 port map( A1 => n31280, A2 => n39655, B1 => n31344, B2 =>
                           n39649, C1 => n31216, C2 => n39643, ZN => n33899);
   U29007 : AOI221_X1 port map( B1 => n39415, B2 => n31098, C1 => n39409, C2 =>
                           n31162, A => n35173, ZN => n35172);
   U29008 : OAI222_X1 port map( A1 => n31280, A2 => n39403, B1 => n31344, B2 =>
                           n39397, C1 => n31216, C2 => n39391, ZN => n35173);
   U29009 : AOI221_X1 port map( B1 => n39667, B2 => n31097, C1 => n39661, C2 =>
                           n31161, A => n33918, ZN => n33917);
   U29010 : OAI222_X1 port map( A1 => n31279, A2 => n39655, B1 => n31343, B2 =>
                           n39649, C1 => n31215, C2 => n39643, ZN => n33918);
   U29011 : AOI221_X1 port map( B1 => n39415, B2 => n31097, C1 => n39409, C2 =>
                           n31161, A => n35192, ZN => n35191);
   U29012 : OAI222_X1 port map( A1 => n31279, A2 => n39403, B1 => n31343, B2 =>
                           n39397, C1 => n31215, C2 => n39391, ZN => n35192);
   U29013 : AOI221_X1 port map( B1 => n39667, B2 => n31096, C1 => n39661, C2 =>
                           n31160, A => n33937, ZN => n33936);
   U29014 : OAI222_X1 port map( A1 => n31278, A2 => n39655, B1 => n31342, B2 =>
                           n39649, C1 => n31214, C2 => n39643, ZN => n33937);
   U29015 : AOI221_X1 port map( B1 => n39415, B2 => n31096, C1 => n39409, C2 =>
                           n31160, A => n35211, ZN => n35210);
   U29016 : OAI222_X1 port map( A1 => n31278, A2 => n39403, B1 => n31342, B2 =>
                           n39397, C1 => n31214, C2 => n39391, ZN => n35211);
   U29017 : AOI221_X1 port map( B1 => n39667, B2 => n31095, C1 => n39661, C2 =>
                           n31159, A => n33956, ZN => n33955);
   U29018 : OAI222_X1 port map( A1 => n31277, A2 => n39655, B1 => n31341, B2 =>
                           n39649, C1 => n31213, C2 => n39643, ZN => n33956);
   U29019 : AOI221_X1 port map( B1 => n39415, B2 => n31095, C1 => n39409, C2 =>
                           n31159, A => n35230, ZN => n35229);
   U29020 : OAI222_X1 port map( A1 => n31277, A2 => n39403, B1 => n31341, B2 =>
                           n39397, C1 => n31213, C2 => n39391, ZN => n35230);
   U29021 : AOI221_X1 port map( B1 => n39667, B2 => n31094, C1 => n39661, C2 =>
                           n31158, A => n33975, ZN => n33974);
   U29022 : OAI222_X1 port map( A1 => n31276, A2 => n39655, B1 => n31340, B2 =>
                           n39649, C1 => n31212, C2 => n39643, ZN => n33975);
   U29023 : AOI221_X1 port map( B1 => n39415, B2 => n31094, C1 => n39409, C2 =>
                           n31158, A => n35249, ZN => n35248);
   U29024 : OAI222_X1 port map( A1 => n31276, A2 => n39403, B1 => n31340, B2 =>
                           n39397, C1 => n31212, C2 => n39391, ZN => n35249);
   U29025 : AOI221_X1 port map( B1 => n39667, B2 => n31093, C1 => n39661, C2 =>
                           n31157, A => n33994, ZN => n33993);
   U29026 : OAI222_X1 port map( A1 => n31275, A2 => n39655, B1 => n31339, B2 =>
                           n39649, C1 => n31211, C2 => n39643, ZN => n33994);
   U29027 : AOI221_X1 port map( B1 => n39415, B2 => n31093, C1 => n39409, C2 =>
                           n31157, A => n35268, ZN => n35267);
   U29028 : OAI222_X1 port map( A1 => n31275, A2 => n39403, B1 => n31339, B2 =>
                           n39397, C1 => n31211, C2 => n39391, ZN => n35268);
   U29029 : AOI221_X1 port map( B1 => n39666, B2 => n31092, C1 => n39660, C2 =>
                           n31156, A => n34013, ZN => n34012);
   U29030 : OAI222_X1 port map( A1 => n31274, A2 => n39654, B1 => n31338, B2 =>
                           n39648, C1 => n31210, C2 => n39642, ZN => n34013);
   U29031 : AOI221_X1 port map( B1 => n39414, B2 => n31092, C1 => n39408, C2 =>
                           n31156, A => n35287, ZN => n35286);
   U29032 : OAI222_X1 port map( A1 => n31274, A2 => n39402, B1 => n31338, B2 =>
                           n39396, C1 => n31210, C2 => n39390, ZN => n35287);
   U29033 : AOI221_X1 port map( B1 => n39666, B2 => n31091, C1 => n39660, C2 =>
                           n31155, A => n34032, ZN => n34031);
   U29034 : OAI222_X1 port map( A1 => n31273, A2 => n39654, B1 => n31337, B2 =>
                           n39648, C1 => n31209, C2 => n39642, ZN => n34032);
   U29035 : AOI221_X1 port map( B1 => n39414, B2 => n31091, C1 => n39408, C2 =>
                           n31155, A => n35306, ZN => n35305);
   U29036 : OAI222_X1 port map( A1 => n31273, A2 => n39402, B1 => n31337, B2 =>
                           n39396, C1 => n31209, C2 => n39390, ZN => n35306);
   U29037 : AOI221_X1 port map( B1 => n39666, B2 => n31090, C1 => n39660, C2 =>
                           n31154, A => n34051, ZN => n34050);
   U29038 : OAI222_X1 port map( A1 => n31272, A2 => n39654, B1 => n31336, B2 =>
                           n39648, C1 => n31208, C2 => n39642, ZN => n34051);
   U29039 : AOI221_X1 port map( B1 => n39414, B2 => n31090, C1 => n39408, C2 =>
                           n31154, A => n35325, ZN => n35324);
   U29040 : OAI222_X1 port map( A1 => n31272, A2 => n39402, B1 => n31336, B2 =>
                           n39396, C1 => n31208, C2 => n39390, ZN => n35325);
   U29041 : AOI221_X1 port map( B1 => n39666, B2 => n31089, C1 => n39660, C2 =>
                           n31153, A => n34070, ZN => n34069);
   U29042 : OAI222_X1 port map( A1 => n31271, A2 => n39654, B1 => n31335, B2 =>
                           n39648, C1 => n31207, C2 => n39642, ZN => n34070);
   U29043 : AOI221_X1 port map( B1 => n39414, B2 => n31089, C1 => n39408, C2 =>
                           n31153, A => n35344, ZN => n35343);
   U29044 : OAI222_X1 port map( A1 => n31271, A2 => n39402, B1 => n31335, B2 =>
                           n39396, C1 => n31207, C2 => n39390, ZN => n35344);
   U29045 : AOI221_X1 port map( B1 => n39666, B2 => n31088, C1 => n39660, C2 =>
                           n31152, A => n34089, ZN => n34088);
   U29046 : OAI222_X1 port map( A1 => n31270, A2 => n39654, B1 => n31334, B2 =>
                           n39648, C1 => n31206, C2 => n39642, ZN => n34089);
   U29047 : AOI221_X1 port map( B1 => n39414, B2 => n31088, C1 => n39408, C2 =>
                           n31152, A => n35363, ZN => n35362);
   U29048 : OAI222_X1 port map( A1 => n31270, A2 => n39402, B1 => n31334, B2 =>
                           n39396, C1 => n31206, C2 => n39390, ZN => n35363);
   U29049 : AOI221_X1 port map( B1 => n39666, B2 => n31087, C1 => n39660, C2 =>
                           n31151, A => n34108, ZN => n34107);
   U29050 : OAI222_X1 port map( A1 => n31269, A2 => n39654, B1 => n31333, B2 =>
                           n39648, C1 => n31205, C2 => n39642, ZN => n34108);
   U29051 : AOI221_X1 port map( B1 => n39414, B2 => n31087, C1 => n39408, C2 =>
                           n31151, A => n35382, ZN => n35381);
   U29052 : OAI222_X1 port map( A1 => n31269, A2 => n39402, B1 => n31333, B2 =>
                           n39396, C1 => n31205, C2 => n39390, ZN => n35382);
   U29053 : AOI221_X1 port map( B1 => n39666, B2 => n31086, C1 => n39660, C2 =>
                           n31150, A => n34127, ZN => n34126);
   U29054 : OAI222_X1 port map( A1 => n31268, A2 => n39654, B1 => n31332, B2 =>
                           n39648, C1 => n31204, C2 => n39642, ZN => n34127);
   U29055 : AOI221_X1 port map( B1 => n39414, B2 => n31086, C1 => n39408, C2 =>
                           n31150, A => n35401, ZN => n35400);
   U29056 : OAI222_X1 port map( A1 => n31268, A2 => n39402, B1 => n31332, B2 =>
                           n39396, C1 => n31204, C2 => n39390, ZN => n35401);
   U29057 : AOI221_X1 port map( B1 => n39666, B2 => n31085, C1 => n39660, C2 =>
                           n31149, A => n34146, ZN => n34145);
   U29058 : OAI222_X1 port map( A1 => n31267, A2 => n39654, B1 => n31331, B2 =>
                           n39648, C1 => n31203, C2 => n39642, ZN => n34146);
   U29059 : AOI221_X1 port map( B1 => n39414, B2 => n31085, C1 => n39408, C2 =>
                           n31149, A => n35420, ZN => n35419);
   U29060 : OAI222_X1 port map( A1 => n31267, A2 => n39402, B1 => n31331, B2 =>
                           n39396, C1 => n31203, C2 => n39390, ZN => n35420);
   U29061 : AOI221_X1 port map( B1 => n39666, B2 => n31084, C1 => n39660, C2 =>
                           n31148, A => n34165, ZN => n34164);
   U29062 : OAI222_X1 port map( A1 => n31266, A2 => n39654, B1 => n31330, B2 =>
                           n39648, C1 => n31202, C2 => n39642, ZN => n34165);
   U29063 : AOI221_X1 port map( B1 => n39414, B2 => n31084, C1 => n39408, C2 =>
                           n31148, A => n35439, ZN => n35438);
   U29064 : OAI222_X1 port map( A1 => n31266, A2 => n39402, B1 => n31330, B2 =>
                           n39396, C1 => n31202, C2 => n39390, ZN => n35439);
   U29065 : AOI221_X1 port map( B1 => n39666, B2 => n31083, C1 => n39660, C2 =>
                           n31147, A => n34184, ZN => n34183);
   U29066 : OAI222_X1 port map( A1 => n31265, A2 => n39654, B1 => n31329, B2 =>
                           n39648, C1 => n31201, C2 => n39642, ZN => n34184);
   U29067 : AOI221_X1 port map( B1 => n39414, B2 => n31083, C1 => n39408, C2 =>
                           n31147, A => n35458, ZN => n35457);
   U29068 : OAI222_X1 port map( A1 => n31265, A2 => n39402, B1 => n31329, B2 =>
                           n39396, C1 => n31201, C2 => n39390, ZN => n35458);
   U29069 : AOI221_X1 port map( B1 => n39666, B2 => n31082, C1 => n39660, C2 =>
                           n31146, A => n34203, ZN => n34202);
   U29070 : OAI222_X1 port map( A1 => n31264, A2 => n39654, B1 => n31328, B2 =>
                           n39648, C1 => n31200, C2 => n39642, ZN => n34203);
   U29071 : AOI221_X1 port map( B1 => n39414, B2 => n31082, C1 => n39408, C2 =>
                           n31146, A => n35477, ZN => n35476);
   U29072 : OAI222_X1 port map( A1 => n31264, A2 => n39402, B1 => n31328, B2 =>
                           n39396, C1 => n31200, C2 => n39390, ZN => n35477);
   U29073 : AOI221_X1 port map( B1 => n39666, B2 => n31081, C1 => n39660, C2 =>
                           n31145, A => n34222, ZN => n34221);
   U29074 : OAI222_X1 port map( A1 => n31263, A2 => n39654, B1 => n31327, B2 =>
                           n39648, C1 => n31199, C2 => n39642, ZN => n34222);
   U29075 : AOI221_X1 port map( B1 => n39414, B2 => n31081, C1 => n39408, C2 =>
                           n31145, A => n35496, ZN => n35495);
   U29076 : OAI222_X1 port map( A1 => n31263, A2 => n39402, B1 => n31327, B2 =>
                           n39396, C1 => n31199, C2 => n39390, ZN => n35496);
   U29077 : AOI221_X1 port map( B1 => n39665, B2 => n31080, C1 => n39659, C2 =>
                           n31144, A => n34241, ZN => n34240);
   U29078 : OAI222_X1 port map( A1 => n31262, A2 => n39653, B1 => n31326, B2 =>
                           n39647, C1 => n31198, C2 => n39641, ZN => n34241);
   U29079 : AOI221_X1 port map( B1 => n39413, B2 => n31080, C1 => n39407, C2 =>
                           n31144, A => n35515, ZN => n35514);
   U29080 : OAI222_X1 port map( A1 => n31262, A2 => n39401, B1 => n31326, B2 =>
                           n39395, C1 => n31198, C2 => n39389, ZN => n35515);
   U29081 : AOI221_X1 port map( B1 => n39665, B2 => n31079, C1 => n39659, C2 =>
                           n31143, A => n34260, ZN => n34259);
   U29082 : OAI222_X1 port map( A1 => n31261, A2 => n39653, B1 => n31325, B2 =>
                           n39647, C1 => n31197, C2 => n39641, ZN => n34260);
   U29083 : AOI221_X1 port map( B1 => n39413, B2 => n31079, C1 => n39407, C2 =>
                           n31143, A => n35534, ZN => n35533);
   U29084 : OAI222_X1 port map( A1 => n31261, A2 => n39401, B1 => n31325, B2 =>
                           n39395, C1 => n31197, C2 => n39389, ZN => n35534);
   U29085 : AOI221_X1 port map( B1 => n39665, B2 => n31078, C1 => n39659, C2 =>
                           n31142, A => n34279, ZN => n34278);
   U29086 : OAI222_X1 port map( A1 => n31260, A2 => n39653, B1 => n31324, B2 =>
                           n39647, C1 => n31196, C2 => n39641, ZN => n34279);
   U29087 : AOI221_X1 port map( B1 => n39413, B2 => n31078, C1 => n39407, C2 =>
                           n31142, A => n35553, ZN => n35552);
   U29088 : OAI222_X1 port map( A1 => n31260, A2 => n39401, B1 => n31324, B2 =>
                           n39395, C1 => n31196, C2 => n39389, ZN => n35553);
   U29089 : AOI221_X1 port map( B1 => n39665, B2 => n31077, C1 => n39659, C2 =>
                           n31141, A => n34298, ZN => n34297);
   U29090 : OAI222_X1 port map( A1 => n31259, A2 => n39653, B1 => n31323, B2 =>
                           n39647, C1 => n31195, C2 => n39641, ZN => n34298);
   U29091 : AOI221_X1 port map( B1 => n39413, B2 => n31077, C1 => n39407, C2 =>
                           n31141, A => n35572, ZN => n35571);
   U29092 : OAI222_X1 port map( A1 => n31259, A2 => n39401, B1 => n31323, B2 =>
                           n39395, C1 => n31195, C2 => n39389, ZN => n35572);
   U29093 : AOI221_X1 port map( B1 => n39665, B2 => n31076, C1 => n39659, C2 =>
                           n31140, A => n34317, ZN => n34316);
   U29094 : OAI222_X1 port map( A1 => n31258, A2 => n39653, B1 => n31322, B2 =>
                           n39647, C1 => n31194, C2 => n39641, ZN => n34317);
   U29095 : AOI221_X1 port map( B1 => n39413, B2 => n31076, C1 => n39407, C2 =>
                           n31140, A => n35591, ZN => n35590);
   U29096 : OAI222_X1 port map( A1 => n31258, A2 => n39401, B1 => n31322, B2 =>
                           n39395, C1 => n31194, C2 => n39389, ZN => n35591);
   U29097 : AOI221_X1 port map( B1 => n39665, B2 => n31075, C1 => n39659, C2 =>
                           n31139, A => n34336, ZN => n34335);
   U29098 : OAI222_X1 port map( A1 => n31257, A2 => n39653, B1 => n31321, B2 =>
                           n39647, C1 => n31193, C2 => n39641, ZN => n34336);
   U29099 : AOI221_X1 port map( B1 => n39413, B2 => n31075, C1 => n39407, C2 =>
                           n31139, A => n35610, ZN => n35609);
   U29100 : OAI222_X1 port map( A1 => n31257, A2 => n39401, B1 => n31321, B2 =>
                           n39395, C1 => n31193, C2 => n39389, ZN => n35610);
   U29101 : AOI221_X1 port map( B1 => n39665, B2 => n31074, C1 => n39659, C2 =>
                           n31138, A => n34355, ZN => n34354);
   U29102 : OAI222_X1 port map( A1 => n31256, A2 => n39653, B1 => n31320, B2 =>
                           n39647, C1 => n31192, C2 => n39641, ZN => n34355);
   U29103 : AOI221_X1 port map( B1 => n39413, B2 => n31074, C1 => n39407, C2 =>
                           n31138, A => n35629, ZN => n35628);
   U29104 : OAI222_X1 port map( A1 => n31256, A2 => n39401, B1 => n31320, B2 =>
                           n39395, C1 => n31192, C2 => n39389, ZN => n35629);
   U29105 : AOI221_X1 port map( B1 => n39665, B2 => n31073, C1 => n39659, C2 =>
                           n31137, A => n34374, ZN => n34373);
   U29106 : OAI222_X1 port map( A1 => n31255, A2 => n39653, B1 => n31319, B2 =>
                           n39647, C1 => n31191, C2 => n39641, ZN => n34374);
   U29107 : AOI221_X1 port map( B1 => n39413, B2 => n31073, C1 => n39407, C2 =>
                           n31137, A => n35648, ZN => n35647);
   U29108 : OAI222_X1 port map( A1 => n31255, A2 => n39401, B1 => n31319, B2 =>
                           n39395, C1 => n31191, C2 => n39389, ZN => n35648);
   U29109 : AOI221_X1 port map( B1 => n39665, B2 => n31072, C1 => n39659, C2 =>
                           n31136, A => n34393, ZN => n34392);
   U29110 : OAI222_X1 port map( A1 => n31254, A2 => n39653, B1 => n31318, B2 =>
                           n39647, C1 => n31190, C2 => n39641, ZN => n34393);
   U29111 : AOI221_X1 port map( B1 => n39413, B2 => n31072, C1 => n39407, C2 =>
                           n31136, A => n35667, ZN => n35666);
   U29112 : OAI222_X1 port map( A1 => n31254, A2 => n39401, B1 => n31318, B2 =>
                           n39395, C1 => n31190, C2 => n39389, ZN => n35667);
   U29113 : AOI221_X1 port map( B1 => n39665, B2 => n31071, C1 => n39659, C2 =>
                           n31135, A => n34412, ZN => n34411);
   U29114 : OAI222_X1 port map( A1 => n31253, A2 => n39653, B1 => n31317, B2 =>
                           n39647, C1 => n31189, C2 => n39641, ZN => n34412);
   U29115 : AOI221_X1 port map( B1 => n39413, B2 => n31071, C1 => n39407, C2 =>
                           n31135, A => n35686, ZN => n35685);
   U29116 : OAI222_X1 port map( A1 => n31253, A2 => n39401, B1 => n31317, B2 =>
                           n39395, C1 => n31189, C2 => n39389, ZN => n35686);
   U29117 : AOI221_X1 port map( B1 => n39665, B2 => n31070, C1 => n39659, C2 =>
                           n31134, A => n34431, ZN => n34430);
   U29118 : OAI222_X1 port map( A1 => n31252, A2 => n39653, B1 => n31316, B2 =>
                           n39647, C1 => n31188, C2 => n39641, ZN => n34431);
   U29119 : AOI221_X1 port map( B1 => n39413, B2 => n31070, C1 => n39407, C2 =>
                           n31134, A => n35705, ZN => n35704);
   U29120 : OAI222_X1 port map( A1 => n31252, A2 => n39401, B1 => n31316, B2 =>
                           n39395, C1 => n31188, C2 => n39389, ZN => n35705);
   U29121 : AOI221_X1 port map( B1 => n39665, B2 => n31069, C1 => n39659, C2 =>
                           n31133, A => n34450, ZN => n34449);
   U29122 : OAI222_X1 port map( A1 => n31251, A2 => n39653, B1 => n31315, B2 =>
                           n39647, C1 => n31187, C2 => n39641, ZN => n34450);
   U29123 : AOI221_X1 port map( B1 => n39413, B2 => n31069, C1 => n39407, C2 =>
                           n31133, A => n35724, ZN => n35723);
   U29124 : OAI222_X1 port map( A1 => n31251, A2 => n39401, B1 => n31315, B2 =>
                           n39395, C1 => n31187, C2 => n39389, ZN => n35724);
   U29125 : AOI221_X1 port map( B1 => n39664, B2 => n31068, C1 => n39658, C2 =>
                           n31132, A => n34469, ZN => n34468);
   U29126 : OAI222_X1 port map( A1 => n31250, A2 => n39652, B1 => n31314, B2 =>
                           n39646, C1 => n31186, C2 => n39640, ZN => n34469);
   U29127 : AOI221_X1 port map( B1 => n39412, B2 => n31068, C1 => n39406, C2 =>
                           n31132, A => n35743, ZN => n35742);
   U29128 : OAI222_X1 port map( A1 => n31250, A2 => n39400, B1 => n31314, B2 =>
                           n39394, C1 => n31186, C2 => n39388, ZN => n35743);
   U29129 : AOI221_X1 port map( B1 => n39664, B2 => n31067, C1 => n39658, C2 =>
                           n31131, A => n34488, ZN => n34487);
   U29130 : OAI222_X1 port map( A1 => n31249, A2 => n39652, B1 => n31313, B2 =>
                           n39646, C1 => n31185, C2 => n39640, ZN => n34488);
   U29131 : AOI221_X1 port map( B1 => n39412, B2 => n31067, C1 => n39406, C2 =>
                           n31131, A => n35762, ZN => n35761);
   U29132 : OAI222_X1 port map( A1 => n31249, A2 => n39400, B1 => n31313, B2 =>
                           n39394, C1 => n31185, C2 => n39388, ZN => n35762);
   U29133 : AOI221_X1 port map( B1 => n39664, B2 => n31066, C1 => n39658, C2 =>
                           n31130, A => n34507, ZN => n34506);
   U29134 : OAI222_X1 port map( A1 => n31248, A2 => n39652, B1 => n31312, B2 =>
                           n39646, C1 => n31184, C2 => n39640, ZN => n34507);
   U29135 : AOI221_X1 port map( B1 => n39412, B2 => n31066, C1 => n39406, C2 =>
                           n31130, A => n35781, ZN => n35780);
   U29136 : OAI222_X1 port map( A1 => n31248, A2 => n39400, B1 => n31312, B2 =>
                           n39394, C1 => n31184, C2 => n39388, ZN => n35781);
   U29137 : AOI221_X1 port map( B1 => n39664, B2 => n31065, C1 => n39658, C2 =>
                           n31129, A => n34526, ZN => n34525);
   U29138 : OAI222_X1 port map( A1 => n31247, A2 => n39652, B1 => n31311, B2 =>
                           n39646, C1 => n31183, C2 => n39640, ZN => n34526);
   U29139 : AOI221_X1 port map( B1 => n39412, B2 => n31065, C1 => n39406, C2 =>
                           n31129, A => n35800, ZN => n35799);
   U29140 : OAI222_X1 port map( A1 => n31247, A2 => n39400, B1 => n31311, B2 =>
                           n39394, C1 => n31183, C2 => n39388, ZN => n35800);
   U29141 : AOI221_X1 port map( B1 => n39664, B2 => n31064, C1 => n39658, C2 =>
                           n31128, A => n34545, ZN => n34544);
   U29142 : OAI222_X1 port map( A1 => n31246, A2 => n39652, B1 => n31310, B2 =>
                           n39646, C1 => n31182, C2 => n39640, ZN => n34545);
   U29143 : AOI221_X1 port map( B1 => n39412, B2 => n31064, C1 => n39406, C2 =>
                           n31128, A => n35819, ZN => n35818);
   U29144 : OAI222_X1 port map( A1 => n31246, A2 => n39400, B1 => n31310, B2 =>
                           n39394, C1 => n31182, C2 => n39388, ZN => n35819);
   U29145 : AOI221_X1 port map( B1 => n39664, B2 => n31063, C1 => n39658, C2 =>
                           n31127, A => n34564, ZN => n34563);
   U29146 : OAI222_X1 port map( A1 => n31245, A2 => n39652, B1 => n31309, B2 =>
                           n39646, C1 => n31181, C2 => n39640, ZN => n34564);
   U29147 : AOI221_X1 port map( B1 => n39412, B2 => n31063, C1 => n39406, C2 =>
                           n31127, A => n35838, ZN => n35837);
   U29148 : OAI222_X1 port map( A1 => n31245, A2 => n39400, B1 => n31309, B2 =>
                           n39394, C1 => n31181, C2 => n39388, ZN => n35838);
   U29149 : AOI221_X1 port map( B1 => n39664, B2 => n31062, C1 => n39658, C2 =>
                           n31126, A => n34583, ZN => n34582);
   U29150 : OAI222_X1 port map( A1 => n31244, A2 => n39652, B1 => n31308, B2 =>
                           n39646, C1 => n31180, C2 => n39640, ZN => n34583);
   U29151 : AOI221_X1 port map( B1 => n39412, B2 => n31062, C1 => n39406, C2 =>
                           n31126, A => n35857, ZN => n35856);
   U29152 : OAI222_X1 port map( A1 => n31244, A2 => n39400, B1 => n31308, B2 =>
                           n39394, C1 => n31180, C2 => n39388, ZN => n35857);
   U29153 : AOI221_X1 port map( B1 => n39664, B2 => n31061, C1 => n39658, C2 =>
                           n31125, A => n34602, ZN => n34601);
   U29154 : OAI222_X1 port map( A1 => n31243, A2 => n39652, B1 => n31307, B2 =>
                           n39646, C1 => n31179, C2 => n39640, ZN => n34602);
   U29155 : AOI221_X1 port map( B1 => n39412, B2 => n31061, C1 => n39406, C2 =>
                           n31125, A => n35876, ZN => n35875);
   U29156 : OAI222_X1 port map( A1 => n31243, A2 => n39400, B1 => n31307, B2 =>
                           n39394, C1 => n31179, C2 => n39388, ZN => n35876);
   U29157 : AOI221_X1 port map( B1 => n39664, B2 => n31060, C1 => n39658, C2 =>
                           n31124, A => n34621, ZN => n34620);
   U29158 : OAI222_X1 port map( A1 => n31242, A2 => n39652, B1 => n31306, B2 =>
                           n39646, C1 => n31178, C2 => n39640, ZN => n34621);
   U29159 : AOI221_X1 port map( B1 => n39412, B2 => n31060, C1 => n39406, C2 =>
                           n31124, A => n35895, ZN => n35894);
   U29160 : OAI222_X1 port map( A1 => n31242, A2 => n39400, B1 => n31306, B2 =>
                           n39394, C1 => n31178, C2 => n39388, ZN => n35895);
   U29161 : AOI221_X1 port map( B1 => n39664, B2 => n31059, C1 => n39658, C2 =>
                           n31123, A => n34640, ZN => n34639);
   U29162 : OAI222_X1 port map( A1 => n31241, A2 => n39652, B1 => n31305, B2 =>
                           n39646, C1 => n31177, C2 => n39640, ZN => n34640);
   U29163 : AOI221_X1 port map( B1 => n39412, B2 => n31059, C1 => n39406, C2 =>
                           n31123, A => n35914, ZN => n35913);
   U29164 : OAI222_X1 port map( A1 => n31241, A2 => n39400, B1 => n31305, B2 =>
                           n39394, C1 => n31177, C2 => n39388, ZN => n35914);
   U29165 : AOI221_X1 port map( B1 => n39664, B2 => n31058, C1 => n39658, C2 =>
                           n31122, A => n34659, ZN => n34658);
   U29166 : OAI222_X1 port map( A1 => n31240, A2 => n39652, B1 => n31304, B2 =>
                           n39646, C1 => n31176, C2 => n39640, ZN => n34659);
   U29167 : AOI221_X1 port map( B1 => n39412, B2 => n31058, C1 => n39406, C2 =>
                           n31122, A => n35933, ZN => n35932);
   U29168 : OAI222_X1 port map( A1 => n31240, A2 => n39400, B1 => n31304, B2 =>
                           n39394, C1 => n31176, C2 => n39388, ZN => n35933);
   U29169 : AOI221_X1 port map( B1 => n39664, B2 => n31057, C1 => n39658, C2 =>
                           n31121, A => n34689, ZN => n34688);
   U29170 : OAI222_X1 port map( A1 => n31239, A2 => n39652, B1 => n31303, B2 =>
                           n39646, C1 => n31175, C2 => n39640, ZN => n34689);
   U29171 : AOI221_X1 port map( B1 => n39412, B2 => n31057, C1 => n39406, C2 =>
                           n31121, A => n35963, ZN => n35962);
   U29172 : OAI222_X1 port map( A1 => n31239, A2 => n39400, B1 => n31303, B2 =>
                           n39394, C1 => n31175, C2 => n39388, ZN => n35963);
   U29173 : AOI221_X1 port map( B1 => n39132, B2 => n32815, C1 => n39126, C2 =>
                           n32767, A => n37025, ZN => n37022);
   U29174 : OAI222_X1 port map( A1 => n30981, A2 => n39120, B1 => n31045, B2 =>
                           n39114, C1 => n30917, C2 => n39108, ZN => n37025);
   U29175 : AOI221_X1 port map( B1 => n39133, B2 => n32814, C1 => n39127, C2 =>
                           n32766, A => n37006, ZN => n37003);
   U29176 : OAI222_X1 port map( A1 => n30980, A2 => n39121, B1 => n31044, B2 =>
                           n39115, C1 => n30916, C2 => n39109, ZN => n37006);
   U29177 : AOI221_X1 port map( B1 => n39133, B2 => n32813, C1 => n39127, C2 =>
                           n32765, A => n36987, ZN => n36984);
   U29178 : OAI222_X1 port map( A1 => n30979, A2 => n39121, B1 => n31043, B2 =>
                           n39115, C1 => n30915, C2 => n39109, ZN => n36987);
   U29179 : AOI221_X1 port map( B1 => n39133, B2 => n32812, C1 => n39127, C2 =>
                           n32764, A => n36968, ZN => n36965);
   U29180 : OAI222_X1 port map( A1 => n30978, A2 => n39121, B1 => n31042, B2 =>
                           n39115, C1 => n30914, C2 => n39109, ZN => n36968);
   U29181 : AOI221_X1 port map( B1 => n39133, B2 => n32811, C1 => n39127, C2 =>
                           n32763, A => n36949, ZN => n36946);
   U29182 : OAI222_X1 port map( A1 => n30977, A2 => n39121, B1 => n31041, B2 =>
                           n39115, C1 => n30913, C2 => n39109, ZN => n36949);
   U29183 : AOI221_X1 port map( B1 => n39133, B2 => n32810, C1 => n39127, C2 =>
                           n32762, A => n36930, ZN => n36927);
   U29184 : OAI222_X1 port map( A1 => n30976, A2 => n39121, B1 => n31040, B2 =>
                           n39115, C1 => n30912, C2 => n39109, ZN => n36930);
   U29185 : AOI221_X1 port map( B1 => n39133, B2 => n32809, C1 => n39127, C2 =>
                           n32761, A => n36911, ZN => n36908);
   U29186 : OAI222_X1 port map( A1 => n30975, A2 => n39121, B1 => n31039, B2 =>
                           n39115, C1 => n30911, C2 => n39109, ZN => n36911);
   U29187 : AOI221_X1 port map( B1 => n39133, B2 => n32808, C1 => n39127, C2 =>
                           n32760, A => n36892, ZN => n36889);
   U29188 : OAI222_X1 port map( A1 => n30974, A2 => n39121, B1 => n31038, B2 =>
                           n39115, C1 => n30910, C2 => n39109, ZN => n36892);
   U29189 : AOI221_X1 port map( B1 => n39133, B2 => n32807, C1 => n39127, C2 =>
                           n32759, A => n36873, ZN => n36870);
   U29190 : OAI222_X1 port map( A1 => n30973, A2 => n39121, B1 => n31037, B2 =>
                           n39115, C1 => n30909, C2 => n39109, ZN => n36873);
   U29191 : AOI221_X1 port map( B1 => n39133, B2 => n32806, C1 => n39127, C2 =>
                           n32758, A => n36854, ZN => n36851);
   U29192 : OAI222_X1 port map( A1 => n30972, A2 => n39121, B1 => n31036, B2 =>
                           n39115, C1 => n30908, C2 => n39109, ZN => n36854);
   U29193 : AOI221_X1 port map( B1 => n39133, B2 => n32805, C1 => n39127, C2 =>
                           n32757, A => n36835, ZN => n36832);
   U29194 : OAI222_X1 port map( A1 => n30971, A2 => n39121, B1 => n31035, B2 =>
                           n39115, C1 => n30907, C2 => n39109, ZN => n36835);
   U29195 : AOI221_X1 port map( B1 => n39133, B2 => n32804, C1 => n39127, C2 =>
                           n32756, A => n36816, ZN => n36813);
   U29196 : OAI222_X1 port map( A1 => n30970, A2 => n39121, B1 => n31034, B2 =>
                           n39115, C1 => n30906, C2 => n39109, ZN => n36816);
   U29197 : AOI221_X1 port map( B1 => n39133, B2 => n32803, C1 => n39127, C2 =>
                           n32755, A => n36797, ZN => n36794);
   U29198 : OAI222_X1 port map( A1 => n30969, A2 => n39121, B1 => n31033, B2 =>
                           n39115, C1 => n30905, C2 => n39109, ZN => n36797);
   U29199 : AOI221_X1 port map( B1 => n39134, B2 => n32802, C1 => n39128, C2 =>
                           n32754, A => n36778, ZN => n36775);
   U29200 : OAI222_X1 port map( A1 => n30968, A2 => n39122, B1 => n31032, B2 =>
                           n39116, C1 => n30904, C2 => n39110, ZN => n36778);
   U29201 : AOI221_X1 port map( B1 => n39134, B2 => n32801, C1 => n39128, C2 =>
                           n32753, A => n36759, ZN => n36756);
   U29202 : OAI222_X1 port map( A1 => n30967, A2 => n39122, B1 => n31031, B2 =>
                           n39116, C1 => n30903, C2 => n39110, ZN => n36759);
   U29203 : AOI221_X1 port map( B1 => n39134, B2 => n32800, C1 => n39128, C2 =>
                           n32752, A => n36740, ZN => n36737);
   U29204 : OAI222_X1 port map( A1 => n30966, A2 => n39122, B1 => n31030, B2 =>
                           n39116, C1 => n30902, C2 => n39110, ZN => n36740);
   U29205 : AOI221_X1 port map( B1 => n39134, B2 => n32799, C1 => n39128, C2 =>
                           n32751, A => n36721, ZN => n36718);
   U29206 : OAI222_X1 port map( A1 => n30965, A2 => n39122, B1 => n31029, B2 =>
                           n39116, C1 => n30901, C2 => n39110, ZN => n36721);
   U29207 : AOI221_X1 port map( B1 => n39134, B2 => n32798, C1 => n39128, C2 =>
                           n32750, A => n36702, ZN => n36699);
   U29208 : OAI222_X1 port map( A1 => n30964, A2 => n39122, B1 => n31028, B2 =>
                           n39116, C1 => n30900, C2 => n39110, ZN => n36702);
   U29209 : AOI221_X1 port map( B1 => n39134, B2 => n32797, C1 => n39128, C2 =>
                           n32749, A => n36683, ZN => n36680);
   U29210 : OAI222_X1 port map( A1 => n30963, A2 => n39122, B1 => n31027, B2 =>
                           n39116, C1 => n30899, C2 => n39110, ZN => n36683);
   U29211 : AOI221_X1 port map( B1 => n39134, B2 => n32796, C1 => n39128, C2 =>
                           n32748, A => n36664, ZN => n36661);
   U29212 : OAI222_X1 port map( A1 => n30962, A2 => n39122, B1 => n31026, B2 =>
                           n39116, C1 => n30898, C2 => n39110, ZN => n36664);
   U29213 : AOI221_X1 port map( B1 => n39134, B2 => n32795, C1 => n39128, C2 =>
                           n32747, A => n36645, ZN => n36642);
   U29214 : OAI222_X1 port map( A1 => n30961, A2 => n39122, B1 => n31025, B2 =>
                           n39116, C1 => n30897, C2 => n39110, ZN => n36645);
   U29215 : AOI221_X1 port map( B1 => n39134, B2 => n32794, C1 => n39128, C2 =>
                           n32746, A => n36626, ZN => n36623);
   U29216 : OAI222_X1 port map( A1 => n30960, A2 => n39122, B1 => n31024, B2 =>
                           n39116, C1 => n30896, C2 => n39110, ZN => n36626);
   U29217 : AOI221_X1 port map( B1 => n39134, B2 => n32793, C1 => n39128, C2 =>
                           n32745, A => n36607, ZN => n36604);
   U29218 : OAI222_X1 port map( A1 => n30959, A2 => n39122, B1 => n31023, B2 =>
                           n39116, C1 => n30895, C2 => n39110, ZN => n36607);
   U29219 : AOI221_X1 port map( B1 => n39134, B2 => n32792, C1 => n39128, C2 =>
                           n32744, A => n36588, ZN => n36585);
   U29220 : OAI222_X1 port map( A1 => n30958, A2 => n39122, B1 => n31022, B2 =>
                           n39116, C1 => n30894, C2 => n39110, ZN => n36588);
   U29221 : AOI221_X1 port map( B1 => n39134, B2 => n32791, C1 => n39128, C2 =>
                           n32743, A => n36569, ZN => n36566);
   U29222 : OAI222_X1 port map( A1 => n30957, A2 => n39122, B1 => n31021, B2 =>
                           n39116, C1 => n30893, C2 => n39110, ZN => n36569);
   U29223 : AOI221_X1 port map( B1 => n39135, B2 => n32790, C1 => n39129, C2 =>
                           n32742, A => n36550, ZN => n36547);
   U29224 : OAI222_X1 port map( A1 => n30956, A2 => n39123, B1 => n31020, B2 =>
                           n39117, C1 => n30892, C2 => n39111, ZN => n36550);
   U29225 : AOI221_X1 port map( B1 => n39135, B2 => n32789, C1 => n39129, C2 =>
                           n32741, A => n36531, ZN => n36528);
   U29226 : OAI222_X1 port map( A1 => n30955, A2 => n39123, B1 => n31019, B2 =>
                           n39117, C1 => n30891, C2 => n39111, ZN => n36531);
   U29227 : AOI221_X1 port map( B1 => n39135, B2 => n32788, C1 => n39129, C2 =>
                           n32740, A => n36512, ZN => n36509);
   U29228 : OAI222_X1 port map( A1 => n30954, A2 => n39123, B1 => n31018, B2 =>
                           n39117, C1 => n30890, C2 => n39111, ZN => n36512);
   U29229 : AOI221_X1 port map( B1 => n39135, B2 => n32787, C1 => n39129, C2 =>
                           n32739, A => n36493, ZN => n36490);
   U29230 : OAI222_X1 port map( A1 => n30953, A2 => n39123, B1 => n31017, B2 =>
                           n39117, C1 => n30889, C2 => n39111, ZN => n36493);
   U29231 : AOI221_X1 port map( B1 => n39135, B2 => n32786, C1 => n39129, C2 =>
                           n32738, A => n36474, ZN => n36471);
   U29232 : OAI222_X1 port map( A1 => n30952, A2 => n39123, B1 => n31016, B2 =>
                           n39117, C1 => n30888, C2 => n39111, ZN => n36474);
   U29233 : AOI221_X1 port map( B1 => n39135, B2 => n32785, C1 => n39129, C2 =>
                           n32737, A => n36455, ZN => n36452);
   U29234 : OAI222_X1 port map( A1 => n30951, A2 => n39123, B1 => n31015, B2 =>
                           n39117, C1 => n30887, C2 => n39111, ZN => n36455);
   U29235 : AOI221_X1 port map( B1 => n39135, B2 => n32784, C1 => n39129, C2 =>
                           n32736, A => n36436, ZN => n36433);
   U29236 : OAI222_X1 port map( A1 => n30950, A2 => n39123, B1 => n31014, B2 =>
                           n39117, C1 => n30886, C2 => n39111, ZN => n36436);
   U29237 : AOI221_X1 port map( B1 => n39135, B2 => n32783, C1 => n39129, C2 =>
                           n32735, A => n36417, ZN => n36414);
   U29238 : OAI222_X1 port map( A1 => n30949, A2 => n39123, B1 => n31013, B2 =>
                           n39117, C1 => n30885, C2 => n39111, ZN => n36417);
   U29239 : AOI221_X1 port map( B1 => n39135, B2 => n32782, C1 => n39129, C2 =>
                           n32734, A => n36398, ZN => n36395);
   U29240 : OAI222_X1 port map( A1 => n30948, A2 => n39123, B1 => n31012, B2 =>
                           n39117, C1 => n30884, C2 => n39111, ZN => n36398);
   U29241 : AOI221_X1 port map( B1 => n39135, B2 => n32781, C1 => n39129, C2 =>
                           n32733, A => n36379, ZN => n36376);
   U29242 : OAI222_X1 port map( A1 => n30947, A2 => n39123, B1 => n31011, B2 =>
                           n39117, C1 => n30883, C2 => n39111, ZN => n36379);
   U29243 : AOI221_X1 port map( B1 => n39135, B2 => n32780, C1 => n39129, C2 =>
                           n32732, A => n36360, ZN => n36357);
   U29244 : OAI222_X1 port map( A1 => n30946, A2 => n39123, B1 => n31010, B2 =>
                           n39117, C1 => n30882, C2 => n39111, ZN => n36360);
   U29245 : AOI221_X1 port map( B1 => n39135, B2 => n32779, C1 => n39129, C2 =>
                           n32731, A => n36341, ZN => n36338);
   U29246 : OAI222_X1 port map( A1 => n30945, A2 => n39123, B1 => n31009, B2 =>
                           n39117, C1 => n30881, C2 => n39111, ZN => n36341);
   U29247 : AOI221_X1 port map( B1 => n39136, B2 => n32778, C1 => n39130, C2 =>
                           n32730, A => n36322, ZN => n36319);
   U29248 : OAI222_X1 port map( A1 => n30944, A2 => n39124, B1 => n31008, B2 =>
                           n39118, C1 => n30880, C2 => n39112, ZN => n36322);
   U29249 : AOI221_X1 port map( B1 => n39136, B2 => n32777, C1 => n39130, C2 =>
                           n32729, A => n36303, ZN => n36300);
   U29250 : OAI222_X1 port map( A1 => n30943, A2 => n39124, B1 => n31007, B2 =>
                           n39118, C1 => n30879, C2 => n39112, ZN => n36303);
   U29251 : AOI221_X1 port map( B1 => n39136, B2 => n32776, C1 => n39130, C2 =>
                           n32728, A => n36284, ZN => n36281);
   U29252 : OAI222_X1 port map( A1 => n30942, A2 => n39124, B1 => n31006, B2 =>
                           n39118, C1 => n30878, C2 => n39112, ZN => n36284);
   U29253 : AOI221_X1 port map( B1 => n39136, B2 => n32775, C1 => n39130, C2 =>
                           n32727, A => n36265, ZN => n36262);
   U29254 : OAI222_X1 port map( A1 => n30941, A2 => n39124, B1 => n31005, B2 =>
                           n39118, C1 => n30877, C2 => n39112, ZN => n36265);
   U29255 : AOI221_X1 port map( B1 => n39136, B2 => n32846, C1 => n39130, C2 =>
                           n32834, A => n36246, ZN => n36243);
   U29256 : OAI222_X1 port map( A1 => n30940, A2 => n39124, B1 => n31004, B2 =>
                           n39118, C1 => n30876, C2 => n39112, ZN => n36246);
   U29257 : AOI221_X1 port map( B1 => n39136, B2 => n32845, C1 => n39130, C2 =>
                           n32833, A => n36227, ZN => n36224);
   U29258 : OAI222_X1 port map( A1 => n30939, A2 => n39124, B1 => n31003, B2 =>
                           n39118, C1 => n30875, C2 => n39112, ZN => n36227);
   U29259 : AOI221_X1 port map( B1 => n39132, B2 => n32474, C1 => n39126, C2 =>
                           n32470, A => n37215, ZN => n37212);
   U29260 : OAI222_X1 port map( A1 => n30991, A2 => n39120, B1 => n31055, B2 =>
                           n39114, C1 => n30927, C2 => n39108, ZN => n37215);
   U29261 : AOI221_X1 port map( B1 => n39132, B2 => n32473, C1 => n39126, C2 =>
                           n32469, A => n37196, ZN => n37193);
   U29262 : OAI222_X1 port map( A1 => n30990, A2 => n39120, B1 => n31054, B2 =>
                           n39114, C1 => n30926, C2 => n39108, ZN => n37196);
   U29263 : AOI221_X1 port map( B1 => n39132, B2 => n32472, C1 => n39126, C2 =>
                           n32468, A => n37177, ZN => n37174);
   U29264 : OAI222_X1 port map( A1 => n30989, A2 => n39120, B1 => n31053, B2 =>
                           n39114, C1 => n30925, C2 => n39108, ZN => n37177);
   U29265 : AOI221_X1 port map( B1 => n39132, B2 => n32822, C1 => n39126, C2 =>
                           n32774, A => n37158, ZN => n37155);
   U29266 : OAI222_X1 port map( A1 => n30988, A2 => n39120, B1 => n31052, B2 =>
                           n39114, C1 => n30924, C2 => n39108, ZN => n37158);
   U29267 : AOI221_X1 port map( B1 => n39132, B2 => n32821, C1 => n39126, C2 =>
                           n32773, A => n37139, ZN => n37136);
   U29268 : OAI222_X1 port map( A1 => n30987, A2 => n39120, B1 => n31051, B2 =>
                           n39114, C1 => n30923, C2 => n39108, ZN => n37139);
   U29269 : AOI221_X1 port map( B1 => n39137, B2 => n32838, C1 => n39131, C2 =>
                           n32826, A => n36094, ZN => n36091);
   U29270 : OAI222_X1 port map( A1 => n30932, A2 => n39125, B1 => n30996, B2 =>
                           n39119, C1 => n30868, C2 => n39113, ZN => n36094);
   U29271 : AOI221_X1 port map( B1 => n39137, B2 => n32837, C1 => n39131, C2 =>
                           n32825, A => n36075, ZN => n36072);
   U29272 : OAI222_X1 port map( A1 => n30931, A2 => n39125, B1 => n30995, B2 =>
                           n39119, C1 => n30867, C2 => n39113, ZN => n36075);
   U29273 : AOI221_X1 port map( B1 => n39137, B2 => n32836, C1 => n39131, C2 =>
                           n32824, A => n36056, ZN => n36053);
   U29274 : OAI222_X1 port map( A1 => n30930, A2 => n39125, B1 => n30994, B2 =>
                           n39119, C1 => n30866, C2 => n39113, ZN => n36056);
   U29275 : AOI221_X1 port map( B1 => n39137, B2 => n32835, C1 => n39131, C2 =>
                           n32823, A => n36024, ZN => n36014);
   U29276 : OAI222_X1 port map( A1 => n30929, A2 => n39125, B1 => n30993, B2 =>
                           n39119, C1 => n30865, C2 => n39113, ZN => n36024);
   U29277 : AOI221_X1 port map( B1 => n39132, B2 => n32475, C1 => n39126, C2 =>
                           n32471, A => n37247, ZN => n37243);
   U29278 : OAI222_X1 port map( A1 => n30992, A2 => n39120, B1 => n31056, B2 =>
                           n39114, C1 => n30928, C2 => n39108, ZN => n37247);
   U29279 : AOI221_X1 port map( B1 => n39132, B2 => n32820, C1 => n39126, C2 =>
                           n32772, A => n37120, ZN => n37117);
   U29280 : OAI222_X1 port map( A1 => n30986, A2 => n39120, B1 => n31050, B2 =>
                           n39114, C1 => n30922, C2 => n39108, ZN => n37120);
   U29281 : AOI221_X1 port map( B1 => n39132, B2 => n32819, C1 => n39126, C2 =>
                           n32771, A => n37101, ZN => n37098);
   U29282 : OAI222_X1 port map( A1 => n30985, A2 => n39120, B1 => n31049, B2 =>
                           n39114, C1 => n30921, C2 => n39108, ZN => n37101);
   U29283 : AOI221_X1 port map( B1 => n39132, B2 => n32818, C1 => n39126, C2 =>
                           n32770, A => n37082, ZN => n37079);
   U29284 : OAI222_X1 port map( A1 => n30984, A2 => n39120, B1 => n31048, B2 =>
                           n39114, C1 => n30920, C2 => n39108, ZN => n37082);
   U29285 : AOI221_X1 port map( B1 => n39132, B2 => n32817, C1 => n39126, C2 =>
                           n32769, A => n37063, ZN => n37060);
   U29286 : OAI222_X1 port map( A1 => n30983, A2 => n39120, B1 => n31047, B2 =>
                           n39114, C1 => n30919, C2 => n39108, ZN => n37063);
   U29287 : AOI221_X1 port map( B1 => n39132, B2 => n32816, C1 => n39126, C2 =>
                           n32768, A => n37044, ZN => n37041);
   U29288 : OAI222_X1 port map( A1 => n30982, A2 => n39120, B1 => n31046, B2 =>
                           n39114, C1 => n30918, C2 => n39108, ZN => n37044);
   U29289 : AOI221_X1 port map( B1 => n39136, B2 => n32844, C1 => n39130, C2 =>
                           n32832, A => n36208, ZN => n36205);
   U29290 : OAI222_X1 port map( A1 => n30938, A2 => n39124, B1 => n31002, B2 =>
                           n39118, C1 => n30874, C2 => n39112, ZN => n36208);
   U29291 : AOI221_X1 port map( B1 => n39136, B2 => n32843, C1 => n39130, C2 =>
                           n32831, A => n36189, ZN => n36186);
   U29292 : OAI222_X1 port map( A1 => n30937, A2 => n39124, B1 => n31001, B2 =>
                           n39118, C1 => n30873, C2 => n39112, ZN => n36189);
   U29293 : AOI221_X1 port map( B1 => n39136, B2 => n32842, C1 => n39130, C2 =>
                           n32830, A => n36170, ZN => n36167);
   U29294 : OAI222_X1 port map( A1 => n30936, A2 => n39124, B1 => n31000, B2 =>
                           n39118, C1 => n30872, C2 => n39112, ZN => n36170);
   U29295 : AOI221_X1 port map( B1 => n39136, B2 => n32841, C1 => n39130, C2 =>
                           n32829, A => n36151, ZN => n36148);
   U29296 : OAI222_X1 port map( A1 => n30935, A2 => n39124, B1 => n30999, B2 =>
                           n39118, C1 => n30871, C2 => n39112, ZN => n36151);
   U29297 : AOI221_X1 port map( B1 => n39136, B2 => n32840, C1 => n39130, C2 =>
                           n32828, A => n36132, ZN => n36129);
   U29298 : OAI222_X1 port map( A1 => n30934, A2 => n39124, B1 => n30998, B2 =>
                           n39118, C1 => n30870, C2 => n39112, ZN => n36132);
   U29299 : AOI221_X1 port map( B1 => n39136, B2 => n32839, C1 => n39130, C2 =>
                           n32827, A => n36113, ZN => n36110);
   U29300 : OAI222_X1 port map( A1 => n30933, A2 => n39124, B1 => n30997, B2 =>
                           n39118, C1 => n30869, C2 => n39112, ZN => n36113);
   U29301 : AOI221_X1 port map( B1 => n39639, B2 => n32475, C1 => n39633, C2 =>
                           n32471, A => n33469, ZN => n33459);
   U29302 : OAI222_X1 port map( A1 => n30992, A2 => n39627, B1 => n31056, B2 =>
                           n39621, C1 => n30928, C2 => n39615, ZN => n33469);
   U29303 : AOI221_X1 port map( B1 => n39387, B2 => n32475, C1 => n39381, C2 =>
                           n32471, A => n34743, ZN => n34733);
   U29304 : OAI222_X1 port map( A1 => n30992, A2 => n39375, B1 => n31056, B2 =>
                           n39369, C1 => n30928, C2 => n39363, ZN => n34743);
   U29305 : AOI221_X1 port map( B1 => n39639, B2 => n32474, C1 => n39633, C2 =>
                           n32470, A => n33501, ZN => n33498);
   U29306 : OAI222_X1 port map( A1 => n30991, A2 => n39627, B1 => n31055, B2 =>
                           n39621, C1 => n30927, C2 => n39615, ZN => n33501);
   U29307 : AOI221_X1 port map( B1 => n39387, B2 => n32474, C1 => n39381, C2 =>
                           n32470, A => n34775, ZN => n34772);
   U29308 : OAI222_X1 port map( A1 => n30991, A2 => n39375, B1 => n31055, B2 =>
                           n39369, C1 => n30927, C2 => n39363, ZN => n34775);
   U29309 : AOI221_X1 port map( B1 => n39639, B2 => n32473, C1 => n39633, C2 =>
                           n32469, A => n33520, ZN => n33517);
   U29310 : OAI222_X1 port map( A1 => n30990, A2 => n39627, B1 => n31054, B2 =>
                           n39621, C1 => n30926, C2 => n39615, ZN => n33520);
   U29311 : AOI221_X1 port map( B1 => n39387, B2 => n32473, C1 => n39381, C2 =>
                           n32469, A => n34794, ZN => n34791);
   U29312 : OAI222_X1 port map( A1 => n30990, A2 => n39375, B1 => n31054, B2 =>
                           n39369, C1 => n30926, C2 => n39363, ZN => n34794);
   U29313 : AOI221_X1 port map( B1 => n39639, B2 => n32472, C1 => n39633, C2 =>
                           n32468, A => n33539, ZN => n33536);
   U29314 : OAI222_X1 port map( A1 => n30989, A2 => n39627, B1 => n31053, B2 =>
                           n39621, C1 => n30925, C2 => n39615, ZN => n33539);
   U29315 : AOI221_X1 port map( B1 => n39387, B2 => n32472, C1 => n39381, C2 =>
                           n32468, A => n34813, ZN => n34810);
   U29316 : OAI222_X1 port map( A1 => n30989, A2 => n39375, B1 => n31053, B2 =>
                           n39369, C1 => n30925, C2 => n39363, ZN => n34813);
   U29317 : OAI222_X1 port map( A1 => n40593, A2 => n40745, B1 => n40586, B2 =>
                           n41129, C1 => n40577, C2 => n32321, ZN => n9866);
   U29318 : OAI222_X1 port map( A1 => n40593, A2 => n40751, B1 => n40586, B2 =>
                           n41135, C1 => n40578, C2 => n32320, ZN => n9865);
   U29319 : OAI222_X1 port map( A1 => n40593, A2 => n40757, B1 => n40586, B2 =>
                           n41141, C1 => n40578, C2 => n32319, ZN => n9864);
   U29320 : OAI222_X1 port map( A1 => n40593, A2 => n40763, B1 => n40586, B2 =>
                           n41147, C1 => n40578, C2 => n32318, ZN => n9863);
   U29321 : OAI222_X1 port map( A1 => n40592, A2 => n40769, B1 => n40585, B2 =>
                           n41153, C1 => n40578, C2 => n32317, ZN => n9862);
   U29322 : OAI222_X1 port map( A1 => n40592, A2 => n40775, B1 => n40585, B2 =>
                           n41159, C1 => n40578, C2 => n32316, ZN => n9861);
   U29323 : OAI222_X1 port map( A1 => n40592, A2 => n40781, B1 => n40585, B2 =>
                           n41165, C1 => n40578, C2 => n32315, ZN => n9860);
   U29324 : OAI222_X1 port map( A1 => n40592, A2 => n40787, B1 => n40585, B2 =>
                           n41171, C1 => n40578, C2 => n32314, ZN => n9859);
   U29325 : OAI222_X1 port map( A1 => n40592, A2 => n40793, B1 => n40585, B2 =>
                           n41177, C1 => n40578, C2 => n32313, ZN => n9858);
   U29326 : OAI222_X1 port map( A1 => n40592, A2 => n40799, B1 => n40585, B2 =>
                           n41183, C1 => n40578, C2 => n32312, ZN => n9857);
   U29327 : OAI222_X1 port map( A1 => n40592, A2 => n40805, B1 => n40585, B2 =>
                           n41189, C1 => n40578, C2 => n32311, ZN => n9856);
   U29328 : OAI222_X1 port map( A1 => n40592, A2 => n40811, B1 => n40585, B2 =>
                           n41195, C1 => n40578, C2 => n32310, ZN => n9855);
   U29329 : OAI222_X1 port map( A1 => n40592, A2 => n40817, B1 => n40585, B2 =>
                           n41201, C1 => n40579, C2 => n32309, ZN => n9854);
   U29330 : OAI222_X1 port map( A1 => n40592, A2 => n40823, B1 => n40585, B2 =>
                           n41207, C1 => n40579, C2 => n32308, ZN => n9853);
   U29331 : OAI222_X1 port map( A1 => n40592, A2 => n40829, B1 => n40585, B2 =>
                           n41213, C1 => n40579, C2 => n32307, ZN => n9852);
   U29332 : OAI222_X1 port map( A1 => n40592, A2 => n40835, B1 => n40585, B2 =>
                           n41219, C1 => n40579, C2 => n32306, ZN => n9851);
   U29333 : OAI222_X1 port map( A1 => n40591, A2 => n40841, B1 => n40584, B2 =>
                           n41225, C1 => n40579, C2 => n32305, ZN => n9850);
   U29334 : OAI222_X1 port map( A1 => n40591, A2 => n40847, B1 => n40584, B2 =>
                           n41231, C1 => n40579, C2 => n32304, ZN => n9849);
   U29335 : OAI222_X1 port map( A1 => n40591, A2 => n40853, B1 => n40584, B2 =>
                           n41237, C1 => n40579, C2 => n32303, ZN => n9848);
   U29336 : OAI222_X1 port map( A1 => n40591, A2 => n40859, B1 => n40584, B2 =>
                           n41243, C1 => n40579, C2 => n32302, ZN => n9847);
   U29337 : OAI222_X1 port map( A1 => n40591, A2 => n40865, B1 => n40584, B2 =>
                           n41249, C1 => n40579, C2 => n32301, ZN => n9846);
   U29338 : OAI222_X1 port map( A1 => n40591, A2 => n40871, B1 => n40584, B2 =>
                           n41255, C1 => n40579, C2 => n32300, ZN => n9845);
   U29339 : OAI222_X1 port map( A1 => n40591, A2 => n40877, B1 => n40584, B2 =>
                           n41261, C1 => n40579, C2 => n32299, ZN => n9844);
   U29340 : OAI222_X1 port map( A1 => n40591, A2 => n40883, B1 => n40584, B2 =>
                           n41267, C1 => n40579, C2 => n32298, ZN => n9843);
   U29341 : OAI222_X1 port map( A1 => n40591, A2 => n40889, B1 => n40584, B2 =>
                           n41273, C1 => n40580, C2 => n32297, ZN => n9842);
   U29342 : OAI222_X1 port map( A1 => n40591, A2 => n40895, B1 => n40584, B2 =>
                           n41279, C1 => n40580, C2 => n32296, ZN => n9841);
   U29343 : OAI222_X1 port map( A1 => n40591, A2 => n40901, B1 => n40584, B2 =>
                           n41285, C1 => n40580, C2 => n32295, ZN => n9840);
   U29344 : OAI222_X1 port map( A1 => n40591, A2 => n40907, B1 => n40584, B2 =>
                           n41291, C1 => n40580, C2 => n32294, ZN => n9839);
   U29345 : OAI222_X1 port map( A1 => n40590, A2 => n40913, B1 => n40583, B2 =>
                           n41297, C1 => n40580, C2 => n32293, ZN => n9838);
   U29346 : OAI222_X1 port map( A1 => n40590, A2 => n40919, B1 => n40583, B2 =>
                           n41303, C1 => n40580, C2 => n32292, ZN => n9837);
   U29347 : OAI222_X1 port map( A1 => n40590, A2 => n40925, B1 => n40583, B2 =>
                           n41309, C1 => n40580, C2 => n32291, ZN => n9836);
   U29348 : OAI222_X1 port map( A1 => n40590, A2 => n40931, B1 => n40583, B2 =>
                           n41315, C1 => n40580, C2 => n32290, ZN => n9835);
   U29349 : OAI222_X1 port map( A1 => n40590, A2 => n40937, B1 => n40583, B2 =>
                           n41321, C1 => n40580, C2 => n32289, ZN => n9834);
   U29350 : OAI222_X1 port map( A1 => n40590, A2 => n40943, B1 => n40583, B2 =>
                           n41327, C1 => n40580, C2 => n32288, ZN => n9833);
   U29351 : OAI222_X1 port map( A1 => n40590, A2 => n40949, B1 => n40583, B2 =>
                           n41333, C1 => n40580, C2 => n32287, ZN => n9832);
   U29352 : OAI222_X1 port map( A1 => n40590, A2 => n40961, B1 => n40583, B2 =>
                           n41345, C1 => n40580, C2 => n32286, ZN => n9830);
   U29353 : OAI222_X1 port map( A1 => n40601, A2 => n40555, B1 => n40985, B2 =>
                           n40548, C1 => n40536, C2 => n32285, ZN => n9762);
   U29354 : OAI222_X1 port map( A1 => n40607, A2 => n40555, B1 => n40991, B2 =>
                           n40548, C1 => n40536, C2 => n32284, ZN => n9761);
   U29355 : OAI222_X1 port map( A1 => n40613, A2 => n40555, B1 => n40997, B2 =>
                           n40548, C1 => n40536, C2 => n32283, ZN => n9760);
   U29356 : OAI222_X1 port map( A1 => n40619, A2 => n40555, B1 => n41003, B2 =>
                           n40548, C1 => n40536, C2 => n32282, ZN => n9759);
   U29357 : OAI222_X1 port map( A1 => n40601, A2 => n40575, B1 => n40985, B2 =>
                           n40568, C1 => n40556, C2 => n32281, ZN => n9826);
   U29358 : OAI222_X1 port map( A1 => n40607, A2 => n40575, B1 => n40991, B2 =>
                           n40568, C1 => n40556, C2 => n32280, ZN => n9825);
   U29359 : OAI222_X1 port map( A1 => n40613, A2 => n40575, B1 => n40997, B2 =>
                           n40568, C1 => n40556, C2 => n32279, ZN => n9824);
   U29360 : OAI222_X1 port map( A1 => n40619, A2 => n40575, B1 => n41003, B2 =>
                           n40568, C1 => n40556, C2 => n32278, ZN => n9823);
   U29361 : OAI222_X1 port map( A1 => n40600, A2 => n40455, B1 => n40984, B2 =>
                           n40448, C1 => n40436, C2 => n32277, ZN => n9442);
   U29362 : OAI222_X1 port map( A1 => n40606, A2 => n40455, B1 => n40990, B2 =>
                           n40448, C1 => n40436, C2 => n32276, ZN => n9441);
   U29363 : OAI222_X1 port map( A1 => n40612, A2 => n40455, B1 => n40996, B2 =>
                           n40448, C1 => n40436, C2 => n32275, ZN => n9440);
   U29364 : OAI222_X1 port map( A1 => n40618, A2 => n40455, B1 => n41002, B2 =>
                           n40448, C1 => n40436, C2 => n32274, ZN => n9439);
   U29365 : OAI222_X1 port map( A1 => n40600, A2 => n40495, B1 => n40984, B2 =>
                           n40488, C1 => n40476, C2 => n32273, ZN => n9570);
   U29366 : OAI222_X1 port map( A1 => n40606, A2 => n40495, B1 => n40990, B2 =>
                           n40488, C1 => n40476, C2 => n32272, ZN => n9569);
   U29367 : OAI222_X1 port map( A1 => n40612, A2 => n40495, B1 => n40996, B2 =>
                           n40488, C1 => n40476, C2 => n32271, ZN => n9568);
   U29368 : OAI222_X1 port map( A1 => n40618, A2 => n40495, B1 => n41002, B2 =>
                           n40488, C1 => n40476, C2 => n32270, ZN => n9567);
   U29369 : OAI222_X1 port map( A1 => n40600, A2 => n40475, B1 => n40984, B2 =>
                           n40468, C1 => n40456, C2 => n32269, ZN => n9506);
   U29370 : OAI222_X1 port map( A1 => n40606, A2 => n40475, B1 => n40990, B2 =>
                           n40468, C1 => n40456, C2 => n32268, ZN => n9505);
   U29371 : OAI222_X1 port map( A1 => n40612, A2 => n40475, B1 => n40996, B2 =>
                           n40468, C1 => n40456, C2 => n32267, ZN => n9504);
   U29372 : OAI222_X1 port map( A1 => n40618, A2 => n40475, B1 => n41002, B2 =>
                           n40468, C1 => n40456, C2 => n32266, ZN => n9503);
   U29373 : OAI222_X1 port map( A1 => n40595, A2 => n40601, B1 => n40588, B2 =>
                           n40985, C1 => n40576, C2 => n32265, ZN => n9890);
   U29374 : OAI222_X1 port map( A1 => n40595, A2 => n40607, B1 => n40588, B2 =>
                           n40991, C1 => n40576, C2 => n32264, ZN => n9889);
   U29375 : OAI222_X1 port map( A1 => n40595, A2 => n40613, B1 => n40588, B2 =>
                           n40997, C1 => n40576, C2 => n32263, ZN => n9888);
   U29376 : OAI222_X1 port map( A1 => n40595, A2 => n40619, B1 => n40588, B2 =>
                           n41003, C1 => n40576, C2 => n32262, ZN => n9887);
   U29377 : OAI222_X1 port map( A1 => n40594, A2 => n40625, B1 => n40587, B2 =>
                           n41009, C1 => n40576, C2 => n32074, ZN => n9886);
   U29378 : OAI222_X1 port map( A1 => n40594, A2 => n40631, B1 => n40587, B2 =>
                           n41015, C1 => n40576, C2 => n32073, ZN => n9885);
   U29379 : OAI222_X1 port map( A1 => n40594, A2 => n40637, B1 => n40587, B2 =>
                           n41021, C1 => n40576, C2 => n32072, ZN => n9884);
   U29380 : OAI222_X1 port map( A1 => n40594, A2 => n40643, B1 => n40587, B2 =>
                           n41027, C1 => n40576, C2 => n32071, ZN => n9883);
   U29381 : OAI222_X1 port map( A1 => n40594, A2 => n40649, B1 => n40587, B2 =>
                           n41033, C1 => n40576, C2 => n32070, ZN => n9882);
   U29382 : OAI222_X1 port map( A1 => n40594, A2 => n40655, B1 => n40587, B2 =>
                           n41039, C1 => n40576, C2 => n32069, ZN => n9881);
   U29383 : OAI222_X1 port map( A1 => n40594, A2 => n40661, B1 => n40587, B2 =>
                           n41045, C1 => n40576, C2 => n32068, ZN => n9880);
   U29384 : OAI222_X1 port map( A1 => n40594, A2 => n40667, B1 => n40587, B2 =>
                           n41051, C1 => n40576, C2 => n32067, ZN => n9879);
   U29385 : OAI222_X1 port map( A1 => n40594, A2 => n40673, B1 => n40587, B2 =>
                           n41057, C1 => n40577, C2 => n32066, ZN => n9878);
   U29386 : OAI222_X1 port map( A1 => n40594, A2 => n40679, B1 => n40587, B2 =>
                           n41063, C1 => n40577, C2 => n32065, ZN => n9877);
   U29387 : OAI222_X1 port map( A1 => n40594, A2 => n40685, B1 => n40587, B2 =>
                           n41069, C1 => n40577, C2 => n32064, ZN => n9876);
   U29388 : OAI222_X1 port map( A1 => n40594, A2 => n40691, B1 => n40587, B2 =>
                           n41075, C1 => n40578, C2 => n32063, ZN => n9875);
   U29389 : OAI222_X1 port map( A1 => n40593, A2 => n40697, B1 => n40586, B2 =>
                           n41081, C1 => n40577, C2 => n32062, ZN => n9874);
   U29390 : OAI222_X1 port map( A1 => n40593, A2 => n40703, B1 => n40586, B2 =>
                           n41087, C1 => n40577, C2 => n32061, ZN => n9873);
   U29391 : OAI222_X1 port map( A1 => n40593, A2 => n40709, B1 => n40586, B2 =>
                           n41093, C1 => n40577, C2 => n32060, ZN => n9872);
   U29392 : OAI222_X1 port map( A1 => n40593, A2 => n40715, B1 => n40586, B2 =>
                           n41099, C1 => n40577, C2 => n32059, ZN => n9871);
   U29393 : OAI222_X1 port map( A1 => n40593, A2 => n40721, B1 => n40586, B2 =>
                           n41105, C1 => n40577, C2 => n32058, ZN => n9870);
   U29394 : OAI222_X1 port map( A1 => n40593, A2 => n40727, B1 => n40586, B2 =>
                           n41111, C1 => n40577, C2 => n32057, ZN => n9869);
   U29395 : OAI222_X1 port map( A1 => n40593, A2 => n40733, B1 => n40586, B2 =>
                           n41117, C1 => n40577, C2 => n32056, ZN => n9868);
   U29396 : OAI222_X1 port map( A1 => n40593, A2 => n40739, B1 => n40586, B2 =>
                           n41123, C1 => n40577, C2 => n32055, ZN => n9867);
   U29397 : OAI222_X1 port map( A1 => n40625, A2 => n40574, B1 => n41009, B2 =>
                           n40567, C1 => n40556, C2 => n32050, ZN => n9822);
   U29398 : OAI222_X1 port map( A1 => n40631, A2 => n40574, B1 => n41015, B2 =>
                           n40567, C1 => n40556, C2 => n32049, ZN => n9821);
   U29399 : OAI222_X1 port map( A1 => n40637, A2 => n40574, B1 => n41021, B2 =>
                           n40567, C1 => n40556, C2 => n32048, ZN => n9820);
   U29400 : OAI222_X1 port map( A1 => n40643, A2 => n40574, B1 => n41027, B2 =>
                           n40567, C1 => n40556, C2 => n32047, ZN => n9819);
   U29401 : OAI222_X1 port map( A1 => n40649, A2 => n40574, B1 => n41033, B2 =>
                           n40567, C1 => n40556, C2 => n32046, ZN => n9818);
   U29402 : OAI222_X1 port map( A1 => n40655, A2 => n40574, B1 => n41039, B2 =>
                           n40567, C1 => n40556, C2 => n32045, ZN => n9817);
   U29403 : OAI222_X1 port map( A1 => n40661, A2 => n40574, B1 => n41045, B2 =>
                           n40567, C1 => n40556, C2 => n32044, ZN => n9816);
   U29404 : OAI222_X1 port map( A1 => n40667, A2 => n40574, B1 => n41051, B2 =>
                           n40567, C1 => n40556, C2 => n32043, ZN => n9815);
   U29405 : OAI222_X1 port map( A1 => n40673, A2 => n40574, B1 => n41057, B2 =>
                           n40567, C1 => n40557, C2 => n32042, ZN => n9814);
   U29406 : OAI222_X1 port map( A1 => n40679, A2 => n40574, B1 => n41063, B2 =>
                           n40567, C1 => n40557, C2 => n32041, ZN => n9813);
   U29407 : OAI222_X1 port map( A1 => n40685, A2 => n40574, B1 => n41069, B2 =>
                           n40567, C1 => n40557, C2 => n32040, ZN => n9812);
   U29408 : OAI222_X1 port map( A1 => n40691, A2 => n40574, B1 => n41075, B2 =>
                           n40567, C1 => n40558, C2 => n32039, ZN => n9811);
   U29409 : OAI222_X1 port map( A1 => n40697, A2 => n40573, B1 => n41081, B2 =>
                           n40566, C1 => n40557, C2 => n32038, ZN => n9810);
   U29410 : OAI222_X1 port map( A1 => n40703, A2 => n40573, B1 => n41087, B2 =>
                           n40566, C1 => n40557, C2 => n32037, ZN => n9809);
   U29411 : OAI222_X1 port map( A1 => n40709, A2 => n40573, B1 => n41093, B2 =>
                           n40566, C1 => n40557, C2 => n32036, ZN => n9808);
   U29412 : OAI222_X1 port map( A1 => n40715, A2 => n40573, B1 => n41099, B2 =>
                           n40566, C1 => n40557, C2 => n32035, ZN => n9807);
   U29413 : OAI222_X1 port map( A1 => n40721, A2 => n40573, B1 => n41105, B2 =>
                           n40566, C1 => n40557, C2 => n32034, ZN => n9806);
   U29414 : OAI222_X1 port map( A1 => n40727, A2 => n40573, B1 => n41111, B2 =>
                           n40566, C1 => n40557, C2 => n32033, ZN => n9805);
   U29415 : OAI222_X1 port map( A1 => n40733, A2 => n40573, B1 => n41117, B2 =>
                           n40566, C1 => n40557, C2 => n32032, ZN => n9804);
   U29416 : OAI222_X1 port map( A1 => n40739, A2 => n40573, B1 => n41123, B2 =>
                           n40566, C1 => n40557, C2 => n32031, ZN => n9803);
   U29417 : OAI222_X1 port map( A1 => n40745, A2 => n40573, B1 => n41129, B2 =>
                           n40566, C1 => n40557, C2 => n32030, ZN => n9802);
   U29418 : OAI222_X1 port map( A1 => n40751, A2 => n40573, B1 => n41135, B2 =>
                           n40566, C1 => n40558, C2 => n32029, ZN => n9801);
   U29419 : OAI222_X1 port map( A1 => n40757, A2 => n40573, B1 => n41141, B2 =>
                           n40566, C1 => n40558, C2 => n32028, ZN => n9800);
   U29420 : OAI222_X1 port map( A1 => n40763, A2 => n40573, B1 => n41147, B2 =>
                           n40566, C1 => n40558, C2 => n32027, ZN => n9799);
   U29421 : OAI222_X1 port map( A1 => n40769, A2 => n40572, B1 => n41153, B2 =>
                           n40565, C1 => n40558, C2 => n32026, ZN => n9798);
   U29422 : OAI222_X1 port map( A1 => n40775, A2 => n40572, B1 => n41159, B2 =>
                           n40565, C1 => n40558, C2 => n32025, ZN => n9797);
   U29423 : OAI222_X1 port map( A1 => n40781, A2 => n40572, B1 => n41165, B2 =>
                           n40565, C1 => n40558, C2 => n32024, ZN => n9796);
   U29424 : OAI222_X1 port map( A1 => n40787, A2 => n40572, B1 => n41171, B2 =>
                           n40565, C1 => n40558, C2 => n32023, ZN => n9795);
   U29425 : OAI222_X1 port map( A1 => n40793, A2 => n40572, B1 => n41177, B2 =>
                           n40565, C1 => n40558, C2 => n32022, ZN => n9794);
   U29426 : OAI222_X1 port map( A1 => n40799, A2 => n40572, B1 => n41183, B2 =>
                           n40565, C1 => n40558, C2 => n32021, ZN => n9793);
   U29427 : OAI222_X1 port map( A1 => n40805, A2 => n40572, B1 => n41189, B2 =>
                           n40565, C1 => n40558, C2 => n32020, ZN => n9792);
   U29428 : OAI222_X1 port map( A1 => n40811, A2 => n40572, B1 => n41195, B2 =>
                           n40565, C1 => n40558, C2 => n32019, ZN => n9791);
   U29429 : OAI222_X1 port map( A1 => n40817, A2 => n40572, B1 => n41201, B2 =>
                           n40565, C1 => n40559, C2 => n32018, ZN => n9790);
   U29430 : OAI222_X1 port map( A1 => n40823, A2 => n40572, B1 => n41207, B2 =>
                           n40565, C1 => n40559, C2 => n32017, ZN => n9789);
   U29431 : OAI222_X1 port map( A1 => n40829, A2 => n40572, B1 => n41213, B2 =>
                           n40565, C1 => n40559, C2 => n32016, ZN => n9788);
   U29432 : OAI222_X1 port map( A1 => n40835, A2 => n40572, B1 => n41219, B2 =>
                           n40565, C1 => n40559, C2 => n32015, ZN => n9787);
   U29433 : OAI222_X1 port map( A1 => n40841, A2 => n40571, B1 => n41225, B2 =>
                           n40564, C1 => n40559, C2 => n32014, ZN => n9786);
   U29434 : OAI222_X1 port map( A1 => n40847, A2 => n40571, B1 => n41231, B2 =>
                           n40564, C1 => n40559, C2 => n32013, ZN => n9785);
   U29435 : OAI222_X1 port map( A1 => n40853, A2 => n40571, B1 => n41237, B2 =>
                           n40564, C1 => n40559, C2 => n32012, ZN => n9784);
   U29436 : OAI222_X1 port map( A1 => n40859, A2 => n40571, B1 => n41243, B2 =>
                           n40564, C1 => n40559, C2 => n32011, ZN => n9783);
   U29437 : OAI222_X1 port map( A1 => n40865, A2 => n40571, B1 => n41249, B2 =>
                           n40564, C1 => n40559, C2 => n32010, ZN => n9782);
   U29438 : OAI222_X1 port map( A1 => n40871, A2 => n40571, B1 => n41255, B2 =>
                           n40564, C1 => n40559, C2 => n32009, ZN => n9781);
   U29439 : OAI222_X1 port map( A1 => n40877, A2 => n40571, B1 => n41261, B2 =>
                           n40564, C1 => n40559, C2 => n32008, ZN => n9780);
   U29440 : OAI222_X1 port map( A1 => n40883, A2 => n40571, B1 => n41267, B2 =>
                           n40564, C1 => n40559, C2 => n32007, ZN => n9779);
   U29441 : OAI222_X1 port map( A1 => n40889, A2 => n40571, B1 => n41273, B2 =>
                           n40564, C1 => n40560, C2 => n32006, ZN => n9778);
   U29442 : OAI222_X1 port map( A1 => n40895, A2 => n40571, B1 => n41279, B2 =>
                           n40564, C1 => n40560, C2 => n32005, ZN => n9777);
   U29443 : OAI222_X1 port map( A1 => n40901, A2 => n40571, B1 => n41285, B2 =>
                           n40564, C1 => n40560, C2 => n32004, ZN => n9776);
   U29444 : OAI222_X1 port map( A1 => n40907, A2 => n40571, B1 => n41291, B2 =>
                           n40564, C1 => n40560, C2 => n32003, ZN => n9775);
   U29445 : OAI222_X1 port map( A1 => n40913, A2 => n40570, B1 => n41297, B2 =>
                           n40563, C1 => n40560, C2 => n32002, ZN => n9774);
   U29446 : OAI222_X1 port map( A1 => n40919, A2 => n40570, B1 => n41303, B2 =>
                           n40563, C1 => n40560, C2 => n32001, ZN => n9773);
   U29447 : OAI222_X1 port map( A1 => n40925, A2 => n40570, B1 => n41309, B2 =>
                           n40563, C1 => n40560, C2 => n32000, ZN => n9772);
   U29448 : OAI222_X1 port map( A1 => n40931, A2 => n40570, B1 => n41315, B2 =>
                           n40563, C1 => n40560, C2 => n31999, ZN => n9771);
   U29449 : OAI222_X1 port map( A1 => n40937, A2 => n40570, B1 => n41321, B2 =>
                           n40563, C1 => n40560, C2 => n31998, ZN => n9770);
   U29450 : OAI222_X1 port map( A1 => n40943, A2 => n40570, B1 => n41327, B2 =>
                           n40563, C1 => n40560, C2 => n31997, ZN => n9769);
   U29451 : OAI222_X1 port map( A1 => n40949, A2 => n40570, B1 => n41333, B2 =>
                           n40563, C1 => n40560, C2 => n31996, ZN => n9768);
   U29452 : OAI222_X1 port map( A1 => n40961, A2 => n40570, B1 => n41345, B2 =>
                           n40563, C1 => n40560, C2 => n31994, ZN => n9766);
   U29453 : OAI222_X1 port map( A1 => n40625, A2 => n40554, B1 => n41009, B2 =>
                           n40547, C1 => n40536, C2 => n31990, ZN => n9758);
   U29454 : OAI222_X1 port map( A1 => n40631, A2 => n40554, B1 => n41015, B2 =>
                           n40547, C1 => n40536, C2 => n31989, ZN => n9757);
   U29455 : OAI222_X1 port map( A1 => n40637, A2 => n40554, B1 => n41021, B2 =>
                           n40547, C1 => n40536, C2 => n31988, ZN => n9756);
   U29456 : OAI222_X1 port map( A1 => n40643, A2 => n40554, B1 => n41027, B2 =>
                           n40547, C1 => n40536, C2 => n31987, ZN => n9755);
   U29457 : OAI222_X1 port map( A1 => n40649, A2 => n40554, B1 => n41033, B2 =>
                           n40547, C1 => n40536, C2 => n31986, ZN => n9754);
   U29458 : OAI222_X1 port map( A1 => n40655, A2 => n40554, B1 => n41039, B2 =>
                           n40547, C1 => n40536, C2 => n31985, ZN => n9753);
   U29459 : OAI222_X1 port map( A1 => n40661, A2 => n40554, B1 => n41045, B2 =>
                           n40547, C1 => n40536, C2 => n31984, ZN => n9752);
   U29460 : OAI222_X1 port map( A1 => n40667, A2 => n40554, B1 => n41051, B2 =>
                           n40547, C1 => n40536, C2 => n31983, ZN => n9751);
   U29461 : OAI222_X1 port map( A1 => n40673, A2 => n40554, B1 => n41057, B2 =>
                           n40547, C1 => n40537, C2 => n31982, ZN => n9750);
   U29462 : OAI222_X1 port map( A1 => n40679, A2 => n40554, B1 => n41063, B2 =>
                           n40547, C1 => n40537, C2 => n31981, ZN => n9749);
   U29463 : OAI222_X1 port map( A1 => n40685, A2 => n40554, B1 => n41069, B2 =>
                           n40547, C1 => n40537, C2 => n31980, ZN => n9748);
   U29464 : OAI222_X1 port map( A1 => n40691, A2 => n40554, B1 => n41075, B2 =>
                           n40547, C1 => n40538, C2 => n31979, ZN => n9747);
   U29465 : OAI222_X1 port map( A1 => n40697, A2 => n40553, B1 => n41081, B2 =>
                           n40546, C1 => n40537, C2 => n31978, ZN => n9746);
   U29466 : OAI222_X1 port map( A1 => n40703, A2 => n40553, B1 => n41087, B2 =>
                           n40546, C1 => n40537, C2 => n31977, ZN => n9745);
   U29467 : OAI222_X1 port map( A1 => n40709, A2 => n40553, B1 => n41093, B2 =>
                           n40546, C1 => n40537, C2 => n31976, ZN => n9744);
   U29468 : OAI222_X1 port map( A1 => n40715, A2 => n40553, B1 => n41099, B2 =>
                           n40546, C1 => n40537, C2 => n31975, ZN => n9743);
   U29469 : OAI222_X1 port map( A1 => n40721, A2 => n40553, B1 => n41105, B2 =>
                           n40546, C1 => n40537, C2 => n31974, ZN => n9742);
   U29470 : OAI222_X1 port map( A1 => n40727, A2 => n40553, B1 => n41111, B2 =>
                           n40546, C1 => n40537, C2 => n31973, ZN => n9741);
   U29471 : OAI222_X1 port map( A1 => n40733, A2 => n40553, B1 => n41117, B2 =>
                           n40546, C1 => n40537, C2 => n31972, ZN => n9740);
   U29472 : OAI222_X1 port map( A1 => n40739, A2 => n40553, B1 => n41123, B2 =>
                           n40546, C1 => n40537, C2 => n31971, ZN => n9739);
   U29473 : OAI222_X1 port map( A1 => n40745, A2 => n40553, B1 => n41129, B2 =>
                           n40546, C1 => n40537, C2 => n31970, ZN => n9738);
   U29474 : OAI222_X1 port map( A1 => n40751, A2 => n40553, B1 => n41135, B2 =>
                           n40546, C1 => n40538, C2 => n31969, ZN => n9737);
   U29475 : OAI222_X1 port map( A1 => n40757, A2 => n40553, B1 => n41141, B2 =>
                           n40546, C1 => n40538, C2 => n31968, ZN => n9736);
   U29476 : OAI222_X1 port map( A1 => n40763, A2 => n40553, B1 => n41147, B2 =>
                           n40546, C1 => n40538, C2 => n31967, ZN => n9735);
   U29477 : OAI222_X1 port map( A1 => n40769, A2 => n40552, B1 => n41153, B2 =>
                           n40545, C1 => n40538, C2 => n31966, ZN => n9734);
   U29478 : OAI222_X1 port map( A1 => n40775, A2 => n40552, B1 => n41159, B2 =>
                           n40545, C1 => n40538, C2 => n31965, ZN => n9733);
   U29479 : OAI222_X1 port map( A1 => n40781, A2 => n40552, B1 => n41165, B2 =>
                           n40545, C1 => n40538, C2 => n31964, ZN => n9732);
   U29480 : OAI222_X1 port map( A1 => n40787, A2 => n40552, B1 => n41171, B2 =>
                           n40545, C1 => n40538, C2 => n31963, ZN => n9731);
   U29481 : OAI222_X1 port map( A1 => n40793, A2 => n40552, B1 => n41177, B2 =>
                           n40545, C1 => n40538, C2 => n31962, ZN => n9730);
   U29482 : OAI222_X1 port map( A1 => n40799, A2 => n40552, B1 => n41183, B2 =>
                           n40545, C1 => n40538, C2 => n31961, ZN => n9729);
   U29483 : OAI222_X1 port map( A1 => n40805, A2 => n40552, B1 => n41189, B2 =>
                           n40545, C1 => n40538, C2 => n31960, ZN => n9728);
   U29484 : OAI222_X1 port map( A1 => n40811, A2 => n40552, B1 => n41195, B2 =>
                           n40545, C1 => n40538, C2 => n31959, ZN => n9727);
   U29485 : OAI222_X1 port map( A1 => n40817, A2 => n40552, B1 => n41201, B2 =>
                           n40545, C1 => n40539, C2 => n31958, ZN => n9726);
   U29486 : OAI222_X1 port map( A1 => n40823, A2 => n40552, B1 => n41207, B2 =>
                           n40545, C1 => n40539, C2 => n31957, ZN => n9725);
   U29487 : OAI222_X1 port map( A1 => n40829, A2 => n40552, B1 => n41213, B2 =>
                           n40545, C1 => n40539, C2 => n31956, ZN => n9724);
   U29488 : OAI222_X1 port map( A1 => n40835, A2 => n40552, B1 => n41219, B2 =>
                           n40545, C1 => n40539, C2 => n31955, ZN => n9723);
   U29489 : OAI222_X1 port map( A1 => n40841, A2 => n40551, B1 => n41225, B2 =>
                           n40544, C1 => n40539, C2 => n31954, ZN => n9722);
   U29490 : OAI222_X1 port map( A1 => n40847, A2 => n40551, B1 => n41231, B2 =>
                           n40544, C1 => n40539, C2 => n31953, ZN => n9721);
   U29491 : OAI222_X1 port map( A1 => n40853, A2 => n40551, B1 => n41237, B2 =>
                           n40544, C1 => n40539, C2 => n31952, ZN => n9720);
   U29492 : OAI222_X1 port map( A1 => n40859, A2 => n40551, B1 => n41243, B2 =>
                           n40544, C1 => n40539, C2 => n31951, ZN => n9719);
   U29493 : OAI222_X1 port map( A1 => n40865, A2 => n40551, B1 => n41249, B2 =>
                           n40544, C1 => n40539, C2 => n31950, ZN => n9718);
   U29494 : OAI222_X1 port map( A1 => n40871, A2 => n40551, B1 => n41255, B2 =>
                           n40544, C1 => n40539, C2 => n31949, ZN => n9717);
   U29495 : OAI222_X1 port map( A1 => n40877, A2 => n40551, B1 => n41261, B2 =>
                           n40544, C1 => n40539, C2 => n31948, ZN => n9716);
   U29496 : OAI222_X1 port map( A1 => n40883, A2 => n40551, B1 => n41267, B2 =>
                           n40544, C1 => n40539, C2 => n31947, ZN => n9715);
   U29497 : OAI222_X1 port map( A1 => n40889, A2 => n40551, B1 => n41273, B2 =>
                           n40544, C1 => n40540, C2 => n31946, ZN => n9714);
   U29498 : OAI222_X1 port map( A1 => n40895, A2 => n40551, B1 => n41279, B2 =>
                           n40544, C1 => n40540, C2 => n31945, ZN => n9713);
   U29499 : OAI222_X1 port map( A1 => n40901, A2 => n40551, B1 => n41285, B2 =>
                           n40544, C1 => n40540, C2 => n31944, ZN => n9712);
   U29500 : OAI222_X1 port map( A1 => n40907, A2 => n40551, B1 => n41291, B2 =>
                           n40544, C1 => n40540, C2 => n31943, ZN => n9711);
   U29501 : OAI222_X1 port map( A1 => n40913, A2 => n40550, B1 => n41297, B2 =>
                           n40543, C1 => n40540, C2 => n31942, ZN => n9710);
   U29502 : OAI222_X1 port map( A1 => n40919, A2 => n40550, B1 => n41303, B2 =>
                           n40543, C1 => n40540, C2 => n31941, ZN => n9709);
   U29503 : OAI222_X1 port map( A1 => n40925, A2 => n40550, B1 => n41309, B2 =>
                           n40543, C1 => n40540, C2 => n31940, ZN => n9708);
   U29504 : OAI222_X1 port map( A1 => n40931, A2 => n40550, B1 => n41315, B2 =>
                           n40543, C1 => n40540, C2 => n31939, ZN => n9707);
   U29505 : OAI222_X1 port map( A1 => n40937, A2 => n40550, B1 => n41321, B2 =>
                           n40543, C1 => n40540, C2 => n31938, ZN => n9706);
   U29506 : OAI222_X1 port map( A1 => n40943, A2 => n40550, B1 => n41327, B2 =>
                           n40543, C1 => n40540, C2 => n31937, ZN => n9705);
   U29507 : OAI222_X1 port map( A1 => n40949, A2 => n40550, B1 => n41333, B2 =>
                           n40543, C1 => n40540, C2 => n31936, ZN => n9704);
   U29508 : OAI222_X1 port map( A1 => n40961, A2 => n40550, B1 => n41345, B2 =>
                           n40543, C1 => n40540, C2 => n31934, ZN => n9702);
   U29509 : OAI222_X1 port map( A1 => n40624, A2 => n40494, B1 => n41008, B2 =>
                           n40487, C1 => n40476, C2 => n31930, ZN => n9566);
   U29510 : OAI222_X1 port map( A1 => n40630, A2 => n40494, B1 => n41014, B2 =>
                           n40487, C1 => n40476, C2 => n31929, ZN => n9565);
   U29511 : OAI222_X1 port map( A1 => n40636, A2 => n40494, B1 => n41020, B2 =>
                           n40487, C1 => n40476, C2 => n31928, ZN => n9564);
   U29512 : OAI222_X1 port map( A1 => n40642, A2 => n40494, B1 => n41026, B2 =>
                           n40487, C1 => n40476, C2 => n31927, ZN => n9563);
   U29513 : OAI222_X1 port map( A1 => n40648, A2 => n40494, B1 => n41032, B2 =>
                           n40487, C1 => n40476, C2 => n31926, ZN => n9562);
   U29514 : OAI222_X1 port map( A1 => n40654, A2 => n40494, B1 => n41038, B2 =>
                           n40487, C1 => n40476, C2 => n31925, ZN => n9561);
   U29515 : OAI222_X1 port map( A1 => n40660, A2 => n40494, B1 => n41044, B2 =>
                           n40487, C1 => n40476, C2 => n31924, ZN => n9560);
   U29516 : OAI222_X1 port map( A1 => n40666, A2 => n40494, B1 => n41050, B2 =>
                           n40487, C1 => n40476, C2 => n31923, ZN => n9559);
   U29517 : OAI222_X1 port map( A1 => n40672, A2 => n40494, B1 => n41056, B2 =>
                           n40487, C1 => n40477, C2 => n31922, ZN => n9558);
   U29518 : OAI222_X1 port map( A1 => n40678, A2 => n40494, B1 => n41062, B2 =>
                           n40487, C1 => n40477, C2 => n31921, ZN => n9557);
   U29519 : OAI222_X1 port map( A1 => n40684, A2 => n40494, B1 => n41068, B2 =>
                           n40487, C1 => n40477, C2 => n31920, ZN => n9556);
   U29520 : OAI222_X1 port map( A1 => n40690, A2 => n40494, B1 => n41074, B2 =>
                           n40487, C1 => n40478, C2 => n31919, ZN => n9555);
   U29521 : OAI222_X1 port map( A1 => n40696, A2 => n40493, B1 => n41080, B2 =>
                           n40486, C1 => n40477, C2 => n31918, ZN => n9554);
   U29522 : OAI222_X1 port map( A1 => n40702, A2 => n40493, B1 => n41086, B2 =>
                           n40486, C1 => n40477, C2 => n31917, ZN => n9553);
   U29523 : OAI222_X1 port map( A1 => n40708, A2 => n40493, B1 => n41092, B2 =>
                           n40486, C1 => n40477, C2 => n31916, ZN => n9552);
   U29524 : OAI222_X1 port map( A1 => n40714, A2 => n40493, B1 => n41098, B2 =>
                           n40486, C1 => n40477, C2 => n31915, ZN => n9551);
   U29525 : OAI222_X1 port map( A1 => n40720, A2 => n40493, B1 => n41104, B2 =>
                           n40486, C1 => n40477, C2 => n31914, ZN => n9550);
   U29526 : OAI222_X1 port map( A1 => n40726, A2 => n40493, B1 => n41110, B2 =>
                           n40486, C1 => n40477, C2 => n31913, ZN => n9549);
   U29527 : OAI222_X1 port map( A1 => n40732, A2 => n40493, B1 => n41116, B2 =>
                           n40486, C1 => n40477, C2 => n31912, ZN => n9548);
   U29528 : OAI222_X1 port map( A1 => n40738, A2 => n40493, B1 => n41122, B2 =>
                           n40486, C1 => n40477, C2 => n31911, ZN => n9547);
   U29529 : OAI222_X1 port map( A1 => n40744, A2 => n40493, B1 => n41128, B2 =>
                           n40486, C1 => n40477, C2 => n31910, ZN => n9546);
   U29530 : OAI222_X1 port map( A1 => n40750, A2 => n40493, B1 => n41134, B2 =>
                           n40486, C1 => n40478, C2 => n31909, ZN => n9545);
   U29531 : OAI222_X1 port map( A1 => n40756, A2 => n40493, B1 => n41140, B2 =>
                           n40486, C1 => n40478, C2 => n31908, ZN => n9544);
   U29532 : OAI222_X1 port map( A1 => n40762, A2 => n40493, B1 => n41146, B2 =>
                           n40486, C1 => n40478, C2 => n31907, ZN => n9543);
   U29533 : OAI222_X1 port map( A1 => n40768, A2 => n40492, B1 => n41152, B2 =>
                           n40485, C1 => n40478, C2 => n31906, ZN => n9542);
   U29534 : OAI222_X1 port map( A1 => n40774, A2 => n40492, B1 => n41158, B2 =>
                           n40485, C1 => n40478, C2 => n31905, ZN => n9541);
   U29535 : OAI222_X1 port map( A1 => n40780, A2 => n40492, B1 => n41164, B2 =>
                           n40485, C1 => n40478, C2 => n31904, ZN => n9540);
   U29536 : OAI222_X1 port map( A1 => n40786, A2 => n40492, B1 => n41170, B2 =>
                           n40485, C1 => n40478, C2 => n31903, ZN => n9539);
   U29537 : OAI222_X1 port map( A1 => n40792, A2 => n40492, B1 => n41176, B2 =>
                           n40485, C1 => n40478, C2 => n31902, ZN => n9538);
   U29538 : OAI222_X1 port map( A1 => n40798, A2 => n40492, B1 => n41182, B2 =>
                           n40485, C1 => n40478, C2 => n31901, ZN => n9537);
   U29539 : OAI222_X1 port map( A1 => n40804, A2 => n40492, B1 => n41188, B2 =>
                           n40485, C1 => n40478, C2 => n31900, ZN => n9536);
   U29540 : OAI222_X1 port map( A1 => n40810, A2 => n40492, B1 => n41194, B2 =>
                           n40485, C1 => n40478, C2 => n31899, ZN => n9535);
   U29541 : OAI222_X1 port map( A1 => n40816, A2 => n40492, B1 => n41200, B2 =>
                           n40485, C1 => n40479, C2 => n31898, ZN => n9534);
   U29542 : OAI222_X1 port map( A1 => n40822, A2 => n40492, B1 => n41206, B2 =>
                           n40485, C1 => n40479, C2 => n31897, ZN => n9533);
   U29543 : OAI222_X1 port map( A1 => n40828, A2 => n40492, B1 => n41212, B2 =>
                           n40485, C1 => n40479, C2 => n31896, ZN => n9532);
   U29544 : OAI222_X1 port map( A1 => n40834, A2 => n40492, B1 => n41218, B2 =>
                           n40485, C1 => n40479, C2 => n31895, ZN => n9531);
   U29545 : OAI222_X1 port map( A1 => n40840, A2 => n40491, B1 => n41224, B2 =>
                           n40484, C1 => n40479, C2 => n31894, ZN => n9530);
   U29546 : OAI222_X1 port map( A1 => n40846, A2 => n40491, B1 => n41230, B2 =>
                           n40484, C1 => n40479, C2 => n31893, ZN => n9529);
   U29547 : OAI222_X1 port map( A1 => n40852, A2 => n40491, B1 => n41236, B2 =>
                           n40484, C1 => n40479, C2 => n31892, ZN => n9528);
   U29548 : OAI222_X1 port map( A1 => n40858, A2 => n40491, B1 => n41242, B2 =>
                           n40484, C1 => n40479, C2 => n31891, ZN => n9527);
   U29549 : OAI222_X1 port map( A1 => n40864, A2 => n40491, B1 => n41248, B2 =>
                           n40484, C1 => n40479, C2 => n31890, ZN => n9526);
   U29550 : OAI222_X1 port map( A1 => n40870, A2 => n40491, B1 => n41254, B2 =>
                           n40484, C1 => n40479, C2 => n31889, ZN => n9525);
   U29551 : OAI222_X1 port map( A1 => n40876, A2 => n40491, B1 => n41260, B2 =>
                           n40484, C1 => n40479, C2 => n31888, ZN => n9524);
   U29552 : OAI222_X1 port map( A1 => n40882, A2 => n40491, B1 => n41266, B2 =>
                           n40484, C1 => n40479, C2 => n31887, ZN => n9523);
   U29553 : OAI222_X1 port map( A1 => n40888, A2 => n40491, B1 => n41272, B2 =>
                           n40484, C1 => n40480, C2 => n31886, ZN => n9522);
   U29554 : OAI222_X1 port map( A1 => n40894, A2 => n40491, B1 => n41278, B2 =>
                           n40484, C1 => n40480, C2 => n31885, ZN => n9521);
   U29555 : OAI222_X1 port map( A1 => n40900, A2 => n40491, B1 => n41284, B2 =>
                           n40484, C1 => n40480, C2 => n31884, ZN => n9520);
   U29556 : OAI222_X1 port map( A1 => n40906, A2 => n40491, B1 => n41290, B2 =>
                           n40484, C1 => n40480, C2 => n31883, ZN => n9519);
   U29557 : OAI222_X1 port map( A1 => n40912, A2 => n40490, B1 => n41296, B2 =>
                           n40483, C1 => n40480, C2 => n31882, ZN => n9518);
   U29558 : OAI222_X1 port map( A1 => n40918, A2 => n40490, B1 => n41302, B2 =>
                           n40483, C1 => n40480, C2 => n31881, ZN => n9517);
   U29559 : OAI222_X1 port map( A1 => n40924, A2 => n40490, B1 => n41308, B2 =>
                           n40483, C1 => n40480, C2 => n31880, ZN => n9516);
   U29560 : OAI222_X1 port map( A1 => n40930, A2 => n40490, B1 => n41314, B2 =>
                           n40483, C1 => n40480, C2 => n31879, ZN => n9515);
   U29561 : OAI222_X1 port map( A1 => n40936, A2 => n40490, B1 => n41320, B2 =>
                           n40483, C1 => n40480, C2 => n31878, ZN => n9514);
   U29562 : OAI222_X1 port map( A1 => n40942, A2 => n40490, B1 => n41326, B2 =>
                           n40483, C1 => n40480, C2 => n31877, ZN => n9513);
   U29563 : OAI222_X1 port map( A1 => n40948, A2 => n40490, B1 => n41332, B2 =>
                           n40483, C1 => n40480, C2 => n31876, ZN => n9512);
   U29564 : OAI222_X1 port map( A1 => n40960, A2 => n40490, B1 => n41344, B2 =>
                           n40483, C1 => n40480, C2 => n31874, ZN => n9510);
   U29565 : OAI222_X1 port map( A1 => n40624, A2 => n40474, B1 => n41008, B2 =>
                           n40467, C1 => n40456, C2 => n31870, ZN => n9502);
   U29566 : OAI222_X1 port map( A1 => n40630, A2 => n40474, B1 => n41014, B2 =>
                           n40467, C1 => n40456, C2 => n31869, ZN => n9501);
   U29567 : OAI222_X1 port map( A1 => n40636, A2 => n40474, B1 => n41020, B2 =>
                           n40467, C1 => n40456, C2 => n31868, ZN => n9500);
   U29568 : OAI222_X1 port map( A1 => n40642, A2 => n40474, B1 => n41026, B2 =>
                           n40467, C1 => n40456, C2 => n31867, ZN => n9499);
   U29569 : OAI222_X1 port map( A1 => n40648, A2 => n40474, B1 => n41032, B2 =>
                           n40467, C1 => n40456, C2 => n31866, ZN => n9498);
   U29570 : OAI222_X1 port map( A1 => n40654, A2 => n40474, B1 => n41038, B2 =>
                           n40467, C1 => n40456, C2 => n31865, ZN => n9497);
   U29571 : OAI222_X1 port map( A1 => n40660, A2 => n40474, B1 => n41044, B2 =>
                           n40467, C1 => n40456, C2 => n31864, ZN => n9496);
   U29572 : OAI222_X1 port map( A1 => n40666, A2 => n40474, B1 => n41050, B2 =>
                           n40467, C1 => n40456, C2 => n31863, ZN => n9495);
   U29573 : OAI222_X1 port map( A1 => n40672, A2 => n40474, B1 => n41056, B2 =>
                           n40467, C1 => n40457, C2 => n31862, ZN => n9494);
   U29574 : OAI222_X1 port map( A1 => n40678, A2 => n40474, B1 => n41062, B2 =>
                           n40467, C1 => n40457, C2 => n31861, ZN => n9493);
   U29575 : OAI222_X1 port map( A1 => n40684, A2 => n40474, B1 => n41068, B2 =>
                           n40467, C1 => n40457, C2 => n31860, ZN => n9492);
   U29576 : OAI222_X1 port map( A1 => n40690, A2 => n40474, B1 => n41074, B2 =>
                           n40467, C1 => n40458, C2 => n31859, ZN => n9491);
   U29577 : OAI222_X1 port map( A1 => n40696, A2 => n40473, B1 => n41080, B2 =>
                           n40466, C1 => n40457, C2 => n31858, ZN => n9490);
   U29578 : OAI222_X1 port map( A1 => n40702, A2 => n40473, B1 => n41086, B2 =>
                           n40466, C1 => n40457, C2 => n31857, ZN => n9489);
   U29579 : OAI222_X1 port map( A1 => n40708, A2 => n40473, B1 => n41092, B2 =>
                           n40466, C1 => n40457, C2 => n31856, ZN => n9488);
   U29580 : OAI222_X1 port map( A1 => n40714, A2 => n40473, B1 => n41098, B2 =>
                           n40466, C1 => n40457, C2 => n31855, ZN => n9487);
   U29581 : OAI222_X1 port map( A1 => n40720, A2 => n40473, B1 => n41104, B2 =>
                           n40466, C1 => n40457, C2 => n31854, ZN => n9486);
   U29582 : OAI222_X1 port map( A1 => n40726, A2 => n40473, B1 => n41110, B2 =>
                           n40466, C1 => n40457, C2 => n31853, ZN => n9485);
   U29583 : OAI222_X1 port map( A1 => n40732, A2 => n40473, B1 => n41116, B2 =>
                           n40466, C1 => n40457, C2 => n31852, ZN => n9484);
   U29584 : OAI222_X1 port map( A1 => n40738, A2 => n40473, B1 => n41122, B2 =>
                           n40466, C1 => n40457, C2 => n31851, ZN => n9483);
   U29585 : OAI222_X1 port map( A1 => n40744, A2 => n40473, B1 => n41128, B2 =>
                           n40466, C1 => n40457, C2 => n31850, ZN => n9482);
   U29586 : OAI222_X1 port map( A1 => n40750, A2 => n40473, B1 => n41134, B2 =>
                           n40466, C1 => n40458, C2 => n31849, ZN => n9481);
   U29587 : OAI222_X1 port map( A1 => n40756, A2 => n40473, B1 => n41140, B2 =>
                           n40466, C1 => n40458, C2 => n31848, ZN => n9480);
   U29588 : OAI222_X1 port map( A1 => n40762, A2 => n40473, B1 => n41146, B2 =>
                           n40466, C1 => n40458, C2 => n31847, ZN => n9479);
   U29589 : OAI222_X1 port map( A1 => n40768, A2 => n40472, B1 => n41152, B2 =>
                           n40465, C1 => n40458, C2 => n31846, ZN => n9478);
   U29590 : OAI222_X1 port map( A1 => n40774, A2 => n40472, B1 => n41158, B2 =>
                           n40465, C1 => n40458, C2 => n31845, ZN => n9477);
   U29591 : OAI222_X1 port map( A1 => n40780, A2 => n40472, B1 => n41164, B2 =>
                           n40465, C1 => n40458, C2 => n31844, ZN => n9476);
   U29592 : OAI222_X1 port map( A1 => n40786, A2 => n40472, B1 => n41170, B2 =>
                           n40465, C1 => n40458, C2 => n31843, ZN => n9475);
   U29593 : OAI222_X1 port map( A1 => n40792, A2 => n40472, B1 => n41176, B2 =>
                           n40465, C1 => n40458, C2 => n31842, ZN => n9474);
   U29594 : OAI222_X1 port map( A1 => n40798, A2 => n40472, B1 => n41182, B2 =>
                           n40465, C1 => n40458, C2 => n31841, ZN => n9473);
   U29595 : OAI222_X1 port map( A1 => n40804, A2 => n40472, B1 => n41188, B2 =>
                           n40465, C1 => n40458, C2 => n31840, ZN => n9472);
   U29596 : OAI222_X1 port map( A1 => n40810, A2 => n40472, B1 => n41194, B2 =>
                           n40465, C1 => n40458, C2 => n31839, ZN => n9471);
   U29597 : OAI222_X1 port map( A1 => n40816, A2 => n40472, B1 => n41200, B2 =>
                           n40465, C1 => n40459, C2 => n31838, ZN => n9470);
   U29598 : OAI222_X1 port map( A1 => n40822, A2 => n40472, B1 => n41206, B2 =>
                           n40465, C1 => n40459, C2 => n31837, ZN => n9469);
   U29599 : OAI222_X1 port map( A1 => n40828, A2 => n40472, B1 => n41212, B2 =>
                           n40465, C1 => n40459, C2 => n31836, ZN => n9468);
   U29600 : OAI222_X1 port map( A1 => n40834, A2 => n40472, B1 => n41218, B2 =>
                           n40465, C1 => n40459, C2 => n31835, ZN => n9467);
   U29601 : OAI222_X1 port map( A1 => n40840, A2 => n40471, B1 => n41224, B2 =>
                           n40464, C1 => n40459, C2 => n31834, ZN => n9466);
   U29602 : OAI222_X1 port map( A1 => n40846, A2 => n40471, B1 => n41230, B2 =>
                           n40464, C1 => n40459, C2 => n31833, ZN => n9465);
   U29603 : OAI222_X1 port map( A1 => n40852, A2 => n40471, B1 => n41236, B2 =>
                           n40464, C1 => n40459, C2 => n31832, ZN => n9464);
   U29604 : OAI222_X1 port map( A1 => n40858, A2 => n40471, B1 => n41242, B2 =>
                           n40464, C1 => n40459, C2 => n31831, ZN => n9463);
   U29605 : OAI222_X1 port map( A1 => n40864, A2 => n40471, B1 => n41248, B2 =>
                           n40464, C1 => n40459, C2 => n31830, ZN => n9462);
   U29606 : OAI222_X1 port map( A1 => n40870, A2 => n40471, B1 => n41254, B2 =>
                           n40464, C1 => n40459, C2 => n31829, ZN => n9461);
   U29607 : OAI222_X1 port map( A1 => n40876, A2 => n40471, B1 => n41260, B2 =>
                           n40464, C1 => n40459, C2 => n31828, ZN => n9460);
   U29608 : OAI222_X1 port map( A1 => n40882, A2 => n40471, B1 => n41266, B2 =>
                           n40464, C1 => n40459, C2 => n31827, ZN => n9459);
   U29609 : OAI222_X1 port map( A1 => n40888, A2 => n40471, B1 => n41272, B2 =>
                           n40464, C1 => n40460, C2 => n31826, ZN => n9458);
   U29610 : OAI222_X1 port map( A1 => n40894, A2 => n40471, B1 => n41278, B2 =>
                           n40464, C1 => n40460, C2 => n31825, ZN => n9457);
   U29611 : OAI222_X1 port map( A1 => n40900, A2 => n40471, B1 => n41284, B2 =>
                           n40464, C1 => n40460, C2 => n31824, ZN => n9456);
   U29612 : OAI222_X1 port map( A1 => n40906, A2 => n40471, B1 => n41290, B2 =>
                           n40464, C1 => n40460, C2 => n31823, ZN => n9455);
   U29613 : OAI222_X1 port map( A1 => n40912, A2 => n40470, B1 => n41296, B2 =>
                           n40463, C1 => n40460, C2 => n31822, ZN => n9454);
   U29614 : OAI222_X1 port map( A1 => n40918, A2 => n40470, B1 => n41302, B2 =>
                           n40463, C1 => n40460, C2 => n31821, ZN => n9453);
   U29615 : OAI222_X1 port map( A1 => n40924, A2 => n40470, B1 => n41308, B2 =>
                           n40463, C1 => n40460, C2 => n31820, ZN => n9452);
   U29616 : OAI222_X1 port map( A1 => n40930, A2 => n40470, B1 => n41314, B2 =>
                           n40463, C1 => n40460, C2 => n31819, ZN => n9451);
   U29617 : OAI222_X1 port map( A1 => n40936, A2 => n40470, B1 => n41320, B2 =>
                           n40463, C1 => n40460, C2 => n31818, ZN => n9450);
   U29618 : OAI222_X1 port map( A1 => n40942, A2 => n40470, B1 => n41326, B2 =>
                           n40463, C1 => n40460, C2 => n31817, ZN => n9449);
   U29619 : OAI222_X1 port map( A1 => n40948, A2 => n40470, B1 => n41332, B2 =>
                           n40463, C1 => n40460, C2 => n31816, ZN => n9448);
   U29620 : OAI222_X1 port map( A1 => n40960, A2 => n40470, B1 => n41344, B2 =>
                           n40463, C1 => n40460, C2 => n31814, ZN => n9446);
   U29621 : OAI222_X1 port map( A1 => n40624, A2 => n40454, B1 => n41008, B2 =>
                           n40447, C1 => n40436, C2 => n31810, ZN => n9438);
   U29622 : OAI222_X1 port map( A1 => n40630, A2 => n40454, B1 => n41014, B2 =>
                           n40447, C1 => n40436, C2 => n31809, ZN => n9437);
   U29623 : OAI222_X1 port map( A1 => n40636, A2 => n40454, B1 => n41020, B2 =>
                           n40447, C1 => n40436, C2 => n31808, ZN => n9436);
   U29624 : OAI222_X1 port map( A1 => n40642, A2 => n40454, B1 => n41026, B2 =>
                           n40447, C1 => n40436, C2 => n31807, ZN => n9435);
   U29625 : OAI222_X1 port map( A1 => n40648, A2 => n40454, B1 => n41032, B2 =>
                           n40447, C1 => n40436, C2 => n31806, ZN => n9434);
   U29626 : OAI222_X1 port map( A1 => n40654, A2 => n40454, B1 => n41038, B2 =>
                           n40447, C1 => n40436, C2 => n31805, ZN => n9433);
   U29627 : OAI222_X1 port map( A1 => n40660, A2 => n40454, B1 => n41044, B2 =>
                           n40447, C1 => n40436, C2 => n31804, ZN => n9432);
   U29628 : OAI222_X1 port map( A1 => n40666, A2 => n40454, B1 => n41050, B2 =>
                           n40447, C1 => n40436, C2 => n31803, ZN => n9431);
   U29629 : OAI222_X1 port map( A1 => n40672, A2 => n40454, B1 => n41056, B2 =>
                           n40447, C1 => n40437, C2 => n31802, ZN => n9430);
   U29630 : OAI222_X1 port map( A1 => n40678, A2 => n40454, B1 => n41062, B2 =>
                           n40447, C1 => n40437, C2 => n31801, ZN => n9429);
   U29631 : OAI222_X1 port map( A1 => n40684, A2 => n40454, B1 => n41068, B2 =>
                           n40447, C1 => n40437, C2 => n31800, ZN => n9428);
   U29632 : OAI222_X1 port map( A1 => n40690, A2 => n40454, B1 => n41074, B2 =>
                           n40447, C1 => n40438, C2 => n31799, ZN => n9427);
   U29633 : OAI222_X1 port map( A1 => n40696, A2 => n40453, B1 => n41080, B2 =>
                           n40446, C1 => n40437, C2 => n31798, ZN => n9426);
   U29634 : OAI222_X1 port map( A1 => n40702, A2 => n40453, B1 => n41086, B2 =>
                           n40446, C1 => n40437, C2 => n31797, ZN => n9425);
   U29635 : OAI222_X1 port map( A1 => n40708, A2 => n40453, B1 => n41092, B2 =>
                           n40446, C1 => n40437, C2 => n31796, ZN => n9424);
   U29636 : OAI222_X1 port map( A1 => n40714, A2 => n40453, B1 => n41098, B2 =>
                           n40446, C1 => n40437, C2 => n31795, ZN => n9423);
   U29637 : OAI222_X1 port map( A1 => n40720, A2 => n40453, B1 => n41104, B2 =>
                           n40446, C1 => n40437, C2 => n31794, ZN => n9422);
   U29638 : OAI222_X1 port map( A1 => n40726, A2 => n40453, B1 => n41110, B2 =>
                           n40446, C1 => n40437, C2 => n31793, ZN => n9421);
   U29639 : OAI222_X1 port map( A1 => n40732, A2 => n40453, B1 => n41116, B2 =>
                           n40446, C1 => n40437, C2 => n31792, ZN => n9420);
   U29640 : OAI222_X1 port map( A1 => n40738, A2 => n40453, B1 => n41122, B2 =>
                           n40446, C1 => n40437, C2 => n31791, ZN => n9419);
   U29641 : OAI222_X1 port map( A1 => n40744, A2 => n40453, B1 => n41128, B2 =>
                           n40446, C1 => n40437, C2 => n31790, ZN => n9418);
   U29642 : OAI222_X1 port map( A1 => n40750, A2 => n40453, B1 => n41134, B2 =>
                           n40446, C1 => n40438, C2 => n31789, ZN => n9417);
   U29643 : OAI222_X1 port map( A1 => n40756, A2 => n40453, B1 => n41140, B2 =>
                           n40446, C1 => n40438, C2 => n31788, ZN => n9416);
   U29644 : OAI222_X1 port map( A1 => n40762, A2 => n40453, B1 => n41146, B2 =>
                           n40446, C1 => n40438, C2 => n31787, ZN => n9415);
   U29645 : OAI222_X1 port map( A1 => n40768, A2 => n40452, B1 => n41152, B2 =>
                           n40445, C1 => n40438, C2 => n31786, ZN => n9414);
   U29646 : OAI222_X1 port map( A1 => n40774, A2 => n40452, B1 => n41158, B2 =>
                           n40445, C1 => n40438, C2 => n31785, ZN => n9413);
   U29647 : OAI222_X1 port map( A1 => n40780, A2 => n40452, B1 => n41164, B2 =>
                           n40445, C1 => n40438, C2 => n31784, ZN => n9412);
   U29648 : OAI222_X1 port map( A1 => n40786, A2 => n40452, B1 => n41170, B2 =>
                           n40445, C1 => n40438, C2 => n31783, ZN => n9411);
   U29649 : OAI222_X1 port map( A1 => n40792, A2 => n40452, B1 => n41176, B2 =>
                           n40445, C1 => n40438, C2 => n31782, ZN => n9410);
   U29650 : OAI222_X1 port map( A1 => n40798, A2 => n40452, B1 => n41182, B2 =>
                           n40445, C1 => n40438, C2 => n31781, ZN => n9409);
   U29651 : OAI222_X1 port map( A1 => n40804, A2 => n40452, B1 => n41188, B2 =>
                           n40445, C1 => n40438, C2 => n31780, ZN => n9408);
   U29652 : OAI222_X1 port map( A1 => n40810, A2 => n40452, B1 => n41194, B2 =>
                           n40445, C1 => n40438, C2 => n31779, ZN => n9407);
   U29653 : OAI222_X1 port map( A1 => n40816, A2 => n40452, B1 => n41200, B2 =>
                           n40445, C1 => n40439, C2 => n31778, ZN => n9406);
   U29654 : OAI222_X1 port map( A1 => n40822, A2 => n40452, B1 => n41206, B2 =>
                           n40445, C1 => n40439, C2 => n31777, ZN => n9405);
   U29655 : OAI222_X1 port map( A1 => n40828, A2 => n40452, B1 => n41212, B2 =>
                           n40445, C1 => n40439, C2 => n31776, ZN => n9404);
   U29656 : OAI222_X1 port map( A1 => n40834, A2 => n40452, B1 => n41218, B2 =>
                           n40445, C1 => n40439, C2 => n31775, ZN => n9403);
   U29657 : OAI222_X1 port map( A1 => n40840, A2 => n40451, B1 => n41224, B2 =>
                           n40444, C1 => n40439, C2 => n31774, ZN => n9402);
   U29658 : OAI222_X1 port map( A1 => n40846, A2 => n40451, B1 => n41230, B2 =>
                           n40444, C1 => n40439, C2 => n31773, ZN => n9401);
   U29659 : OAI222_X1 port map( A1 => n40852, A2 => n40451, B1 => n41236, B2 =>
                           n40444, C1 => n40439, C2 => n31772, ZN => n9400);
   U29660 : OAI222_X1 port map( A1 => n40858, A2 => n40451, B1 => n41242, B2 =>
                           n40444, C1 => n40439, C2 => n31771, ZN => n9399);
   U29661 : OAI222_X1 port map( A1 => n40864, A2 => n40451, B1 => n41248, B2 =>
                           n40444, C1 => n40439, C2 => n31770, ZN => n9398);
   U29662 : OAI222_X1 port map( A1 => n40870, A2 => n40451, B1 => n41254, B2 =>
                           n40444, C1 => n40439, C2 => n31769, ZN => n9397);
   U29663 : OAI222_X1 port map( A1 => n40876, A2 => n40451, B1 => n41260, B2 =>
                           n40444, C1 => n40439, C2 => n31768, ZN => n9396);
   U29664 : OAI222_X1 port map( A1 => n40882, A2 => n40451, B1 => n41266, B2 =>
                           n40444, C1 => n40439, C2 => n31767, ZN => n9395);
   U29665 : OAI222_X1 port map( A1 => n40888, A2 => n40451, B1 => n41272, B2 =>
                           n40444, C1 => n40440, C2 => n31766, ZN => n9394);
   U29666 : OAI222_X1 port map( A1 => n40894, A2 => n40451, B1 => n41278, B2 =>
                           n40444, C1 => n40440, C2 => n31765, ZN => n9393);
   U29667 : OAI222_X1 port map( A1 => n40900, A2 => n40451, B1 => n41284, B2 =>
                           n40444, C1 => n40440, C2 => n31764, ZN => n9392);
   U29668 : OAI222_X1 port map( A1 => n40906, A2 => n40451, B1 => n41290, B2 =>
                           n40444, C1 => n40440, C2 => n31763, ZN => n9391);
   U29669 : OAI222_X1 port map( A1 => n40912, A2 => n40450, B1 => n41296, B2 =>
                           n40443, C1 => n40440, C2 => n31762, ZN => n9390);
   U29670 : OAI222_X1 port map( A1 => n40918, A2 => n40450, B1 => n41302, B2 =>
                           n40443, C1 => n40440, C2 => n31761, ZN => n9389);
   U29671 : OAI222_X1 port map( A1 => n40924, A2 => n40450, B1 => n41308, B2 =>
                           n40443, C1 => n40440, C2 => n31760, ZN => n9388);
   U29672 : OAI222_X1 port map( A1 => n40930, A2 => n40450, B1 => n41314, B2 =>
                           n40443, C1 => n40440, C2 => n31759, ZN => n9387);
   U29673 : OAI222_X1 port map( A1 => n40936, A2 => n40450, B1 => n41320, B2 =>
                           n40443, C1 => n40440, C2 => n31758, ZN => n9386);
   U29674 : OAI222_X1 port map( A1 => n40942, A2 => n40450, B1 => n41326, B2 =>
                           n40443, C1 => n40440, C2 => n31757, ZN => n9385);
   U29675 : OAI222_X1 port map( A1 => n40948, A2 => n40450, B1 => n41332, B2 =>
                           n40443, C1 => n40440, C2 => n31756, ZN => n9384);
   U29676 : OAI222_X1 port map( A1 => n40960, A2 => n40450, B1 => n41344, B2 =>
                           n40443, C1 => n40440, C2 => n31754, ZN => n9382);
   U29677 : OAI222_X1 port map( A1 => n40600, A2 => n40395, B1 => n40984, B2 =>
                           n40388, C1 => n40376, C2 => n31750, ZN => n9250);
   U29678 : OAI222_X1 port map( A1 => n40606, A2 => n40395, B1 => n40990, B2 =>
                           n40388, C1 => n40376, C2 => n31749, ZN => n9249);
   U29679 : OAI222_X1 port map( A1 => n40612, A2 => n40395, B1 => n40996, B2 =>
                           n40388, C1 => n40376, C2 => n31748, ZN => n9248);
   U29680 : OAI222_X1 port map( A1 => n40618, A2 => n40395, B1 => n41002, B2 =>
                           n40388, C1 => n40376, C2 => n31747, ZN => n9247);
   U29681 : OAI222_X1 port map( A1 => n40624, A2 => n40394, B1 => n41008, B2 =>
                           n40387, C1 => n40376, C2 => n31746, ZN => n9246);
   U29682 : OAI222_X1 port map( A1 => n40630, A2 => n40394, B1 => n41014, B2 =>
                           n40387, C1 => n40376, C2 => n31745, ZN => n9245);
   U29683 : OAI222_X1 port map( A1 => n40636, A2 => n40394, B1 => n41020, B2 =>
                           n40387, C1 => n40376, C2 => n31744, ZN => n9244);
   U29684 : OAI222_X1 port map( A1 => n40642, A2 => n40394, B1 => n41026, B2 =>
                           n40387, C1 => n40376, C2 => n31743, ZN => n9243);
   U29685 : OAI222_X1 port map( A1 => n40648, A2 => n40394, B1 => n41032, B2 =>
                           n40387, C1 => n40376, C2 => n31742, ZN => n9242);
   U29686 : OAI222_X1 port map( A1 => n40654, A2 => n40394, B1 => n41038, B2 =>
                           n40387, C1 => n40376, C2 => n31741, ZN => n9241);
   U29687 : OAI222_X1 port map( A1 => n40660, A2 => n40394, B1 => n41044, B2 =>
                           n40387, C1 => n40376, C2 => n31740, ZN => n9240);
   U29688 : OAI222_X1 port map( A1 => n40666, A2 => n40394, B1 => n41050, B2 =>
                           n40387, C1 => n40376, C2 => n31739, ZN => n9239);
   U29689 : OAI222_X1 port map( A1 => n40672, A2 => n40394, B1 => n41056, B2 =>
                           n40387, C1 => n40377, C2 => n31738, ZN => n9238);
   U29690 : OAI222_X1 port map( A1 => n40678, A2 => n40394, B1 => n41062, B2 =>
                           n40387, C1 => n40377, C2 => n31737, ZN => n9237);
   U29691 : OAI222_X1 port map( A1 => n40684, A2 => n40394, B1 => n41068, B2 =>
                           n40387, C1 => n40377, C2 => n31736, ZN => n9236);
   U29692 : OAI222_X1 port map( A1 => n40690, A2 => n40394, B1 => n41074, B2 =>
                           n40387, C1 => n40378, C2 => n31735, ZN => n9235);
   U29693 : OAI222_X1 port map( A1 => n40696, A2 => n40393, B1 => n41080, B2 =>
                           n40386, C1 => n40377, C2 => n31734, ZN => n9234);
   U29694 : OAI222_X1 port map( A1 => n40702, A2 => n40393, B1 => n41086, B2 =>
                           n40386, C1 => n40377, C2 => n31733, ZN => n9233);
   U29695 : OAI222_X1 port map( A1 => n40708, A2 => n40393, B1 => n41092, B2 =>
                           n40386, C1 => n40377, C2 => n31732, ZN => n9232);
   U29696 : OAI222_X1 port map( A1 => n40714, A2 => n40393, B1 => n41098, B2 =>
                           n40386, C1 => n40377, C2 => n31731, ZN => n9231);
   U29697 : OAI222_X1 port map( A1 => n40720, A2 => n40393, B1 => n41104, B2 =>
                           n40386, C1 => n40377, C2 => n31730, ZN => n9230);
   U29698 : OAI222_X1 port map( A1 => n40726, A2 => n40393, B1 => n41110, B2 =>
                           n40386, C1 => n40377, C2 => n31729, ZN => n9229);
   U29699 : OAI222_X1 port map( A1 => n40732, A2 => n40393, B1 => n41116, B2 =>
                           n40386, C1 => n40377, C2 => n31728, ZN => n9228);
   U29700 : OAI222_X1 port map( A1 => n40738, A2 => n40393, B1 => n41122, B2 =>
                           n40386, C1 => n40377, C2 => n31727, ZN => n9227);
   U29701 : OAI222_X1 port map( A1 => n40744, A2 => n40393, B1 => n41128, B2 =>
                           n40386, C1 => n40377, C2 => n31726, ZN => n9226);
   U29702 : OAI222_X1 port map( A1 => n40750, A2 => n40393, B1 => n41134, B2 =>
                           n40386, C1 => n40378, C2 => n31725, ZN => n9225);
   U29703 : OAI222_X1 port map( A1 => n40756, A2 => n40393, B1 => n41140, B2 =>
                           n40386, C1 => n40378, C2 => n31724, ZN => n9224);
   U29704 : OAI222_X1 port map( A1 => n40762, A2 => n40393, B1 => n41146, B2 =>
                           n40386, C1 => n40378, C2 => n31723, ZN => n9223);
   U29705 : OAI222_X1 port map( A1 => n40768, A2 => n40392, B1 => n41152, B2 =>
                           n40385, C1 => n40378, C2 => n31722, ZN => n9222);
   U29706 : OAI222_X1 port map( A1 => n40774, A2 => n40392, B1 => n41158, B2 =>
                           n40385, C1 => n40378, C2 => n31721, ZN => n9221);
   U29707 : OAI222_X1 port map( A1 => n40780, A2 => n40392, B1 => n41164, B2 =>
                           n40385, C1 => n40378, C2 => n31720, ZN => n9220);
   U29708 : OAI222_X1 port map( A1 => n40786, A2 => n40392, B1 => n41170, B2 =>
                           n40385, C1 => n40378, C2 => n31719, ZN => n9219);
   U29709 : OAI222_X1 port map( A1 => n40792, A2 => n40392, B1 => n41176, B2 =>
                           n40385, C1 => n40378, C2 => n31718, ZN => n9218);
   U29710 : OAI222_X1 port map( A1 => n40798, A2 => n40392, B1 => n41182, B2 =>
                           n40385, C1 => n40378, C2 => n31717, ZN => n9217);
   U29711 : OAI222_X1 port map( A1 => n40804, A2 => n40392, B1 => n41188, B2 =>
                           n40385, C1 => n40378, C2 => n31716, ZN => n9216);
   U29712 : OAI222_X1 port map( A1 => n40810, A2 => n40392, B1 => n41194, B2 =>
                           n40385, C1 => n40378, C2 => n31715, ZN => n9215);
   U29713 : OAI222_X1 port map( A1 => n40816, A2 => n40392, B1 => n41200, B2 =>
                           n40385, C1 => n40379, C2 => n31714, ZN => n9214);
   U29714 : OAI222_X1 port map( A1 => n40822, A2 => n40392, B1 => n41206, B2 =>
                           n40385, C1 => n40379, C2 => n31713, ZN => n9213);
   U29715 : OAI222_X1 port map( A1 => n40828, A2 => n40392, B1 => n41212, B2 =>
                           n40385, C1 => n40379, C2 => n31712, ZN => n9212);
   U29716 : OAI222_X1 port map( A1 => n40834, A2 => n40392, B1 => n41218, B2 =>
                           n40385, C1 => n40379, C2 => n31711, ZN => n9211);
   U29717 : OAI222_X1 port map( A1 => n40840, A2 => n40391, B1 => n41224, B2 =>
                           n40384, C1 => n40379, C2 => n31710, ZN => n9210);
   U29718 : OAI222_X1 port map( A1 => n40846, A2 => n40391, B1 => n41230, B2 =>
                           n40384, C1 => n40379, C2 => n31709, ZN => n9209);
   U29719 : OAI222_X1 port map( A1 => n40852, A2 => n40391, B1 => n41236, B2 =>
                           n40384, C1 => n40379, C2 => n31708, ZN => n9208);
   U29720 : OAI222_X1 port map( A1 => n40858, A2 => n40391, B1 => n41242, B2 =>
                           n40384, C1 => n40379, C2 => n31707, ZN => n9207);
   U29721 : OAI222_X1 port map( A1 => n40864, A2 => n40391, B1 => n41248, B2 =>
                           n40384, C1 => n40379, C2 => n31706, ZN => n9206);
   U29722 : OAI222_X1 port map( A1 => n40870, A2 => n40391, B1 => n41254, B2 =>
                           n40384, C1 => n40379, C2 => n31705, ZN => n9205);
   U29723 : OAI222_X1 port map( A1 => n40876, A2 => n40391, B1 => n41260, B2 =>
                           n40384, C1 => n40379, C2 => n31704, ZN => n9204);
   U29724 : OAI222_X1 port map( A1 => n40882, A2 => n40391, B1 => n41266, B2 =>
                           n40384, C1 => n40379, C2 => n31703, ZN => n9203);
   U29725 : OAI222_X1 port map( A1 => n40888, A2 => n40391, B1 => n41272, B2 =>
                           n40384, C1 => n40380, C2 => n31702, ZN => n9202);
   U29726 : OAI222_X1 port map( A1 => n40894, A2 => n40391, B1 => n41278, B2 =>
                           n40384, C1 => n40380, C2 => n31701, ZN => n9201);
   U29727 : OAI222_X1 port map( A1 => n40900, A2 => n40391, B1 => n41284, B2 =>
                           n40384, C1 => n40380, C2 => n31700, ZN => n9200);
   U29728 : OAI222_X1 port map( A1 => n40906, A2 => n40391, B1 => n41290, B2 =>
                           n40384, C1 => n40380, C2 => n31699, ZN => n9199);
   U29729 : OAI222_X1 port map( A1 => n40912, A2 => n40390, B1 => n41296, B2 =>
                           n40383, C1 => n40380, C2 => n31698, ZN => n9198);
   U29730 : OAI222_X1 port map( A1 => n40918, A2 => n40390, B1 => n41302, B2 =>
                           n40383, C1 => n40380, C2 => n31697, ZN => n9197);
   U29731 : OAI222_X1 port map( A1 => n40924, A2 => n40390, B1 => n41308, B2 =>
                           n40383, C1 => n40380, C2 => n31696, ZN => n9196);
   U29732 : OAI222_X1 port map( A1 => n40930, A2 => n40390, B1 => n41314, B2 =>
                           n40383, C1 => n40380, C2 => n31695, ZN => n9195);
   U29733 : OAI222_X1 port map( A1 => n40936, A2 => n40390, B1 => n41320, B2 =>
                           n40383, C1 => n40380, C2 => n31694, ZN => n9194);
   U29734 : OAI222_X1 port map( A1 => n40942, A2 => n40390, B1 => n41326, B2 =>
                           n40383, C1 => n40380, C2 => n31693, ZN => n9193);
   U29735 : OAI222_X1 port map( A1 => n40948, A2 => n40390, B1 => n41332, B2 =>
                           n40383, C1 => n40380, C2 => n31692, ZN => n9192);
   U29736 : OAI222_X1 port map( A1 => n40960, A2 => n40390, B1 => n41344, B2 =>
                           n40383, C1 => n40380, C2 => n31690, ZN => n9190);
   U29737 : OAI222_X1 port map( A1 => n40600, A2 => n40375, B1 => n40984, B2 =>
                           n40368, C1 => n40356, C2 => n31686, ZN => n9186);
   U29738 : OAI222_X1 port map( A1 => n40606, A2 => n40375, B1 => n40990, B2 =>
                           n40368, C1 => n40356, C2 => n31685, ZN => n9185);
   U29739 : OAI222_X1 port map( A1 => n40612, A2 => n40375, B1 => n40996, B2 =>
                           n40368, C1 => n40356, C2 => n31684, ZN => n9184);
   U29740 : OAI222_X1 port map( A1 => n40618, A2 => n40375, B1 => n41002, B2 =>
                           n40368, C1 => n40356, C2 => n31683, ZN => n9183);
   U29741 : OAI222_X1 port map( A1 => n40624, A2 => n40374, B1 => n41008, B2 =>
                           n40367, C1 => n40356, C2 => n31682, ZN => n9182);
   U29742 : OAI222_X1 port map( A1 => n40630, A2 => n40374, B1 => n41014, B2 =>
                           n40367, C1 => n40356, C2 => n31681, ZN => n9181);
   U29743 : OAI222_X1 port map( A1 => n40636, A2 => n40374, B1 => n41020, B2 =>
                           n40367, C1 => n40356, C2 => n31680, ZN => n9180);
   U29744 : OAI222_X1 port map( A1 => n40642, A2 => n40374, B1 => n41026, B2 =>
                           n40367, C1 => n40356, C2 => n31679, ZN => n9179);
   U29745 : OAI222_X1 port map( A1 => n40648, A2 => n40374, B1 => n41032, B2 =>
                           n40367, C1 => n40356, C2 => n31678, ZN => n9178);
   U29746 : OAI222_X1 port map( A1 => n40654, A2 => n40374, B1 => n41038, B2 =>
                           n40367, C1 => n40356, C2 => n31677, ZN => n9177);
   U29747 : OAI222_X1 port map( A1 => n40660, A2 => n40374, B1 => n41044, B2 =>
                           n40367, C1 => n40356, C2 => n31676, ZN => n9176);
   U29748 : OAI222_X1 port map( A1 => n40666, A2 => n40374, B1 => n41050, B2 =>
                           n40367, C1 => n40356, C2 => n31675, ZN => n9175);
   U29749 : OAI222_X1 port map( A1 => n40672, A2 => n40374, B1 => n41056, B2 =>
                           n40367, C1 => n40357, C2 => n31674, ZN => n9174);
   U29750 : OAI222_X1 port map( A1 => n40678, A2 => n40374, B1 => n41062, B2 =>
                           n40367, C1 => n40357, C2 => n31673, ZN => n9173);
   U29751 : OAI222_X1 port map( A1 => n40684, A2 => n40374, B1 => n41068, B2 =>
                           n40367, C1 => n40357, C2 => n31672, ZN => n9172);
   U29752 : OAI222_X1 port map( A1 => n40690, A2 => n40374, B1 => n41074, B2 =>
                           n40367, C1 => n40358, C2 => n31671, ZN => n9171);
   U29753 : OAI222_X1 port map( A1 => n40696, A2 => n40373, B1 => n41080, B2 =>
                           n40366, C1 => n40357, C2 => n31670, ZN => n9170);
   U29754 : OAI222_X1 port map( A1 => n40702, A2 => n40373, B1 => n41086, B2 =>
                           n40366, C1 => n40357, C2 => n31669, ZN => n9169);
   U29755 : OAI222_X1 port map( A1 => n40708, A2 => n40373, B1 => n41092, B2 =>
                           n40366, C1 => n40357, C2 => n31668, ZN => n9168);
   U29756 : OAI222_X1 port map( A1 => n40714, A2 => n40373, B1 => n41098, B2 =>
                           n40366, C1 => n40357, C2 => n31667, ZN => n9167);
   U29757 : OAI222_X1 port map( A1 => n40720, A2 => n40373, B1 => n41104, B2 =>
                           n40366, C1 => n40357, C2 => n31666, ZN => n9166);
   U29758 : OAI222_X1 port map( A1 => n40726, A2 => n40373, B1 => n41110, B2 =>
                           n40366, C1 => n40357, C2 => n31665, ZN => n9165);
   U29759 : OAI222_X1 port map( A1 => n40732, A2 => n40373, B1 => n41116, B2 =>
                           n40366, C1 => n40357, C2 => n31664, ZN => n9164);
   U29760 : OAI222_X1 port map( A1 => n40738, A2 => n40373, B1 => n41122, B2 =>
                           n40366, C1 => n40357, C2 => n31663, ZN => n9163);
   U29761 : OAI222_X1 port map( A1 => n40744, A2 => n40373, B1 => n41128, B2 =>
                           n40366, C1 => n40357, C2 => n31662, ZN => n9162);
   U29762 : OAI222_X1 port map( A1 => n40750, A2 => n40373, B1 => n41134, B2 =>
                           n40366, C1 => n40358, C2 => n31661, ZN => n9161);
   U29763 : OAI222_X1 port map( A1 => n40756, A2 => n40373, B1 => n41140, B2 =>
                           n40366, C1 => n40358, C2 => n31660, ZN => n9160);
   U29764 : OAI222_X1 port map( A1 => n40762, A2 => n40373, B1 => n41146, B2 =>
                           n40366, C1 => n40358, C2 => n31659, ZN => n9159);
   U29765 : OAI222_X1 port map( A1 => n40768, A2 => n40372, B1 => n41152, B2 =>
                           n40365, C1 => n40358, C2 => n31658, ZN => n9158);
   U29766 : OAI222_X1 port map( A1 => n40774, A2 => n40372, B1 => n41158, B2 =>
                           n40365, C1 => n40358, C2 => n31657, ZN => n9157);
   U29767 : OAI222_X1 port map( A1 => n40780, A2 => n40372, B1 => n41164, B2 =>
                           n40365, C1 => n40358, C2 => n31656, ZN => n9156);
   U29768 : OAI222_X1 port map( A1 => n40786, A2 => n40372, B1 => n41170, B2 =>
                           n40365, C1 => n40358, C2 => n31655, ZN => n9155);
   U29769 : OAI222_X1 port map( A1 => n40792, A2 => n40372, B1 => n41176, B2 =>
                           n40365, C1 => n40358, C2 => n31654, ZN => n9154);
   U29770 : OAI222_X1 port map( A1 => n40798, A2 => n40372, B1 => n41182, B2 =>
                           n40365, C1 => n40358, C2 => n31653, ZN => n9153);
   U29771 : OAI222_X1 port map( A1 => n40804, A2 => n40372, B1 => n41188, B2 =>
                           n40365, C1 => n40358, C2 => n31652, ZN => n9152);
   U29772 : OAI222_X1 port map( A1 => n40810, A2 => n40372, B1 => n41194, B2 =>
                           n40365, C1 => n40358, C2 => n31651, ZN => n9151);
   U29773 : OAI222_X1 port map( A1 => n40816, A2 => n40372, B1 => n41200, B2 =>
                           n40365, C1 => n40359, C2 => n31650, ZN => n9150);
   U29774 : OAI222_X1 port map( A1 => n40822, A2 => n40372, B1 => n41206, B2 =>
                           n40365, C1 => n40359, C2 => n31649, ZN => n9149);
   U29775 : OAI222_X1 port map( A1 => n40828, A2 => n40372, B1 => n41212, B2 =>
                           n40365, C1 => n40359, C2 => n31648, ZN => n9148);
   U29776 : OAI222_X1 port map( A1 => n40834, A2 => n40372, B1 => n41218, B2 =>
                           n40365, C1 => n40359, C2 => n31647, ZN => n9147);
   U29777 : OAI222_X1 port map( A1 => n40840, A2 => n40371, B1 => n41224, B2 =>
                           n40364, C1 => n40359, C2 => n31646, ZN => n9146);
   U29778 : OAI222_X1 port map( A1 => n40846, A2 => n40371, B1 => n41230, B2 =>
                           n40364, C1 => n40359, C2 => n31645, ZN => n9145);
   U29779 : OAI222_X1 port map( A1 => n40852, A2 => n40371, B1 => n41236, B2 =>
                           n40364, C1 => n40359, C2 => n31644, ZN => n9144);
   U29780 : OAI222_X1 port map( A1 => n40858, A2 => n40371, B1 => n41242, B2 =>
                           n40364, C1 => n40359, C2 => n31643, ZN => n9143);
   U29781 : OAI222_X1 port map( A1 => n40864, A2 => n40371, B1 => n41248, B2 =>
                           n40364, C1 => n40359, C2 => n31642, ZN => n9142);
   U29782 : OAI222_X1 port map( A1 => n40870, A2 => n40371, B1 => n41254, B2 =>
                           n40364, C1 => n40359, C2 => n31641, ZN => n9141);
   U29783 : OAI222_X1 port map( A1 => n40876, A2 => n40371, B1 => n41260, B2 =>
                           n40364, C1 => n40359, C2 => n31640, ZN => n9140);
   U29784 : OAI222_X1 port map( A1 => n40882, A2 => n40371, B1 => n41266, B2 =>
                           n40364, C1 => n40359, C2 => n31639, ZN => n9139);
   U29785 : OAI222_X1 port map( A1 => n40888, A2 => n40371, B1 => n41272, B2 =>
                           n40364, C1 => n40360, C2 => n31638, ZN => n9138);
   U29786 : OAI222_X1 port map( A1 => n40894, A2 => n40371, B1 => n41278, B2 =>
                           n40364, C1 => n40360, C2 => n31637, ZN => n9137);
   U29787 : OAI222_X1 port map( A1 => n40900, A2 => n40371, B1 => n41284, B2 =>
                           n40364, C1 => n40360, C2 => n31636, ZN => n9136);
   U29788 : OAI222_X1 port map( A1 => n40906, A2 => n40371, B1 => n41290, B2 =>
                           n40364, C1 => n40360, C2 => n31635, ZN => n9135);
   U29789 : OAI222_X1 port map( A1 => n40912, A2 => n40370, B1 => n41296, B2 =>
                           n40363, C1 => n40360, C2 => n31634, ZN => n9134);
   U29790 : OAI222_X1 port map( A1 => n40918, A2 => n40370, B1 => n41302, B2 =>
                           n40363, C1 => n40360, C2 => n31633, ZN => n9133);
   U29791 : OAI222_X1 port map( A1 => n40924, A2 => n40370, B1 => n41308, B2 =>
                           n40363, C1 => n40360, C2 => n31632, ZN => n9132);
   U29792 : OAI222_X1 port map( A1 => n40930, A2 => n40370, B1 => n41314, B2 =>
                           n40363, C1 => n40360, C2 => n31631, ZN => n9131);
   U29793 : OAI222_X1 port map( A1 => n40936, A2 => n40370, B1 => n41320, B2 =>
                           n40363, C1 => n40360, C2 => n31630, ZN => n9130);
   U29794 : OAI222_X1 port map( A1 => n40942, A2 => n40370, B1 => n41326, B2 =>
                           n40363, C1 => n40360, C2 => n31629, ZN => n9129);
   U29795 : OAI222_X1 port map( A1 => n40948, A2 => n40370, B1 => n41332, B2 =>
                           n40363, C1 => n40360, C2 => n31628, ZN => n9128);
   U29796 : OAI222_X1 port map( A1 => n40960, A2 => n40370, B1 => n41344, B2 =>
                           n40363, C1 => n40360, C2 => n31626, ZN => n9126);
   U29797 : OAI222_X1 port map( A1 => n40600, A2 => n40355, B1 => n40984, B2 =>
                           n40348, C1 => n40336, C2 => n31622, ZN => n9122);
   U29798 : OAI222_X1 port map( A1 => n40606, A2 => n40355, B1 => n40990, B2 =>
                           n40348, C1 => n40336, C2 => n31621, ZN => n9121);
   U29799 : OAI222_X1 port map( A1 => n40612, A2 => n40355, B1 => n40996, B2 =>
                           n40348, C1 => n40336, C2 => n31620, ZN => n9120);
   U29800 : OAI222_X1 port map( A1 => n40618, A2 => n40355, B1 => n41002, B2 =>
                           n40348, C1 => n40336, C2 => n31619, ZN => n9119);
   U29801 : OAI222_X1 port map( A1 => n40624, A2 => n40354, B1 => n41008, B2 =>
                           n40347, C1 => n40336, C2 => n31618, ZN => n9118);
   U29802 : OAI222_X1 port map( A1 => n40630, A2 => n40354, B1 => n41014, B2 =>
                           n40347, C1 => n40336, C2 => n31617, ZN => n9117);
   U29803 : OAI222_X1 port map( A1 => n40636, A2 => n40354, B1 => n41020, B2 =>
                           n40347, C1 => n40336, C2 => n31616, ZN => n9116);
   U29804 : OAI222_X1 port map( A1 => n40642, A2 => n40354, B1 => n41026, B2 =>
                           n40347, C1 => n40336, C2 => n31615, ZN => n9115);
   U29805 : OAI222_X1 port map( A1 => n40648, A2 => n40354, B1 => n41032, B2 =>
                           n40347, C1 => n40336, C2 => n31614, ZN => n9114);
   U29806 : OAI222_X1 port map( A1 => n40654, A2 => n40354, B1 => n41038, B2 =>
                           n40347, C1 => n40336, C2 => n31613, ZN => n9113);
   U29807 : OAI222_X1 port map( A1 => n40660, A2 => n40354, B1 => n41044, B2 =>
                           n40347, C1 => n40336, C2 => n31612, ZN => n9112);
   U29808 : OAI222_X1 port map( A1 => n40666, A2 => n40354, B1 => n41050, B2 =>
                           n40347, C1 => n40336, C2 => n31611, ZN => n9111);
   U29809 : OAI222_X1 port map( A1 => n40672, A2 => n40354, B1 => n41056, B2 =>
                           n40347, C1 => n40337, C2 => n31610, ZN => n9110);
   U29810 : OAI222_X1 port map( A1 => n40678, A2 => n40354, B1 => n41062, B2 =>
                           n40347, C1 => n40337, C2 => n31609, ZN => n9109);
   U29811 : OAI222_X1 port map( A1 => n40684, A2 => n40354, B1 => n41068, B2 =>
                           n40347, C1 => n40337, C2 => n31608, ZN => n9108);
   U29812 : OAI222_X1 port map( A1 => n40690, A2 => n40354, B1 => n41074, B2 =>
                           n40347, C1 => n40338, C2 => n31607, ZN => n9107);
   U29813 : OAI222_X1 port map( A1 => n40696, A2 => n40353, B1 => n41080, B2 =>
                           n40346, C1 => n40337, C2 => n31606, ZN => n9106);
   U29814 : OAI222_X1 port map( A1 => n40702, A2 => n40353, B1 => n41086, B2 =>
                           n40346, C1 => n40337, C2 => n31605, ZN => n9105);
   U29815 : OAI222_X1 port map( A1 => n40708, A2 => n40353, B1 => n41092, B2 =>
                           n40346, C1 => n40337, C2 => n31604, ZN => n9104);
   U29816 : OAI222_X1 port map( A1 => n40714, A2 => n40353, B1 => n41098, B2 =>
                           n40346, C1 => n40337, C2 => n31603, ZN => n9103);
   U29817 : OAI222_X1 port map( A1 => n40720, A2 => n40353, B1 => n41104, B2 =>
                           n40346, C1 => n40337, C2 => n31602, ZN => n9102);
   U29818 : OAI222_X1 port map( A1 => n40726, A2 => n40353, B1 => n41110, B2 =>
                           n40346, C1 => n40337, C2 => n31601, ZN => n9101);
   U29819 : OAI222_X1 port map( A1 => n40732, A2 => n40353, B1 => n41116, B2 =>
                           n40346, C1 => n40337, C2 => n31600, ZN => n9100);
   U29820 : OAI222_X1 port map( A1 => n40738, A2 => n40353, B1 => n41122, B2 =>
                           n40346, C1 => n40337, C2 => n31599, ZN => n9099);
   U29821 : OAI222_X1 port map( A1 => n40744, A2 => n40353, B1 => n41128, B2 =>
                           n40346, C1 => n40337, C2 => n31598, ZN => n9098);
   U29822 : OAI222_X1 port map( A1 => n40750, A2 => n40353, B1 => n41134, B2 =>
                           n40346, C1 => n40338, C2 => n31597, ZN => n9097);
   U29823 : OAI222_X1 port map( A1 => n40756, A2 => n40353, B1 => n41140, B2 =>
                           n40346, C1 => n40338, C2 => n31596, ZN => n9096);
   U29824 : OAI222_X1 port map( A1 => n40762, A2 => n40353, B1 => n41146, B2 =>
                           n40346, C1 => n40338, C2 => n31595, ZN => n9095);
   U29825 : OAI222_X1 port map( A1 => n40768, A2 => n40352, B1 => n41152, B2 =>
                           n40345, C1 => n40338, C2 => n31594, ZN => n9094);
   U29826 : OAI222_X1 port map( A1 => n40774, A2 => n40352, B1 => n41158, B2 =>
                           n40345, C1 => n40338, C2 => n31593, ZN => n9093);
   U29827 : OAI222_X1 port map( A1 => n40780, A2 => n40352, B1 => n41164, B2 =>
                           n40345, C1 => n40338, C2 => n31592, ZN => n9092);
   U29828 : OAI222_X1 port map( A1 => n40786, A2 => n40352, B1 => n41170, B2 =>
                           n40345, C1 => n40338, C2 => n31591, ZN => n9091);
   U29829 : OAI222_X1 port map( A1 => n40792, A2 => n40352, B1 => n41176, B2 =>
                           n40345, C1 => n40338, C2 => n31590, ZN => n9090);
   U29830 : OAI222_X1 port map( A1 => n40798, A2 => n40352, B1 => n41182, B2 =>
                           n40345, C1 => n40338, C2 => n31589, ZN => n9089);
   U29831 : OAI222_X1 port map( A1 => n40804, A2 => n40352, B1 => n41188, B2 =>
                           n40345, C1 => n40338, C2 => n31588, ZN => n9088);
   U29832 : OAI222_X1 port map( A1 => n40810, A2 => n40352, B1 => n41194, B2 =>
                           n40345, C1 => n40338, C2 => n31587, ZN => n9087);
   U29833 : OAI222_X1 port map( A1 => n40816, A2 => n40352, B1 => n41200, B2 =>
                           n40345, C1 => n40339, C2 => n31586, ZN => n9086);
   U29834 : OAI222_X1 port map( A1 => n40822, A2 => n40352, B1 => n41206, B2 =>
                           n40345, C1 => n40339, C2 => n31585, ZN => n9085);
   U29835 : OAI222_X1 port map( A1 => n40828, A2 => n40352, B1 => n41212, B2 =>
                           n40345, C1 => n40339, C2 => n31584, ZN => n9084);
   U29836 : OAI222_X1 port map( A1 => n40834, A2 => n40352, B1 => n41218, B2 =>
                           n40345, C1 => n40339, C2 => n31583, ZN => n9083);
   U29837 : OAI222_X1 port map( A1 => n40840, A2 => n40351, B1 => n41224, B2 =>
                           n40344, C1 => n40339, C2 => n31582, ZN => n9082);
   U29838 : OAI222_X1 port map( A1 => n40846, A2 => n40351, B1 => n41230, B2 =>
                           n40344, C1 => n40339, C2 => n31581, ZN => n9081);
   U29839 : OAI222_X1 port map( A1 => n40852, A2 => n40351, B1 => n41236, B2 =>
                           n40344, C1 => n40339, C2 => n31580, ZN => n9080);
   U29840 : OAI222_X1 port map( A1 => n40858, A2 => n40351, B1 => n41242, B2 =>
                           n40344, C1 => n40339, C2 => n31579, ZN => n9079);
   U29841 : OAI222_X1 port map( A1 => n40864, A2 => n40351, B1 => n41248, B2 =>
                           n40344, C1 => n40339, C2 => n31578, ZN => n9078);
   U29842 : OAI222_X1 port map( A1 => n40870, A2 => n40351, B1 => n41254, B2 =>
                           n40344, C1 => n40339, C2 => n31577, ZN => n9077);
   U29843 : OAI222_X1 port map( A1 => n40876, A2 => n40351, B1 => n41260, B2 =>
                           n40344, C1 => n40339, C2 => n31576, ZN => n9076);
   U29844 : OAI222_X1 port map( A1 => n40882, A2 => n40351, B1 => n41266, B2 =>
                           n40344, C1 => n40339, C2 => n31575, ZN => n9075);
   U29845 : OAI222_X1 port map( A1 => n40888, A2 => n40351, B1 => n41272, B2 =>
                           n40344, C1 => n40340, C2 => n31574, ZN => n9074);
   U29846 : OAI222_X1 port map( A1 => n40894, A2 => n40351, B1 => n41278, B2 =>
                           n40344, C1 => n40340, C2 => n31573, ZN => n9073);
   U29847 : OAI222_X1 port map( A1 => n40900, A2 => n40351, B1 => n41284, B2 =>
                           n40344, C1 => n40340, C2 => n31572, ZN => n9072);
   U29848 : OAI222_X1 port map( A1 => n40906, A2 => n40351, B1 => n41290, B2 =>
                           n40344, C1 => n40340, C2 => n31571, ZN => n9071);
   U29849 : OAI222_X1 port map( A1 => n40912, A2 => n40350, B1 => n41296, B2 =>
                           n40343, C1 => n40340, C2 => n31570, ZN => n9070);
   U29850 : OAI222_X1 port map( A1 => n40918, A2 => n40350, B1 => n41302, B2 =>
                           n40343, C1 => n40340, C2 => n31569, ZN => n9069);
   U29851 : OAI222_X1 port map( A1 => n40924, A2 => n40350, B1 => n41308, B2 =>
                           n40343, C1 => n40340, C2 => n31568, ZN => n9068);
   U29852 : OAI222_X1 port map( A1 => n40930, A2 => n40350, B1 => n41314, B2 =>
                           n40343, C1 => n40340, C2 => n31567, ZN => n9067);
   U29853 : OAI222_X1 port map( A1 => n40936, A2 => n40350, B1 => n41320, B2 =>
                           n40343, C1 => n40340, C2 => n31566, ZN => n9066);
   U29854 : OAI222_X1 port map( A1 => n40942, A2 => n40350, B1 => n41326, B2 =>
                           n40343, C1 => n40340, C2 => n31565, ZN => n9065);
   U29855 : OAI222_X1 port map( A1 => n40948, A2 => n40350, B1 => n41332, B2 =>
                           n40343, C1 => n40340, C2 => n31564, ZN => n9064);
   U29856 : OAI222_X1 port map( A1 => n40960, A2 => n40350, B1 => n41344, B2 =>
                           n40343, C1 => n40340, C2 => n31562, ZN => n9062);
   U29857 : OAI222_X1 port map( A1 => n40600, A2 => n40295, B1 => n40984, B2 =>
                           n40288, C1 => n40276, C2 => n31558, ZN => n8930);
   U29858 : OAI222_X1 port map( A1 => n40606, A2 => n40295, B1 => n40990, B2 =>
                           n40288, C1 => n40276, C2 => n31557, ZN => n8929);
   U29859 : OAI222_X1 port map( A1 => n40612, A2 => n40295, B1 => n40996, B2 =>
                           n40288, C1 => n40276, C2 => n31556, ZN => n8928);
   U29860 : OAI222_X1 port map( A1 => n40618, A2 => n40295, B1 => n41002, B2 =>
                           n40288, C1 => n40276, C2 => n31555, ZN => n8927);
   U29861 : OAI222_X1 port map( A1 => n40624, A2 => n40294, B1 => n41008, B2 =>
                           n40287, C1 => n40276, C2 => n31554, ZN => n8926);
   U29862 : OAI222_X1 port map( A1 => n40630, A2 => n40294, B1 => n41014, B2 =>
                           n40287, C1 => n40276, C2 => n31553, ZN => n8925);
   U29863 : OAI222_X1 port map( A1 => n40636, A2 => n40294, B1 => n41020, B2 =>
                           n40287, C1 => n40276, C2 => n31552, ZN => n8924);
   U29864 : OAI222_X1 port map( A1 => n40642, A2 => n40294, B1 => n41026, B2 =>
                           n40287, C1 => n40276, C2 => n31551, ZN => n8923);
   U29865 : OAI222_X1 port map( A1 => n40648, A2 => n40294, B1 => n41032, B2 =>
                           n40287, C1 => n40276, C2 => n31550, ZN => n8922);
   U29866 : OAI222_X1 port map( A1 => n40654, A2 => n40294, B1 => n41038, B2 =>
                           n40287, C1 => n40276, C2 => n31549, ZN => n8921);
   U29867 : OAI222_X1 port map( A1 => n40660, A2 => n40294, B1 => n41044, B2 =>
                           n40287, C1 => n40276, C2 => n31548, ZN => n8920);
   U29868 : OAI222_X1 port map( A1 => n40666, A2 => n40294, B1 => n41050, B2 =>
                           n40287, C1 => n40276, C2 => n31547, ZN => n8919);
   U29869 : OAI222_X1 port map( A1 => n40672, A2 => n40294, B1 => n41056, B2 =>
                           n40287, C1 => n40277, C2 => n31546, ZN => n8918);
   U29870 : OAI222_X1 port map( A1 => n40678, A2 => n40294, B1 => n41062, B2 =>
                           n40287, C1 => n40277, C2 => n31545, ZN => n8917);
   U29871 : OAI222_X1 port map( A1 => n40684, A2 => n40294, B1 => n41068, B2 =>
                           n40287, C1 => n40277, C2 => n31544, ZN => n8916);
   U29872 : OAI222_X1 port map( A1 => n40690, A2 => n40294, B1 => n41074, B2 =>
                           n40287, C1 => n40278, C2 => n31543, ZN => n8915);
   U29873 : OAI222_X1 port map( A1 => n40696, A2 => n40293, B1 => n41080, B2 =>
                           n40286, C1 => n40277, C2 => n31542, ZN => n8914);
   U29874 : OAI222_X1 port map( A1 => n40702, A2 => n40293, B1 => n41086, B2 =>
                           n40286, C1 => n40277, C2 => n31541, ZN => n8913);
   U29875 : OAI222_X1 port map( A1 => n40708, A2 => n40293, B1 => n41092, B2 =>
                           n40286, C1 => n40277, C2 => n31540, ZN => n8912);
   U29876 : OAI222_X1 port map( A1 => n40714, A2 => n40293, B1 => n41098, B2 =>
                           n40286, C1 => n40277, C2 => n31539, ZN => n8911);
   U29877 : OAI222_X1 port map( A1 => n40720, A2 => n40293, B1 => n41104, B2 =>
                           n40286, C1 => n40277, C2 => n31538, ZN => n8910);
   U29878 : OAI222_X1 port map( A1 => n40726, A2 => n40293, B1 => n41110, B2 =>
                           n40286, C1 => n40277, C2 => n31537, ZN => n8909);
   U29879 : OAI222_X1 port map( A1 => n40732, A2 => n40293, B1 => n41116, B2 =>
                           n40286, C1 => n40277, C2 => n31536, ZN => n8908);
   U29880 : OAI222_X1 port map( A1 => n40738, A2 => n40293, B1 => n41122, B2 =>
                           n40286, C1 => n40277, C2 => n31535, ZN => n8907);
   U29881 : OAI222_X1 port map( A1 => n40744, A2 => n40293, B1 => n41128, B2 =>
                           n40286, C1 => n40277, C2 => n31534, ZN => n8906);
   U29882 : OAI222_X1 port map( A1 => n40750, A2 => n40293, B1 => n41134, B2 =>
                           n40286, C1 => n40278, C2 => n31533, ZN => n8905);
   U29883 : OAI222_X1 port map( A1 => n40756, A2 => n40293, B1 => n41140, B2 =>
                           n40286, C1 => n40278, C2 => n31532, ZN => n8904);
   U29884 : OAI222_X1 port map( A1 => n40762, A2 => n40293, B1 => n41146, B2 =>
                           n40286, C1 => n40278, C2 => n31531, ZN => n8903);
   U29885 : OAI222_X1 port map( A1 => n40768, A2 => n40292, B1 => n41152, B2 =>
                           n40285, C1 => n40278, C2 => n31530, ZN => n8902);
   U29886 : OAI222_X1 port map( A1 => n40774, A2 => n40292, B1 => n41158, B2 =>
                           n40285, C1 => n40278, C2 => n31529, ZN => n8901);
   U29887 : OAI222_X1 port map( A1 => n40780, A2 => n40292, B1 => n41164, B2 =>
                           n40285, C1 => n40278, C2 => n31528, ZN => n8900);
   U29888 : OAI222_X1 port map( A1 => n40786, A2 => n40292, B1 => n41170, B2 =>
                           n40285, C1 => n40278, C2 => n31527, ZN => n8899);
   U29889 : OAI222_X1 port map( A1 => n40792, A2 => n40292, B1 => n41176, B2 =>
                           n40285, C1 => n40278, C2 => n31526, ZN => n8898);
   U29890 : OAI222_X1 port map( A1 => n40798, A2 => n40292, B1 => n41182, B2 =>
                           n40285, C1 => n40278, C2 => n31525, ZN => n8897);
   U29891 : OAI222_X1 port map( A1 => n40804, A2 => n40292, B1 => n41188, B2 =>
                           n40285, C1 => n40278, C2 => n31524, ZN => n8896);
   U29892 : OAI222_X1 port map( A1 => n40810, A2 => n40292, B1 => n41194, B2 =>
                           n40285, C1 => n40278, C2 => n31523, ZN => n8895);
   U29893 : OAI222_X1 port map( A1 => n40816, A2 => n40292, B1 => n41200, B2 =>
                           n40285, C1 => n40279, C2 => n31522, ZN => n8894);
   U29894 : OAI222_X1 port map( A1 => n40822, A2 => n40292, B1 => n41206, B2 =>
                           n40285, C1 => n40279, C2 => n31521, ZN => n8893);
   U29895 : OAI222_X1 port map( A1 => n40828, A2 => n40292, B1 => n41212, B2 =>
                           n40285, C1 => n40279, C2 => n31520, ZN => n8892);
   U29896 : OAI222_X1 port map( A1 => n40834, A2 => n40292, B1 => n41218, B2 =>
                           n40285, C1 => n40279, C2 => n31519, ZN => n8891);
   U29897 : OAI222_X1 port map( A1 => n40840, A2 => n40291, B1 => n41224, B2 =>
                           n40284, C1 => n40279, C2 => n31518, ZN => n8890);
   U29898 : OAI222_X1 port map( A1 => n40846, A2 => n40291, B1 => n41230, B2 =>
                           n40284, C1 => n40279, C2 => n31517, ZN => n8889);
   U29899 : OAI222_X1 port map( A1 => n40852, A2 => n40291, B1 => n41236, B2 =>
                           n40284, C1 => n40279, C2 => n31516, ZN => n8888);
   U29900 : OAI222_X1 port map( A1 => n40858, A2 => n40291, B1 => n41242, B2 =>
                           n40284, C1 => n40279, C2 => n31515, ZN => n8887);
   U29901 : OAI222_X1 port map( A1 => n40864, A2 => n40291, B1 => n41248, B2 =>
                           n40284, C1 => n40279, C2 => n31514, ZN => n8886);
   U29902 : OAI222_X1 port map( A1 => n40870, A2 => n40291, B1 => n41254, B2 =>
                           n40284, C1 => n40279, C2 => n31513, ZN => n8885);
   U29903 : OAI222_X1 port map( A1 => n40876, A2 => n40291, B1 => n41260, B2 =>
                           n40284, C1 => n40279, C2 => n31512, ZN => n8884);
   U29904 : OAI222_X1 port map( A1 => n40882, A2 => n40291, B1 => n41266, B2 =>
                           n40284, C1 => n40279, C2 => n31511, ZN => n8883);
   U29905 : OAI222_X1 port map( A1 => n40888, A2 => n40291, B1 => n41272, B2 =>
                           n40284, C1 => n40280, C2 => n31510, ZN => n8882);
   U29906 : OAI222_X1 port map( A1 => n40894, A2 => n40291, B1 => n41278, B2 =>
                           n40284, C1 => n40280, C2 => n31509, ZN => n8881);
   U29907 : OAI222_X1 port map( A1 => n40900, A2 => n40291, B1 => n41284, B2 =>
                           n40284, C1 => n40280, C2 => n31508, ZN => n8880);
   U29908 : OAI222_X1 port map( A1 => n40906, A2 => n40291, B1 => n41290, B2 =>
                           n40284, C1 => n40280, C2 => n31507, ZN => n8879);
   U29909 : OAI222_X1 port map( A1 => n40912, A2 => n40290, B1 => n41296, B2 =>
                           n40283, C1 => n40280, C2 => n31506, ZN => n8878);
   U29910 : OAI222_X1 port map( A1 => n40918, A2 => n40290, B1 => n41302, B2 =>
                           n40283, C1 => n40280, C2 => n31505, ZN => n8877);
   U29911 : OAI222_X1 port map( A1 => n40924, A2 => n40290, B1 => n41308, B2 =>
                           n40283, C1 => n40280, C2 => n31504, ZN => n8876);
   U29912 : OAI222_X1 port map( A1 => n40930, A2 => n40290, B1 => n41314, B2 =>
                           n40283, C1 => n40280, C2 => n31503, ZN => n8875);
   U29913 : OAI222_X1 port map( A1 => n40936, A2 => n40290, B1 => n41320, B2 =>
                           n40283, C1 => n40280, C2 => n31502, ZN => n8874);
   U29914 : OAI222_X1 port map( A1 => n40942, A2 => n40290, B1 => n41326, B2 =>
                           n40283, C1 => n40280, C2 => n31501, ZN => n8873);
   U29915 : OAI222_X1 port map( A1 => n40948, A2 => n40290, B1 => n41332, B2 =>
                           n40283, C1 => n40280, C2 => n31500, ZN => n8872);
   U29916 : OAI222_X1 port map( A1 => n40960, A2 => n40290, B1 => n41344, B2 =>
                           n40283, C1 => n40280, C2 => n31498, ZN => n8870);
   U29917 : OAI222_X1 port map( A1 => n40599, A2 => n40275, B1 => n40983, B2 =>
                           n40268, C1 => n40256, C2 => n31494, ZN => n8866);
   U29918 : OAI222_X1 port map( A1 => n40605, A2 => n40275, B1 => n40989, B2 =>
                           n40268, C1 => n40256, C2 => n31493, ZN => n8865);
   U29919 : OAI222_X1 port map( A1 => n40611, A2 => n40275, B1 => n40995, B2 =>
                           n40268, C1 => n40256, C2 => n31492, ZN => n8864);
   U29920 : OAI222_X1 port map( A1 => n40617, A2 => n40275, B1 => n41001, B2 =>
                           n40268, C1 => n40256, C2 => n31491, ZN => n8863);
   U29921 : OAI222_X1 port map( A1 => n40623, A2 => n40274, B1 => n41007, B2 =>
                           n40267, C1 => n40256, C2 => n31490, ZN => n8862);
   U29922 : OAI222_X1 port map( A1 => n40629, A2 => n40274, B1 => n41013, B2 =>
                           n40267, C1 => n40256, C2 => n31489, ZN => n8861);
   U29923 : OAI222_X1 port map( A1 => n40635, A2 => n40274, B1 => n41019, B2 =>
                           n40267, C1 => n40256, C2 => n31488, ZN => n8860);
   U29924 : OAI222_X1 port map( A1 => n40641, A2 => n40274, B1 => n41025, B2 =>
                           n40267, C1 => n40256, C2 => n31487, ZN => n8859);
   U29925 : OAI222_X1 port map( A1 => n40647, A2 => n40274, B1 => n41031, B2 =>
                           n40267, C1 => n40256, C2 => n31486, ZN => n8858);
   U29926 : OAI222_X1 port map( A1 => n40653, A2 => n40274, B1 => n41037, B2 =>
                           n40267, C1 => n40256, C2 => n31485, ZN => n8857);
   U29927 : OAI222_X1 port map( A1 => n40659, A2 => n40274, B1 => n41043, B2 =>
                           n40267, C1 => n40256, C2 => n31484, ZN => n8856);
   U29928 : OAI222_X1 port map( A1 => n40665, A2 => n40274, B1 => n41049, B2 =>
                           n40267, C1 => n40256, C2 => n31483, ZN => n8855);
   U29929 : OAI222_X1 port map( A1 => n40671, A2 => n40274, B1 => n41055, B2 =>
                           n40267, C1 => n40257, C2 => n31482, ZN => n8854);
   U29930 : OAI222_X1 port map( A1 => n40677, A2 => n40274, B1 => n41061, B2 =>
                           n40267, C1 => n40257, C2 => n31481, ZN => n8853);
   U29931 : OAI222_X1 port map( A1 => n40683, A2 => n40274, B1 => n41067, B2 =>
                           n40267, C1 => n40257, C2 => n31480, ZN => n8852);
   U29932 : OAI222_X1 port map( A1 => n40689, A2 => n40274, B1 => n41073, B2 =>
                           n40267, C1 => n40258, C2 => n31479, ZN => n8851);
   U29933 : OAI222_X1 port map( A1 => n40695, A2 => n40273, B1 => n41079, B2 =>
                           n40266, C1 => n40257, C2 => n31478, ZN => n8850);
   U29934 : OAI222_X1 port map( A1 => n40701, A2 => n40273, B1 => n41085, B2 =>
                           n40266, C1 => n40257, C2 => n31477, ZN => n8849);
   U29935 : OAI222_X1 port map( A1 => n40707, A2 => n40273, B1 => n41091, B2 =>
                           n40266, C1 => n40257, C2 => n31476, ZN => n8848);
   U29936 : OAI222_X1 port map( A1 => n40713, A2 => n40273, B1 => n41097, B2 =>
                           n40266, C1 => n40257, C2 => n31475, ZN => n8847);
   U29937 : OAI222_X1 port map( A1 => n40719, A2 => n40273, B1 => n41103, B2 =>
                           n40266, C1 => n40257, C2 => n31474, ZN => n8846);
   U29938 : OAI222_X1 port map( A1 => n40725, A2 => n40273, B1 => n41109, B2 =>
                           n40266, C1 => n40257, C2 => n31473, ZN => n8845);
   U29939 : OAI222_X1 port map( A1 => n40731, A2 => n40273, B1 => n41115, B2 =>
                           n40266, C1 => n40257, C2 => n31472, ZN => n8844);
   U29940 : OAI222_X1 port map( A1 => n40737, A2 => n40273, B1 => n41121, B2 =>
                           n40266, C1 => n40257, C2 => n31471, ZN => n8843);
   U29941 : OAI222_X1 port map( A1 => n40743, A2 => n40273, B1 => n41127, B2 =>
                           n40266, C1 => n40257, C2 => n31470, ZN => n8842);
   U29942 : OAI222_X1 port map( A1 => n40749, A2 => n40273, B1 => n41133, B2 =>
                           n40266, C1 => n40258, C2 => n31469, ZN => n8841);
   U29943 : OAI222_X1 port map( A1 => n40755, A2 => n40273, B1 => n41139, B2 =>
                           n40266, C1 => n40258, C2 => n31468, ZN => n8840);
   U29944 : OAI222_X1 port map( A1 => n40761, A2 => n40273, B1 => n41145, B2 =>
                           n40266, C1 => n40258, C2 => n31467, ZN => n8839);
   U29945 : OAI222_X1 port map( A1 => n40767, A2 => n40272, B1 => n41151, B2 =>
                           n40265, C1 => n40258, C2 => n31466, ZN => n8838);
   U29946 : OAI222_X1 port map( A1 => n40773, A2 => n40272, B1 => n41157, B2 =>
                           n40265, C1 => n40258, C2 => n31465, ZN => n8837);
   U29947 : OAI222_X1 port map( A1 => n40779, A2 => n40272, B1 => n41163, B2 =>
                           n40265, C1 => n40258, C2 => n31464, ZN => n8836);
   U29948 : OAI222_X1 port map( A1 => n40785, A2 => n40272, B1 => n41169, B2 =>
                           n40265, C1 => n40258, C2 => n31463, ZN => n8835);
   U29949 : OAI222_X1 port map( A1 => n40791, A2 => n40272, B1 => n41175, B2 =>
                           n40265, C1 => n40258, C2 => n31462, ZN => n8834);
   U29950 : OAI222_X1 port map( A1 => n40797, A2 => n40272, B1 => n41181, B2 =>
                           n40265, C1 => n40258, C2 => n31461, ZN => n8833);
   U29951 : OAI222_X1 port map( A1 => n40803, A2 => n40272, B1 => n41187, B2 =>
                           n40265, C1 => n40258, C2 => n31460, ZN => n8832);
   U29952 : OAI222_X1 port map( A1 => n40809, A2 => n40272, B1 => n41193, B2 =>
                           n40265, C1 => n40258, C2 => n31459, ZN => n8831);
   U29953 : OAI222_X1 port map( A1 => n40815, A2 => n40272, B1 => n41199, B2 =>
                           n40265, C1 => n40259, C2 => n31458, ZN => n8830);
   U29954 : OAI222_X1 port map( A1 => n40821, A2 => n40272, B1 => n41205, B2 =>
                           n40265, C1 => n40259, C2 => n31457, ZN => n8829);
   U29955 : OAI222_X1 port map( A1 => n40827, A2 => n40272, B1 => n41211, B2 =>
                           n40265, C1 => n40259, C2 => n31456, ZN => n8828);
   U29956 : OAI222_X1 port map( A1 => n40833, A2 => n40272, B1 => n41217, B2 =>
                           n40265, C1 => n40259, C2 => n31455, ZN => n8827);
   U29957 : OAI222_X1 port map( A1 => n40839, A2 => n40271, B1 => n41223, B2 =>
                           n40264, C1 => n40259, C2 => n31454, ZN => n8826);
   U29958 : OAI222_X1 port map( A1 => n40845, A2 => n40271, B1 => n41229, B2 =>
                           n40264, C1 => n40259, C2 => n31453, ZN => n8825);
   U29959 : OAI222_X1 port map( A1 => n40851, A2 => n40271, B1 => n41235, B2 =>
                           n40264, C1 => n40259, C2 => n31452, ZN => n8824);
   U29960 : OAI222_X1 port map( A1 => n40857, A2 => n40271, B1 => n41241, B2 =>
                           n40264, C1 => n40259, C2 => n31451, ZN => n8823);
   U29961 : OAI222_X1 port map( A1 => n40863, A2 => n40271, B1 => n41247, B2 =>
                           n40264, C1 => n40259, C2 => n31450, ZN => n8822);
   U29962 : OAI222_X1 port map( A1 => n40869, A2 => n40271, B1 => n41253, B2 =>
                           n40264, C1 => n40259, C2 => n31449, ZN => n8821);
   U29963 : OAI222_X1 port map( A1 => n40875, A2 => n40271, B1 => n41259, B2 =>
                           n40264, C1 => n40259, C2 => n31448, ZN => n8820);
   U29964 : OAI222_X1 port map( A1 => n40881, A2 => n40271, B1 => n41265, B2 =>
                           n40264, C1 => n40259, C2 => n31447, ZN => n8819);
   U29965 : OAI222_X1 port map( A1 => n40887, A2 => n40271, B1 => n41271, B2 =>
                           n40264, C1 => n40260, C2 => n31446, ZN => n8818);
   U29966 : OAI222_X1 port map( A1 => n40893, A2 => n40271, B1 => n41277, B2 =>
                           n40264, C1 => n40260, C2 => n31445, ZN => n8817);
   U29967 : OAI222_X1 port map( A1 => n40899, A2 => n40271, B1 => n41283, B2 =>
                           n40264, C1 => n40260, C2 => n31444, ZN => n8816);
   U29968 : OAI222_X1 port map( A1 => n40905, A2 => n40271, B1 => n41289, B2 =>
                           n40264, C1 => n40260, C2 => n31443, ZN => n8815);
   U29969 : OAI222_X1 port map( A1 => n40911, A2 => n40270, B1 => n41295, B2 =>
                           n40263, C1 => n40260, C2 => n31442, ZN => n8814);
   U29970 : OAI222_X1 port map( A1 => n40917, A2 => n40270, B1 => n41301, B2 =>
                           n40263, C1 => n40260, C2 => n31441, ZN => n8813);
   U29971 : OAI222_X1 port map( A1 => n40923, A2 => n40270, B1 => n41307, B2 =>
                           n40263, C1 => n40260, C2 => n31440, ZN => n8812);
   U29972 : OAI222_X1 port map( A1 => n40929, A2 => n40270, B1 => n41313, B2 =>
                           n40263, C1 => n40260, C2 => n31439, ZN => n8811);
   U29973 : OAI222_X1 port map( A1 => n40935, A2 => n40270, B1 => n41319, B2 =>
                           n40263, C1 => n40260, C2 => n31438, ZN => n8810);
   U29974 : OAI222_X1 port map( A1 => n40941, A2 => n40270, B1 => n41325, B2 =>
                           n40263, C1 => n40260, C2 => n31437, ZN => n8809);
   U29975 : OAI222_X1 port map( A1 => n40947, A2 => n40270, B1 => n41331, B2 =>
                           n40263, C1 => n40260, C2 => n31436, ZN => n8808);
   U29976 : OAI222_X1 port map( A1 => n40959, A2 => n40270, B1 => n41343, B2 =>
                           n40263, C1 => n40260, C2 => n31434, ZN => n8806);
   U29977 : OAI222_X1 port map( A1 => n40599, A2 => n40255, B1 => n40983, B2 =>
                           n40248, C1 => n40236, C2 => n31430, ZN => n8802);
   U29978 : OAI222_X1 port map( A1 => n40605, A2 => n40255, B1 => n40989, B2 =>
                           n40248, C1 => n40236, C2 => n31429, ZN => n8801);
   U29979 : OAI222_X1 port map( A1 => n40611, A2 => n40255, B1 => n40995, B2 =>
                           n40248, C1 => n40236, C2 => n31428, ZN => n8800);
   U29980 : OAI222_X1 port map( A1 => n40617, A2 => n40255, B1 => n41001, B2 =>
                           n40248, C1 => n40236, C2 => n31427, ZN => n8799);
   U29981 : OAI222_X1 port map( A1 => n40623, A2 => n40254, B1 => n41007, B2 =>
                           n40247, C1 => n40236, C2 => n31426, ZN => n8798);
   U29982 : OAI222_X1 port map( A1 => n40629, A2 => n40254, B1 => n41013, B2 =>
                           n40247, C1 => n40236, C2 => n31425, ZN => n8797);
   U29983 : OAI222_X1 port map( A1 => n40635, A2 => n40254, B1 => n41019, B2 =>
                           n40247, C1 => n40236, C2 => n31424, ZN => n8796);
   U29984 : OAI222_X1 port map( A1 => n40641, A2 => n40254, B1 => n41025, B2 =>
                           n40247, C1 => n40236, C2 => n31423, ZN => n8795);
   U29985 : OAI222_X1 port map( A1 => n40647, A2 => n40254, B1 => n41031, B2 =>
                           n40247, C1 => n40236, C2 => n31422, ZN => n8794);
   U29986 : OAI222_X1 port map( A1 => n40653, A2 => n40254, B1 => n41037, B2 =>
                           n40247, C1 => n40236, C2 => n31421, ZN => n8793);
   U29987 : OAI222_X1 port map( A1 => n40659, A2 => n40254, B1 => n41043, B2 =>
                           n40247, C1 => n40236, C2 => n31420, ZN => n8792);
   U29988 : OAI222_X1 port map( A1 => n40665, A2 => n40254, B1 => n41049, B2 =>
                           n40247, C1 => n40236, C2 => n31419, ZN => n8791);
   U29989 : OAI222_X1 port map( A1 => n40671, A2 => n40254, B1 => n41055, B2 =>
                           n40247, C1 => n40237, C2 => n31418, ZN => n8790);
   U29990 : OAI222_X1 port map( A1 => n40677, A2 => n40254, B1 => n41061, B2 =>
                           n40247, C1 => n40237, C2 => n31417, ZN => n8789);
   U29991 : OAI222_X1 port map( A1 => n40683, A2 => n40254, B1 => n41067, B2 =>
                           n40247, C1 => n40237, C2 => n31416, ZN => n8788);
   U29992 : OAI222_X1 port map( A1 => n40689, A2 => n40254, B1 => n41073, B2 =>
                           n40247, C1 => n40238, C2 => n31415, ZN => n8787);
   U29993 : OAI222_X1 port map( A1 => n40695, A2 => n40253, B1 => n41079, B2 =>
                           n40246, C1 => n40237, C2 => n31414, ZN => n8786);
   U29994 : OAI222_X1 port map( A1 => n40701, A2 => n40253, B1 => n41085, B2 =>
                           n40246, C1 => n40237, C2 => n31413, ZN => n8785);
   U29995 : OAI222_X1 port map( A1 => n40707, A2 => n40253, B1 => n41091, B2 =>
                           n40246, C1 => n40237, C2 => n31412, ZN => n8784);
   U29996 : OAI222_X1 port map( A1 => n40713, A2 => n40253, B1 => n41097, B2 =>
                           n40246, C1 => n40237, C2 => n31411, ZN => n8783);
   U29997 : OAI222_X1 port map( A1 => n40719, A2 => n40253, B1 => n41103, B2 =>
                           n40246, C1 => n40237, C2 => n31410, ZN => n8782);
   U29998 : OAI222_X1 port map( A1 => n40725, A2 => n40253, B1 => n41109, B2 =>
                           n40246, C1 => n40237, C2 => n31409, ZN => n8781);
   U29999 : OAI222_X1 port map( A1 => n40731, A2 => n40253, B1 => n41115, B2 =>
                           n40246, C1 => n40237, C2 => n31408, ZN => n8780);
   U30000 : OAI222_X1 port map( A1 => n40737, A2 => n40253, B1 => n41121, B2 =>
                           n40246, C1 => n40237, C2 => n31407, ZN => n8779);
   U30001 : OAI222_X1 port map( A1 => n40743, A2 => n40253, B1 => n41127, B2 =>
                           n40246, C1 => n40237, C2 => n31406, ZN => n8778);
   U30002 : OAI222_X1 port map( A1 => n40749, A2 => n40253, B1 => n41133, B2 =>
                           n40246, C1 => n40238, C2 => n31405, ZN => n8777);
   U30003 : OAI222_X1 port map( A1 => n40755, A2 => n40253, B1 => n41139, B2 =>
                           n40246, C1 => n40238, C2 => n31404, ZN => n8776);
   U30004 : OAI222_X1 port map( A1 => n40761, A2 => n40253, B1 => n41145, B2 =>
                           n40246, C1 => n40238, C2 => n31403, ZN => n8775);
   U30005 : OAI222_X1 port map( A1 => n40767, A2 => n40252, B1 => n41151, B2 =>
                           n40245, C1 => n40238, C2 => n31402, ZN => n8774);
   U30006 : OAI222_X1 port map( A1 => n40773, A2 => n40252, B1 => n41157, B2 =>
                           n40245, C1 => n40238, C2 => n31401, ZN => n8773);
   U30007 : OAI222_X1 port map( A1 => n40779, A2 => n40252, B1 => n41163, B2 =>
                           n40245, C1 => n40238, C2 => n31400, ZN => n8772);
   U30008 : OAI222_X1 port map( A1 => n40785, A2 => n40252, B1 => n41169, B2 =>
                           n40245, C1 => n40238, C2 => n31399, ZN => n8771);
   U30009 : OAI222_X1 port map( A1 => n40791, A2 => n40252, B1 => n41175, B2 =>
                           n40245, C1 => n40238, C2 => n31398, ZN => n8770);
   U30010 : OAI222_X1 port map( A1 => n40797, A2 => n40252, B1 => n41181, B2 =>
                           n40245, C1 => n40238, C2 => n31397, ZN => n8769);
   U30011 : OAI222_X1 port map( A1 => n40803, A2 => n40252, B1 => n41187, B2 =>
                           n40245, C1 => n40238, C2 => n31396, ZN => n8768);
   U30012 : OAI222_X1 port map( A1 => n40809, A2 => n40252, B1 => n41193, B2 =>
                           n40245, C1 => n40238, C2 => n31395, ZN => n8767);
   U30013 : OAI222_X1 port map( A1 => n40815, A2 => n40252, B1 => n41199, B2 =>
                           n40245, C1 => n40239, C2 => n31394, ZN => n8766);
   U30014 : OAI222_X1 port map( A1 => n40821, A2 => n40252, B1 => n41205, B2 =>
                           n40245, C1 => n40239, C2 => n31393, ZN => n8765);
   U30015 : OAI222_X1 port map( A1 => n40827, A2 => n40252, B1 => n41211, B2 =>
                           n40245, C1 => n40239, C2 => n31392, ZN => n8764);
   U30016 : OAI222_X1 port map( A1 => n40833, A2 => n40252, B1 => n41217, B2 =>
                           n40245, C1 => n40239, C2 => n31391, ZN => n8763);
   U30017 : OAI222_X1 port map( A1 => n40839, A2 => n40251, B1 => n41223, B2 =>
                           n40244, C1 => n40239, C2 => n31390, ZN => n8762);
   U30018 : OAI222_X1 port map( A1 => n40845, A2 => n40251, B1 => n41229, B2 =>
                           n40244, C1 => n40239, C2 => n31389, ZN => n8761);
   U30019 : OAI222_X1 port map( A1 => n40851, A2 => n40251, B1 => n41235, B2 =>
                           n40244, C1 => n40239, C2 => n31388, ZN => n8760);
   U30020 : OAI222_X1 port map( A1 => n40857, A2 => n40251, B1 => n41241, B2 =>
                           n40244, C1 => n40239, C2 => n31387, ZN => n8759);
   U30021 : OAI222_X1 port map( A1 => n40863, A2 => n40251, B1 => n41247, B2 =>
                           n40244, C1 => n40239, C2 => n31386, ZN => n8758);
   U30022 : OAI222_X1 port map( A1 => n40869, A2 => n40251, B1 => n41253, B2 =>
                           n40244, C1 => n40239, C2 => n31385, ZN => n8757);
   U30023 : OAI222_X1 port map( A1 => n40875, A2 => n40251, B1 => n41259, B2 =>
                           n40244, C1 => n40239, C2 => n31384, ZN => n8756);
   U30024 : OAI222_X1 port map( A1 => n40881, A2 => n40251, B1 => n41265, B2 =>
                           n40244, C1 => n40239, C2 => n31383, ZN => n8755);
   U30025 : OAI222_X1 port map( A1 => n40887, A2 => n40251, B1 => n41271, B2 =>
                           n40244, C1 => n40240, C2 => n31382, ZN => n8754);
   U30026 : OAI222_X1 port map( A1 => n40893, A2 => n40251, B1 => n41277, B2 =>
                           n40244, C1 => n40240, C2 => n31381, ZN => n8753);
   U30027 : OAI222_X1 port map( A1 => n40899, A2 => n40251, B1 => n41283, B2 =>
                           n40244, C1 => n40240, C2 => n31380, ZN => n8752);
   U30028 : OAI222_X1 port map( A1 => n40905, A2 => n40251, B1 => n41289, B2 =>
                           n40244, C1 => n40240, C2 => n31379, ZN => n8751);
   U30029 : OAI222_X1 port map( A1 => n40911, A2 => n40250, B1 => n41295, B2 =>
                           n40243, C1 => n40240, C2 => n31378, ZN => n8750);
   U30030 : OAI222_X1 port map( A1 => n40917, A2 => n40250, B1 => n41301, B2 =>
                           n40243, C1 => n40240, C2 => n31377, ZN => n8749);
   U30031 : OAI222_X1 port map( A1 => n40923, A2 => n40250, B1 => n41307, B2 =>
                           n40243, C1 => n40240, C2 => n31376, ZN => n8748);
   U30032 : OAI222_X1 port map( A1 => n40929, A2 => n40250, B1 => n41313, B2 =>
                           n40243, C1 => n40240, C2 => n31375, ZN => n8747);
   U30033 : OAI222_X1 port map( A1 => n40935, A2 => n40250, B1 => n41319, B2 =>
                           n40243, C1 => n40240, C2 => n31374, ZN => n8746);
   U30034 : OAI222_X1 port map( A1 => n40941, A2 => n40250, B1 => n41325, B2 =>
                           n40243, C1 => n40240, C2 => n31373, ZN => n8745);
   U30035 : OAI222_X1 port map( A1 => n40947, A2 => n40250, B1 => n41331, B2 =>
                           n40243, C1 => n40240, C2 => n31372, ZN => n8744);
   U30036 : OAI222_X1 port map( A1 => n40959, A2 => n40250, B1 => n41343, B2 =>
                           n40243, C1 => n40240, C2 => n31370, ZN => n8742);
   U30037 : OAI222_X1 port map( A1 => n40599, A2 => n40195, B1 => n40983, B2 =>
                           n40188, C1 => n40176, C2 => n31366, ZN => n8610);
   U30038 : OAI222_X1 port map( A1 => n40605, A2 => n40195, B1 => n40989, B2 =>
                           n40188, C1 => n40176, C2 => n31365, ZN => n8609);
   U30039 : OAI222_X1 port map( A1 => n40611, A2 => n40195, B1 => n40995, B2 =>
                           n40188, C1 => n40176, C2 => n31364, ZN => n8608);
   U30040 : OAI222_X1 port map( A1 => n40617, A2 => n40195, B1 => n41001, B2 =>
                           n40188, C1 => n40176, C2 => n31363, ZN => n8607);
   U30041 : OAI222_X1 port map( A1 => n40623, A2 => n40194, B1 => n41007, B2 =>
                           n40187, C1 => n40176, C2 => n31362, ZN => n8606);
   U30042 : OAI222_X1 port map( A1 => n40629, A2 => n40194, B1 => n41013, B2 =>
                           n40187, C1 => n40176, C2 => n31361, ZN => n8605);
   U30043 : OAI222_X1 port map( A1 => n40635, A2 => n40194, B1 => n41019, B2 =>
                           n40187, C1 => n40176, C2 => n31360, ZN => n8604);
   U30044 : OAI222_X1 port map( A1 => n40641, A2 => n40194, B1 => n41025, B2 =>
                           n40187, C1 => n40176, C2 => n31359, ZN => n8603);
   U30045 : OAI222_X1 port map( A1 => n40647, A2 => n40194, B1 => n41031, B2 =>
                           n40187, C1 => n40176, C2 => n31358, ZN => n8602);
   U30046 : OAI222_X1 port map( A1 => n40653, A2 => n40194, B1 => n41037, B2 =>
                           n40187, C1 => n40176, C2 => n31357, ZN => n8601);
   U30047 : OAI222_X1 port map( A1 => n40659, A2 => n40194, B1 => n41043, B2 =>
                           n40187, C1 => n40176, C2 => n31356, ZN => n8600);
   U30048 : OAI222_X1 port map( A1 => n40665, A2 => n40194, B1 => n41049, B2 =>
                           n40187, C1 => n40176, C2 => n31355, ZN => n8599);
   U30049 : OAI222_X1 port map( A1 => n40671, A2 => n40194, B1 => n41055, B2 =>
                           n40187, C1 => n40177, C2 => n31354, ZN => n8598);
   U30050 : OAI222_X1 port map( A1 => n40677, A2 => n40194, B1 => n41061, B2 =>
                           n40187, C1 => n40177, C2 => n31353, ZN => n8597);
   U30051 : OAI222_X1 port map( A1 => n40683, A2 => n40194, B1 => n41067, B2 =>
                           n40187, C1 => n40177, C2 => n31352, ZN => n8596);
   U30052 : OAI222_X1 port map( A1 => n40689, A2 => n40194, B1 => n41073, B2 =>
                           n40187, C1 => n40178, C2 => n31351, ZN => n8595);
   U30053 : OAI222_X1 port map( A1 => n40695, A2 => n40193, B1 => n41079, B2 =>
                           n40186, C1 => n40177, C2 => n31350, ZN => n8594);
   U30054 : OAI222_X1 port map( A1 => n40701, A2 => n40193, B1 => n41085, B2 =>
                           n40186, C1 => n40177, C2 => n31349, ZN => n8593);
   U30055 : OAI222_X1 port map( A1 => n40707, A2 => n40193, B1 => n41091, B2 =>
                           n40186, C1 => n40177, C2 => n31348, ZN => n8592);
   U30056 : OAI222_X1 port map( A1 => n40713, A2 => n40193, B1 => n41097, B2 =>
                           n40186, C1 => n40177, C2 => n31347, ZN => n8591);
   U30057 : OAI222_X1 port map( A1 => n40719, A2 => n40193, B1 => n41103, B2 =>
                           n40186, C1 => n40177, C2 => n31346, ZN => n8590);
   U30058 : OAI222_X1 port map( A1 => n40725, A2 => n40193, B1 => n41109, B2 =>
                           n40186, C1 => n40177, C2 => n31345, ZN => n8589);
   U30059 : OAI222_X1 port map( A1 => n40731, A2 => n40193, B1 => n41115, B2 =>
                           n40186, C1 => n40177, C2 => n31344, ZN => n8588);
   U30060 : OAI222_X1 port map( A1 => n40737, A2 => n40193, B1 => n41121, B2 =>
                           n40186, C1 => n40177, C2 => n31343, ZN => n8587);
   U30061 : OAI222_X1 port map( A1 => n40743, A2 => n40193, B1 => n41127, B2 =>
                           n40186, C1 => n40177, C2 => n31342, ZN => n8586);
   U30062 : OAI222_X1 port map( A1 => n40749, A2 => n40193, B1 => n41133, B2 =>
                           n40186, C1 => n40178, C2 => n31341, ZN => n8585);
   U30063 : OAI222_X1 port map( A1 => n40755, A2 => n40193, B1 => n41139, B2 =>
                           n40186, C1 => n40178, C2 => n31340, ZN => n8584);
   U30064 : OAI222_X1 port map( A1 => n40761, A2 => n40193, B1 => n41145, B2 =>
                           n40186, C1 => n40178, C2 => n31339, ZN => n8583);
   U30065 : OAI222_X1 port map( A1 => n40767, A2 => n40192, B1 => n41151, B2 =>
                           n40185, C1 => n40178, C2 => n31338, ZN => n8582);
   U30066 : OAI222_X1 port map( A1 => n40773, A2 => n40192, B1 => n41157, B2 =>
                           n40185, C1 => n40178, C2 => n31337, ZN => n8581);
   U30067 : OAI222_X1 port map( A1 => n40779, A2 => n40192, B1 => n41163, B2 =>
                           n40185, C1 => n40178, C2 => n31336, ZN => n8580);
   U30068 : OAI222_X1 port map( A1 => n40785, A2 => n40192, B1 => n41169, B2 =>
                           n40185, C1 => n40178, C2 => n31335, ZN => n8579);
   U30069 : OAI222_X1 port map( A1 => n40791, A2 => n40192, B1 => n41175, B2 =>
                           n40185, C1 => n40178, C2 => n31334, ZN => n8578);
   U30070 : OAI222_X1 port map( A1 => n40797, A2 => n40192, B1 => n41181, B2 =>
                           n40185, C1 => n40178, C2 => n31333, ZN => n8577);
   U30071 : OAI222_X1 port map( A1 => n40803, A2 => n40192, B1 => n41187, B2 =>
                           n40185, C1 => n40178, C2 => n31332, ZN => n8576);
   U30072 : OAI222_X1 port map( A1 => n40809, A2 => n40192, B1 => n41193, B2 =>
                           n40185, C1 => n40178, C2 => n31331, ZN => n8575);
   U30073 : OAI222_X1 port map( A1 => n40815, A2 => n40192, B1 => n41199, B2 =>
                           n40185, C1 => n40179, C2 => n31330, ZN => n8574);
   U30074 : OAI222_X1 port map( A1 => n40821, A2 => n40192, B1 => n41205, B2 =>
                           n40185, C1 => n40179, C2 => n31329, ZN => n8573);
   U30075 : OAI222_X1 port map( A1 => n40827, A2 => n40192, B1 => n41211, B2 =>
                           n40185, C1 => n40179, C2 => n31328, ZN => n8572);
   U30076 : OAI222_X1 port map( A1 => n40833, A2 => n40192, B1 => n41217, B2 =>
                           n40185, C1 => n40179, C2 => n31327, ZN => n8571);
   U30077 : OAI222_X1 port map( A1 => n40839, A2 => n40191, B1 => n41223, B2 =>
                           n40184, C1 => n40179, C2 => n31326, ZN => n8570);
   U30078 : OAI222_X1 port map( A1 => n40845, A2 => n40191, B1 => n41229, B2 =>
                           n40184, C1 => n40179, C2 => n31325, ZN => n8569);
   U30079 : OAI222_X1 port map( A1 => n40851, A2 => n40191, B1 => n41235, B2 =>
                           n40184, C1 => n40179, C2 => n31324, ZN => n8568);
   U30080 : OAI222_X1 port map( A1 => n40857, A2 => n40191, B1 => n41241, B2 =>
                           n40184, C1 => n40179, C2 => n31323, ZN => n8567);
   U30081 : OAI222_X1 port map( A1 => n40863, A2 => n40191, B1 => n41247, B2 =>
                           n40184, C1 => n40179, C2 => n31322, ZN => n8566);
   U30082 : OAI222_X1 port map( A1 => n40869, A2 => n40191, B1 => n41253, B2 =>
                           n40184, C1 => n40179, C2 => n31321, ZN => n8565);
   U30083 : OAI222_X1 port map( A1 => n40875, A2 => n40191, B1 => n41259, B2 =>
                           n40184, C1 => n40179, C2 => n31320, ZN => n8564);
   U30084 : OAI222_X1 port map( A1 => n40881, A2 => n40191, B1 => n41265, B2 =>
                           n40184, C1 => n40179, C2 => n31319, ZN => n8563);
   U30085 : OAI222_X1 port map( A1 => n40887, A2 => n40191, B1 => n41271, B2 =>
                           n40184, C1 => n40180, C2 => n31318, ZN => n8562);
   U30086 : OAI222_X1 port map( A1 => n40893, A2 => n40191, B1 => n41277, B2 =>
                           n40184, C1 => n40180, C2 => n31317, ZN => n8561);
   U30087 : OAI222_X1 port map( A1 => n40899, A2 => n40191, B1 => n41283, B2 =>
                           n40184, C1 => n40180, C2 => n31316, ZN => n8560);
   U30088 : OAI222_X1 port map( A1 => n40905, A2 => n40191, B1 => n41289, B2 =>
                           n40184, C1 => n40180, C2 => n31315, ZN => n8559);
   U30089 : OAI222_X1 port map( A1 => n40911, A2 => n40190, B1 => n41295, B2 =>
                           n40183, C1 => n40180, C2 => n31314, ZN => n8558);
   U30090 : OAI222_X1 port map( A1 => n40917, A2 => n40190, B1 => n41301, B2 =>
                           n40183, C1 => n40180, C2 => n31313, ZN => n8557);
   U30091 : OAI222_X1 port map( A1 => n40923, A2 => n40190, B1 => n41307, B2 =>
                           n40183, C1 => n40180, C2 => n31312, ZN => n8556);
   U30092 : OAI222_X1 port map( A1 => n40929, A2 => n40190, B1 => n41313, B2 =>
                           n40183, C1 => n40180, C2 => n31311, ZN => n8555);
   U30093 : OAI222_X1 port map( A1 => n40935, A2 => n40190, B1 => n41319, B2 =>
                           n40183, C1 => n40180, C2 => n31310, ZN => n8554);
   U30094 : OAI222_X1 port map( A1 => n40941, A2 => n40190, B1 => n41325, B2 =>
                           n40183, C1 => n40180, C2 => n31309, ZN => n8553);
   U30095 : OAI222_X1 port map( A1 => n40947, A2 => n40190, B1 => n41331, B2 =>
                           n40183, C1 => n40180, C2 => n31308, ZN => n8552);
   U30096 : OAI222_X1 port map( A1 => n40959, A2 => n40190, B1 => n41343, B2 =>
                           n40183, C1 => n40180, C2 => n31306, ZN => n8550);
   U30097 : OAI222_X1 port map( A1 => n40599, A2 => n40175, B1 => n40983, B2 =>
                           n40168, C1 => n40156, C2 => n31302, ZN => n8546);
   U30098 : OAI222_X1 port map( A1 => n40605, A2 => n40175, B1 => n40989, B2 =>
                           n40168, C1 => n40156, C2 => n31301, ZN => n8545);
   U30099 : OAI222_X1 port map( A1 => n40611, A2 => n40175, B1 => n40995, B2 =>
                           n40168, C1 => n40156, C2 => n31300, ZN => n8544);
   U30100 : OAI222_X1 port map( A1 => n40617, A2 => n40175, B1 => n41001, B2 =>
                           n40168, C1 => n40156, C2 => n31299, ZN => n8543);
   U30101 : OAI222_X1 port map( A1 => n40623, A2 => n40174, B1 => n41007, B2 =>
                           n40167, C1 => n40156, C2 => n31298, ZN => n8542);
   U30102 : OAI222_X1 port map( A1 => n40629, A2 => n40174, B1 => n41013, B2 =>
                           n40167, C1 => n40156, C2 => n31297, ZN => n8541);
   U30103 : OAI222_X1 port map( A1 => n40635, A2 => n40174, B1 => n41019, B2 =>
                           n40167, C1 => n40156, C2 => n31296, ZN => n8540);
   U30104 : OAI222_X1 port map( A1 => n40641, A2 => n40174, B1 => n41025, B2 =>
                           n40167, C1 => n40156, C2 => n31295, ZN => n8539);
   U30105 : OAI222_X1 port map( A1 => n40647, A2 => n40174, B1 => n41031, B2 =>
                           n40167, C1 => n40156, C2 => n31294, ZN => n8538);
   U30106 : OAI222_X1 port map( A1 => n40653, A2 => n40174, B1 => n41037, B2 =>
                           n40167, C1 => n40156, C2 => n31293, ZN => n8537);
   U30107 : OAI222_X1 port map( A1 => n40659, A2 => n40174, B1 => n41043, B2 =>
                           n40167, C1 => n40156, C2 => n31292, ZN => n8536);
   U30108 : OAI222_X1 port map( A1 => n40665, A2 => n40174, B1 => n41049, B2 =>
                           n40167, C1 => n40156, C2 => n31291, ZN => n8535);
   U30109 : OAI222_X1 port map( A1 => n40671, A2 => n40174, B1 => n41055, B2 =>
                           n40167, C1 => n40157, C2 => n31290, ZN => n8534);
   U30110 : OAI222_X1 port map( A1 => n40677, A2 => n40174, B1 => n41061, B2 =>
                           n40167, C1 => n40157, C2 => n31289, ZN => n8533);
   U30111 : OAI222_X1 port map( A1 => n40683, A2 => n40174, B1 => n41067, B2 =>
                           n40167, C1 => n40157, C2 => n31288, ZN => n8532);
   U30112 : OAI222_X1 port map( A1 => n40689, A2 => n40174, B1 => n41073, B2 =>
                           n40167, C1 => n40158, C2 => n31287, ZN => n8531);
   U30113 : OAI222_X1 port map( A1 => n40695, A2 => n40173, B1 => n41079, B2 =>
                           n40166, C1 => n40157, C2 => n31286, ZN => n8530);
   U30114 : OAI222_X1 port map( A1 => n40701, A2 => n40173, B1 => n41085, B2 =>
                           n40166, C1 => n40157, C2 => n31285, ZN => n8529);
   U30115 : OAI222_X1 port map( A1 => n40707, A2 => n40173, B1 => n41091, B2 =>
                           n40166, C1 => n40157, C2 => n31284, ZN => n8528);
   U30116 : OAI222_X1 port map( A1 => n40713, A2 => n40173, B1 => n41097, B2 =>
                           n40166, C1 => n40157, C2 => n31283, ZN => n8527);
   U30117 : OAI222_X1 port map( A1 => n40719, A2 => n40173, B1 => n41103, B2 =>
                           n40166, C1 => n40157, C2 => n31282, ZN => n8526);
   U30118 : OAI222_X1 port map( A1 => n40725, A2 => n40173, B1 => n41109, B2 =>
                           n40166, C1 => n40157, C2 => n31281, ZN => n8525);
   U30119 : OAI222_X1 port map( A1 => n40731, A2 => n40173, B1 => n41115, B2 =>
                           n40166, C1 => n40157, C2 => n31280, ZN => n8524);
   U30120 : OAI222_X1 port map( A1 => n40737, A2 => n40173, B1 => n41121, B2 =>
                           n40166, C1 => n40157, C2 => n31279, ZN => n8523);
   U30121 : OAI222_X1 port map( A1 => n40743, A2 => n40173, B1 => n41127, B2 =>
                           n40166, C1 => n40157, C2 => n31278, ZN => n8522);
   U30122 : OAI222_X1 port map( A1 => n40749, A2 => n40173, B1 => n41133, B2 =>
                           n40166, C1 => n40158, C2 => n31277, ZN => n8521);
   U30123 : OAI222_X1 port map( A1 => n40755, A2 => n40173, B1 => n41139, B2 =>
                           n40166, C1 => n40158, C2 => n31276, ZN => n8520);
   U30124 : OAI222_X1 port map( A1 => n40761, A2 => n40173, B1 => n41145, B2 =>
                           n40166, C1 => n40158, C2 => n31275, ZN => n8519);
   U30125 : OAI222_X1 port map( A1 => n40767, A2 => n40172, B1 => n41151, B2 =>
                           n40165, C1 => n40158, C2 => n31274, ZN => n8518);
   U30126 : OAI222_X1 port map( A1 => n40773, A2 => n40172, B1 => n41157, B2 =>
                           n40165, C1 => n40158, C2 => n31273, ZN => n8517);
   U30127 : OAI222_X1 port map( A1 => n40779, A2 => n40172, B1 => n41163, B2 =>
                           n40165, C1 => n40158, C2 => n31272, ZN => n8516);
   U30128 : OAI222_X1 port map( A1 => n40785, A2 => n40172, B1 => n41169, B2 =>
                           n40165, C1 => n40158, C2 => n31271, ZN => n8515);
   U30129 : OAI222_X1 port map( A1 => n40791, A2 => n40172, B1 => n41175, B2 =>
                           n40165, C1 => n40158, C2 => n31270, ZN => n8514);
   U30130 : OAI222_X1 port map( A1 => n40797, A2 => n40172, B1 => n41181, B2 =>
                           n40165, C1 => n40158, C2 => n31269, ZN => n8513);
   U30131 : OAI222_X1 port map( A1 => n40803, A2 => n40172, B1 => n41187, B2 =>
                           n40165, C1 => n40158, C2 => n31268, ZN => n8512);
   U30132 : OAI222_X1 port map( A1 => n40809, A2 => n40172, B1 => n41193, B2 =>
                           n40165, C1 => n40158, C2 => n31267, ZN => n8511);
   U30133 : OAI222_X1 port map( A1 => n40815, A2 => n40172, B1 => n41199, B2 =>
                           n40165, C1 => n40159, C2 => n31266, ZN => n8510);
   U30134 : OAI222_X1 port map( A1 => n40821, A2 => n40172, B1 => n41205, B2 =>
                           n40165, C1 => n40159, C2 => n31265, ZN => n8509);
   U30135 : OAI222_X1 port map( A1 => n40827, A2 => n40172, B1 => n41211, B2 =>
                           n40165, C1 => n40159, C2 => n31264, ZN => n8508);
   U30136 : OAI222_X1 port map( A1 => n40833, A2 => n40172, B1 => n41217, B2 =>
                           n40165, C1 => n40159, C2 => n31263, ZN => n8507);
   U30137 : OAI222_X1 port map( A1 => n40839, A2 => n40171, B1 => n41223, B2 =>
                           n40164, C1 => n40159, C2 => n31262, ZN => n8506);
   U30138 : OAI222_X1 port map( A1 => n40845, A2 => n40171, B1 => n41229, B2 =>
                           n40164, C1 => n40159, C2 => n31261, ZN => n8505);
   U30139 : OAI222_X1 port map( A1 => n40851, A2 => n40171, B1 => n41235, B2 =>
                           n40164, C1 => n40159, C2 => n31260, ZN => n8504);
   U30140 : OAI222_X1 port map( A1 => n40857, A2 => n40171, B1 => n41241, B2 =>
                           n40164, C1 => n40159, C2 => n31259, ZN => n8503);
   U30141 : OAI222_X1 port map( A1 => n40863, A2 => n40171, B1 => n41247, B2 =>
                           n40164, C1 => n40159, C2 => n31258, ZN => n8502);
   U30142 : OAI222_X1 port map( A1 => n40869, A2 => n40171, B1 => n41253, B2 =>
                           n40164, C1 => n40159, C2 => n31257, ZN => n8501);
   U30143 : OAI222_X1 port map( A1 => n40875, A2 => n40171, B1 => n41259, B2 =>
                           n40164, C1 => n40159, C2 => n31256, ZN => n8500);
   U30144 : OAI222_X1 port map( A1 => n40881, A2 => n40171, B1 => n41265, B2 =>
                           n40164, C1 => n40159, C2 => n31255, ZN => n8499);
   U30145 : OAI222_X1 port map( A1 => n40887, A2 => n40171, B1 => n41271, B2 =>
                           n40164, C1 => n40160, C2 => n31254, ZN => n8498);
   U30146 : OAI222_X1 port map( A1 => n40893, A2 => n40171, B1 => n41277, B2 =>
                           n40164, C1 => n40160, C2 => n31253, ZN => n8497);
   U30147 : OAI222_X1 port map( A1 => n40899, A2 => n40171, B1 => n41283, B2 =>
                           n40164, C1 => n40160, C2 => n31252, ZN => n8496);
   U30148 : OAI222_X1 port map( A1 => n40905, A2 => n40171, B1 => n41289, B2 =>
                           n40164, C1 => n40160, C2 => n31251, ZN => n8495);
   U30149 : OAI222_X1 port map( A1 => n40911, A2 => n40170, B1 => n41295, B2 =>
                           n40163, C1 => n40160, C2 => n31250, ZN => n8494);
   U30150 : OAI222_X1 port map( A1 => n40917, A2 => n40170, B1 => n41301, B2 =>
                           n40163, C1 => n40160, C2 => n31249, ZN => n8493);
   U30151 : OAI222_X1 port map( A1 => n40923, A2 => n40170, B1 => n41307, B2 =>
                           n40163, C1 => n40160, C2 => n31248, ZN => n8492);
   U30152 : OAI222_X1 port map( A1 => n40929, A2 => n40170, B1 => n41313, B2 =>
                           n40163, C1 => n40160, C2 => n31247, ZN => n8491);
   U30153 : OAI222_X1 port map( A1 => n40935, A2 => n40170, B1 => n41319, B2 =>
                           n40163, C1 => n40160, C2 => n31246, ZN => n8490);
   U30154 : OAI222_X1 port map( A1 => n40941, A2 => n40170, B1 => n41325, B2 =>
                           n40163, C1 => n40160, C2 => n31245, ZN => n8489);
   U30155 : OAI222_X1 port map( A1 => n40947, A2 => n40170, B1 => n41331, B2 =>
                           n40163, C1 => n40160, C2 => n31244, ZN => n8488);
   U30156 : OAI222_X1 port map( A1 => n40959, A2 => n40170, B1 => n41343, B2 =>
                           n40163, C1 => n40160, C2 => n31242, ZN => n8486);
   U30157 : OAI222_X1 port map( A1 => n40599, A2 => n40155, B1 => n40983, B2 =>
                           n40148, C1 => n40136, C2 => n31238, ZN => n8482);
   U30158 : OAI222_X1 port map( A1 => n40605, A2 => n40155, B1 => n40989, B2 =>
                           n40148, C1 => n40136, C2 => n31237, ZN => n8481);
   U30159 : OAI222_X1 port map( A1 => n40611, A2 => n40155, B1 => n40995, B2 =>
                           n40148, C1 => n40136, C2 => n31236, ZN => n8480);
   U30160 : OAI222_X1 port map( A1 => n40617, A2 => n40155, B1 => n41001, B2 =>
                           n40148, C1 => n40136, C2 => n31235, ZN => n8479);
   U30161 : OAI222_X1 port map( A1 => n40623, A2 => n40154, B1 => n41007, B2 =>
                           n40147, C1 => n40136, C2 => n31234, ZN => n8478);
   U30162 : OAI222_X1 port map( A1 => n40629, A2 => n40154, B1 => n41013, B2 =>
                           n40147, C1 => n40136, C2 => n31233, ZN => n8477);
   U30163 : OAI222_X1 port map( A1 => n40635, A2 => n40154, B1 => n41019, B2 =>
                           n40147, C1 => n40136, C2 => n31232, ZN => n8476);
   U30164 : OAI222_X1 port map( A1 => n40641, A2 => n40154, B1 => n41025, B2 =>
                           n40147, C1 => n40136, C2 => n31231, ZN => n8475);
   U30165 : OAI222_X1 port map( A1 => n40647, A2 => n40154, B1 => n41031, B2 =>
                           n40147, C1 => n40136, C2 => n31230, ZN => n8474);
   U30166 : OAI222_X1 port map( A1 => n40653, A2 => n40154, B1 => n41037, B2 =>
                           n40147, C1 => n40136, C2 => n31229, ZN => n8473);
   U30167 : OAI222_X1 port map( A1 => n40659, A2 => n40154, B1 => n41043, B2 =>
                           n40147, C1 => n40136, C2 => n31228, ZN => n8472);
   U30168 : OAI222_X1 port map( A1 => n40665, A2 => n40154, B1 => n41049, B2 =>
                           n40147, C1 => n40136, C2 => n31227, ZN => n8471);
   U30169 : OAI222_X1 port map( A1 => n40671, A2 => n40154, B1 => n41055, B2 =>
                           n40147, C1 => n40137, C2 => n31226, ZN => n8470);
   U30170 : OAI222_X1 port map( A1 => n40677, A2 => n40154, B1 => n41061, B2 =>
                           n40147, C1 => n40137, C2 => n31225, ZN => n8469);
   U30171 : OAI222_X1 port map( A1 => n40683, A2 => n40154, B1 => n41067, B2 =>
                           n40147, C1 => n40137, C2 => n31224, ZN => n8468);
   U30172 : OAI222_X1 port map( A1 => n40689, A2 => n40154, B1 => n41073, B2 =>
                           n40147, C1 => n40138, C2 => n31223, ZN => n8467);
   U30173 : OAI222_X1 port map( A1 => n40695, A2 => n40153, B1 => n41079, B2 =>
                           n40146, C1 => n40137, C2 => n31222, ZN => n8466);
   U30174 : OAI222_X1 port map( A1 => n40701, A2 => n40153, B1 => n41085, B2 =>
                           n40146, C1 => n40137, C2 => n31221, ZN => n8465);
   U30175 : OAI222_X1 port map( A1 => n40707, A2 => n40153, B1 => n41091, B2 =>
                           n40146, C1 => n40137, C2 => n31220, ZN => n8464);
   U30176 : OAI222_X1 port map( A1 => n40713, A2 => n40153, B1 => n41097, B2 =>
                           n40146, C1 => n40137, C2 => n31219, ZN => n8463);
   U30177 : OAI222_X1 port map( A1 => n40719, A2 => n40153, B1 => n41103, B2 =>
                           n40146, C1 => n40137, C2 => n31218, ZN => n8462);
   U30178 : OAI222_X1 port map( A1 => n40725, A2 => n40153, B1 => n41109, B2 =>
                           n40146, C1 => n40137, C2 => n31217, ZN => n8461);
   U30179 : OAI222_X1 port map( A1 => n40731, A2 => n40153, B1 => n41115, B2 =>
                           n40146, C1 => n40137, C2 => n31216, ZN => n8460);
   U30180 : OAI222_X1 port map( A1 => n40737, A2 => n40153, B1 => n41121, B2 =>
                           n40146, C1 => n40137, C2 => n31215, ZN => n8459);
   U30181 : OAI222_X1 port map( A1 => n40743, A2 => n40153, B1 => n41127, B2 =>
                           n40146, C1 => n40137, C2 => n31214, ZN => n8458);
   U30182 : OAI222_X1 port map( A1 => n40749, A2 => n40153, B1 => n41133, B2 =>
                           n40146, C1 => n40138, C2 => n31213, ZN => n8457);
   U30183 : OAI222_X1 port map( A1 => n40755, A2 => n40153, B1 => n41139, B2 =>
                           n40146, C1 => n40138, C2 => n31212, ZN => n8456);
   U30184 : OAI222_X1 port map( A1 => n40761, A2 => n40153, B1 => n41145, B2 =>
                           n40146, C1 => n40138, C2 => n31211, ZN => n8455);
   U30185 : OAI222_X1 port map( A1 => n40767, A2 => n40152, B1 => n41151, B2 =>
                           n40145, C1 => n40138, C2 => n31210, ZN => n8454);
   U30186 : OAI222_X1 port map( A1 => n40773, A2 => n40152, B1 => n41157, B2 =>
                           n40145, C1 => n40138, C2 => n31209, ZN => n8453);
   U30187 : OAI222_X1 port map( A1 => n40779, A2 => n40152, B1 => n41163, B2 =>
                           n40145, C1 => n40138, C2 => n31208, ZN => n8452);
   U30188 : OAI222_X1 port map( A1 => n40785, A2 => n40152, B1 => n41169, B2 =>
                           n40145, C1 => n40138, C2 => n31207, ZN => n8451);
   U30189 : OAI222_X1 port map( A1 => n40791, A2 => n40152, B1 => n41175, B2 =>
                           n40145, C1 => n40138, C2 => n31206, ZN => n8450);
   U30190 : OAI222_X1 port map( A1 => n40797, A2 => n40152, B1 => n41181, B2 =>
                           n40145, C1 => n40138, C2 => n31205, ZN => n8449);
   U30191 : OAI222_X1 port map( A1 => n40803, A2 => n40152, B1 => n41187, B2 =>
                           n40145, C1 => n40138, C2 => n31204, ZN => n8448);
   U30192 : OAI222_X1 port map( A1 => n40809, A2 => n40152, B1 => n41193, B2 =>
                           n40145, C1 => n40138, C2 => n31203, ZN => n8447);
   U30193 : OAI222_X1 port map( A1 => n40815, A2 => n40152, B1 => n41199, B2 =>
                           n40145, C1 => n40139, C2 => n31202, ZN => n8446);
   U30194 : OAI222_X1 port map( A1 => n40821, A2 => n40152, B1 => n41205, B2 =>
                           n40145, C1 => n40139, C2 => n31201, ZN => n8445);
   U30195 : OAI222_X1 port map( A1 => n40827, A2 => n40152, B1 => n41211, B2 =>
                           n40145, C1 => n40139, C2 => n31200, ZN => n8444);
   U30196 : OAI222_X1 port map( A1 => n40833, A2 => n40152, B1 => n41217, B2 =>
                           n40145, C1 => n40139, C2 => n31199, ZN => n8443);
   U30197 : OAI222_X1 port map( A1 => n40839, A2 => n40151, B1 => n41223, B2 =>
                           n40144, C1 => n40139, C2 => n31198, ZN => n8442);
   U30198 : OAI222_X1 port map( A1 => n40845, A2 => n40151, B1 => n41229, B2 =>
                           n40144, C1 => n40139, C2 => n31197, ZN => n8441);
   U30199 : OAI222_X1 port map( A1 => n40851, A2 => n40151, B1 => n41235, B2 =>
                           n40144, C1 => n40139, C2 => n31196, ZN => n8440);
   U30200 : OAI222_X1 port map( A1 => n40857, A2 => n40151, B1 => n41241, B2 =>
                           n40144, C1 => n40139, C2 => n31195, ZN => n8439);
   U30201 : OAI222_X1 port map( A1 => n40863, A2 => n40151, B1 => n41247, B2 =>
                           n40144, C1 => n40139, C2 => n31194, ZN => n8438);
   U30202 : OAI222_X1 port map( A1 => n40869, A2 => n40151, B1 => n41253, B2 =>
                           n40144, C1 => n40139, C2 => n31193, ZN => n8437);
   U30203 : OAI222_X1 port map( A1 => n40875, A2 => n40151, B1 => n41259, B2 =>
                           n40144, C1 => n40139, C2 => n31192, ZN => n8436);
   U30204 : OAI222_X1 port map( A1 => n40881, A2 => n40151, B1 => n41265, B2 =>
                           n40144, C1 => n40139, C2 => n31191, ZN => n8435);
   U30205 : OAI222_X1 port map( A1 => n40887, A2 => n40151, B1 => n41271, B2 =>
                           n40144, C1 => n40140, C2 => n31190, ZN => n8434);
   U30206 : OAI222_X1 port map( A1 => n40893, A2 => n40151, B1 => n41277, B2 =>
                           n40144, C1 => n40140, C2 => n31189, ZN => n8433);
   U30207 : OAI222_X1 port map( A1 => n40899, A2 => n40151, B1 => n41283, B2 =>
                           n40144, C1 => n40140, C2 => n31188, ZN => n8432);
   U30208 : OAI222_X1 port map( A1 => n40905, A2 => n40151, B1 => n41289, B2 =>
                           n40144, C1 => n40140, C2 => n31187, ZN => n8431);
   U30209 : OAI222_X1 port map( A1 => n40911, A2 => n40150, B1 => n41295, B2 =>
                           n40143, C1 => n40140, C2 => n31186, ZN => n8430);
   U30210 : OAI222_X1 port map( A1 => n40917, A2 => n40150, B1 => n41301, B2 =>
                           n40143, C1 => n40140, C2 => n31185, ZN => n8429);
   U30211 : OAI222_X1 port map( A1 => n40923, A2 => n40150, B1 => n41307, B2 =>
                           n40143, C1 => n40140, C2 => n31184, ZN => n8428);
   U30212 : OAI222_X1 port map( A1 => n40929, A2 => n40150, B1 => n41313, B2 =>
                           n40143, C1 => n40140, C2 => n31183, ZN => n8427);
   U30213 : OAI222_X1 port map( A1 => n40935, A2 => n40150, B1 => n41319, B2 =>
                           n40143, C1 => n40140, C2 => n31182, ZN => n8426);
   U30214 : OAI222_X1 port map( A1 => n40941, A2 => n40150, B1 => n41325, B2 =>
                           n40143, C1 => n40140, C2 => n31181, ZN => n8425);
   U30215 : OAI222_X1 port map( A1 => n40947, A2 => n40150, B1 => n41331, B2 =>
                           n40143, C1 => n40140, C2 => n31180, ZN => n8424);
   U30216 : OAI222_X1 port map( A1 => n40959, A2 => n40150, B1 => n41343, B2 =>
                           n40143, C1 => n40140, C2 => n31178, ZN => n8422);
   U30217 : OAI222_X1 port map( A1 => n40599, A2 => n40096, B1 => n40983, B2 =>
                           n40089, C1 => n40077, C2 => n31056, ZN => n8290);
   U30218 : OAI222_X1 port map( A1 => n40605, A2 => n40096, B1 => n40989, B2 =>
                           n40089, C1 => n40077, C2 => n31055, ZN => n8289);
   U30219 : OAI222_X1 port map( A1 => n40611, A2 => n40096, B1 => n40995, B2 =>
                           n40089, C1 => n40077, C2 => n31054, ZN => n8288);
   U30220 : OAI222_X1 port map( A1 => n40617, A2 => n40096, B1 => n41001, B2 =>
                           n40089, C1 => n40077, C2 => n31053, ZN => n8287);
   U30221 : OAI222_X1 port map( A1 => n40623, A2 => n40095, B1 => n41007, B2 =>
                           n40088, C1 => n40077, C2 => n31052, ZN => n8286);
   U30222 : OAI222_X1 port map( A1 => n40629, A2 => n40095, B1 => n41013, B2 =>
                           n40088, C1 => n40077, C2 => n31051, ZN => n8285);
   U30223 : OAI222_X1 port map( A1 => n40635, A2 => n40095, B1 => n41019, B2 =>
                           n40088, C1 => n40077, C2 => n31050, ZN => n8284);
   U30224 : OAI222_X1 port map( A1 => n40641, A2 => n40095, B1 => n41025, B2 =>
                           n40088, C1 => n40077, C2 => n31049, ZN => n8283);
   U30225 : OAI222_X1 port map( A1 => n40647, A2 => n40095, B1 => n41031, B2 =>
                           n40088, C1 => n40077, C2 => n31048, ZN => n8282);
   U30226 : OAI222_X1 port map( A1 => n40653, A2 => n40095, B1 => n41037, B2 =>
                           n40088, C1 => n40077, C2 => n31047, ZN => n8281);
   U30227 : OAI222_X1 port map( A1 => n40659, A2 => n40095, B1 => n41043, B2 =>
                           n40088, C1 => n40077, C2 => n31046, ZN => n8280);
   U30228 : OAI222_X1 port map( A1 => n40665, A2 => n40095, B1 => n41049, B2 =>
                           n40088, C1 => n40077, C2 => n31045, ZN => n8279);
   U30229 : OAI222_X1 port map( A1 => n40671, A2 => n40095, B1 => n41055, B2 =>
                           n40088, C1 => n40078, C2 => n31044, ZN => n8278);
   U30230 : OAI222_X1 port map( A1 => n40677, A2 => n40095, B1 => n41061, B2 =>
                           n40088, C1 => n40078, C2 => n31043, ZN => n8277);
   U30231 : OAI222_X1 port map( A1 => n40683, A2 => n40095, B1 => n41067, B2 =>
                           n40088, C1 => n40078, C2 => n31042, ZN => n8276);
   U30232 : OAI222_X1 port map( A1 => n40689, A2 => n40095, B1 => n41073, B2 =>
                           n40088, C1 => n40079, C2 => n31041, ZN => n8275);
   U30233 : OAI222_X1 port map( A1 => n40695, A2 => n40094, B1 => n41079, B2 =>
                           n40087, C1 => n40078, C2 => n31040, ZN => n8274);
   U30234 : OAI222_X1 port map( A1 => n40701, A2 => n40094, B1 => n41085, B2 =>
                           n40087, C1 => n40078, C2 => n31039, ZN => n8273);
   U30235 : OAI222_X1 port map( A1 => n40707, A2 => n40094, B1 => n41091, B2 =>
                           n40087, C1 => n40078, C2 => n31038, ZN => n8272);
   U30236 : OAI222_X1 port map( A1 => n40713, A2 => n40094, B1 => n41097, B2 =>
                           n40087, C1 => n40078, C2 => n31037, ZN => n8271);
   U30237 : OAI222_X1 port map( A1 => n40719, A2 => n40094, B1 => n41103, B2 =>
                           n40087, C1 => n40078, C2 => n31036, ZN => n8270);
   U30238 : OAI222_X1 port map( A1 => n40725, A2 => n40094, B1 => n41109, B2 =>
                           n40087, C1 => n40078, C2 => n31035, ZN => n8269);
   U30239 : OAI222_X1 port map( A1 => n40731, A2 => n40094, B1 => n41115, B2 =>
                           n40087, C1 => n40078, C2 => n31034, ZN => n8268);
   U30240 : OAI222_X1 port map( A1 => n40737, A2 => n40094, B1 => n41121, B2 =>
                           n40087, C1 => n40078, C2 => n31033, ZN => n8267);
   U30241 : OAI222_X1 port map( A1 => n40743, A2 => n40094, B1 => n41127, B2 =>
                           n40087, C1 => n40078, C2 => n31032, ZN => n8266);
   U30242 : OAI222_X1 port map( A1 => n40749, A2 => n40094, B1 => n41133, B2 =>
                           n40087, C1 => n40079, C2 => n31031, ZN => n8265);
   U30243 : OAI222_X1 port map( A1 => n40755, A2 => n40094, B1 => n41139, B2 =>
                           n40087, C1 => n40079, C2 => n31030, ZN => n8264);
   U30244 : OAI222_X1 port map( A1 => n40761, A2 => n40094, B1 => n41145, B2 =>
                           n40087, C1 => n40079, C2 => n31029, ZN => n8263);
   U30245 : OAI222_X1 port map( A1 => n40767, A2 => n40093, B1 => n41151, B2 =>
                           n40086, C1 => n40079, C2 => n31028, ZN => n8262);
   U30246 : OAI222_X1 port map( A1 => n40773, A2 => n40093, B1 => n41157, B2 =>
                           n40086, C1 => n40079, C2 => n31027, ZN => n8261);
   U30247 : OAI222_X1 port map( A1 => n40779, A2 => n40093, B1 => n41163, B2 =>
                           n40086, C1 => n40079, C2 => n31026, ZN => n8260);
   U30248 : OAI222_X1 port map( A1 => n40785, A2 => n40093, B1 => n41169, B2 =>
                           n40086, C1 => n40079, C2 => n31025, ZN => n8259);
   U30249 : OAI222_X1 port map( A1 => n40791, A2 => n40093, B1 => n41175, B2 =>
                           n40086, C1 => n40079, C2 => n31024, ZN => n8258);
   U30250 : OAI222_X1 port map( A1 => n40797, A2 => n40093, B1 => n41181, B2 =>
                           n40086, C1 => n40079, C2 => n31023, ZN => n8257);
   U30251 : OAI222_X1 port map( A1 => n40803, A2 => n40093, B1 => n41187, B2 =>
                           n40086, C1 => n40079, C2 => n31022, ZN => n8256);
   U30252 : OAI222_X1 port map( A1 => n40809, A2 => n40093, B1 => n41193, B2 =>
                           n40086, C1 => n40079, C2 => n31021, ZN => n8255);
   U30253 : OAI222_X1 port map( A1 => n40815, A2 => n40093, B1 => n41199, B2 =>
                           n40086, C1 => n40080, C2 => n31020, ZN => n8254);
   U30254 : OAI222_X1 port map( A1 => n40821, A2 => n40093, B1 => n41205, B2 =>
                           n40086, C1 => n40080, C2 => n31019, ZN => n8253);
   U30255 : OAI222_X1 port map( A1 => n40827, A2 => n40093, B1 => n41211, B2 =>
                           n40086, C1 => n40080, C2 => n31018, ZN => n8252);
   U30256 : OAI222_X1 port map( A1 => n40833, A2 => n40093, B1 => n41217, B2 =>
                           n40086, C1 => n40080, C2 => n31017, ZN => n8251);
   U30257 : OAI222_X1 port map( A1 => n40839, A2 => n40092, B1 => n41223, B2 =>
                           n40085, C1 => n40080, C2 => n31016, ZN => n8250);
   U30258 : OAI222_X1 port map( A1 => n40845, A2 => n40092, B1 => n41229, B2 =>
                           n40085, C1 => n40080, C2 => n31015, ZN => n8249);
   U30259 : OAI222_X1 port map( A1 => n40851, A2 => n40092, B1 => n41235, B2 =>
                           n40085, C1 => n40080, C2 => n31014, ZN => n8248);
   U30260 : OAI222_X1 port map( A1 => n40857, A2 => n40092, B1 => n41241, B2 =>
                           n40085, C1 => n40080, C2 => n31013, ZN => n8247);
   U30261 : OAI222_X1 port map( A1 => n40863, A2 => n40092, B1 => n41247, B2 =>
                           n40085, C1 => n40080, C2 => n31012, ZN => n8246);
   U30262 : OAI222_X1 port map( A1 => n40869, A2 => n40092, B1 => n41253, B2 =>
                           n40085, C1 => n40080, C2 => n31011, ZN => n8245);
   U30263 : OAI222_X1 port map( A1 => n40875, A2 => n40092, B1 => n41259, B2 =>
                           n40085, C1 => n40080, C2 => n31010, ZN => n8244);
   U30264 : OAI222_X1 port map( A1 => n40881, A2 => n40092, B1 => n41265, B2 =>
                           n40085, C1 => n40080, C2 => n31009, ZN => n8243);
   U30265 : OAI222_X1 port map( A1 => n40887, A2 => n40092, B1 => n41271, B2 =>
                           n40085, C1 => n40081, C2 => n31008, ZN => n8242);
   U30266 : OAI222_X1 port map( A1 => n40893, A2 => n40092, B1 => n41277, B2 =>
                           n40085, C1 => n40081, C2 => n31007, ZN => n8241);
   U30267 : OAI222_X1 port map( A1 => n40899, A2 => n40092, B1 => n41283, B2 =>
                           n40085, C1 => n40081, C2 => n31006, ZN => n8240);
   U30268 : OAI222_X1 port map( A1 => n40905, A2 => n40092, B1 => n41289, B2 =>
                           n40085, C1 => n40081, C2 => n31005, ZN => n8239);
   U30269 : OAI222_X1 port map( A1 => n40911, A2 => n40091, B1 => n41295, B2 =>
                           n40084, C1 => n40081, C2 => n31004, ZN => n8238);
   U30270 : OAI222_X1 port map( A1 => n40917, A2 => n40091, B1 => n41301, B2 =>
                           n40084, C1 => n40081, C2 => n31003, ZN => n8237);
   U30271 : OAI222_X1 port map( A1 => n40923, A2 => n40091, B1 => n41307, B2 =>
                           n40084, C1 => n40081, C2 => n31002, ZN => n8236);
   U30272 : OAI222_X1 port map( A1 => n40929, A2 => n40091, B1 => n41313, B2 =>
                           n40084, C1 => n40081, C2 => n31001, ZN => n8235);
   U30273 : OAI222_X1 port map( A1 => n40935, A2 => n40091, B1 => n41319, B2 =>
                           n40084, C1 => n40081, C2 => n31000, ZN => n8234);
   U30274 : OAI222_X1 port map( A1 => n40941, A2 => n40091, B1 => n41325, B2 =>
                           n40084, C1 => n40081, C2 => n30999, ZN => n8233);
   U30275 : OAI222_X1 port map( A1 => n40947, A2 => n40091, B1 => n41331, B2 =>
                           n40084, C1 => n40081, C2 => n30998, ZN => n8232);
   U30276 : OAI222_X1 port map( A1 => n40959, A2 => n40091, B1 => n41343, B2 =>
                           n40084, C1 => n40081, C2 => n30996, ZN => n8230);
   U30277 : OAI222_X1 port map( A1 => n40599, A2 => n40076, B1 => n40983, B2 =>
                           n40069, C1 => n40057, C2 => n30992, ZN => n8226);
   U30278 : OAI222_X1 port map( A1 => n40605, A2 => n40076, B1 => n40989, B2 =>
                           n40069, C1 => n40057, C2 => n30991, ZN => n8225);
   U30279 : OAI222_X1 port map( A1 => n40611, A2 => n40076, B1 => n40995, B2 =>
                           n40069, C1 => n40057, C2 => n30990, ZN => n8224);
   U30280 : OAI222_X1 port map( A1 => n40617, A2 => n40076, B1 => n41001, B2 =>
                           n40069, C1 => n40057, C2 => n30989, ZN => n8223);
   U30281 : OAI222_X1 port map( A1 => n40623, A2 => n40075, B1 => n41007, B2 =>
                           n40068, C1 => n40057, C2 => n30988, ZN => n8222);
   U30282 : OAI222_X1 port map( A1 => n40629, A2 => n40075, B1 => n41013, B2 =>
                           n40068, C1 => n40057, C2 => n30987, ZN => n8221);
   U30283 : OAI222_X1 port map( A1 => n40635, A2 => n40075, B1 => n41019, B2 =>
                           n40068, C1 => n40057, C2 => n30986, ZN => n8220);
   U30284 : OAI222_X1 port map( A1 => n40641, A2 => n40075, B1 => n41025, B2 =>
                           n40068, C1 => n40057, C2 => n30985, ZN => n8219);
   U30285 : OAI222_X1 port map( A1 => n40647, A2 => n40075, B1 => n41031, B2 =>
                           n40068, C1 => n40057, C2 => n30984, ZN => n8218);
   U30286 : OAI222_X1 port map( A1 => n40653, A2 => n40075, B1 => n41037, B2 =>
                           n40068, C1 => n40057, C2 => n30983, ZN => n8217);
   U30287 : OAI222_X1 port map( A1 => n40659, A2 => n40075, B1 => n41043, B2 =>
                           n40068, C1 => n40057, C2 => n30982, ZN => n8216);
   U30288 : OAI222_X1 port map( A1 => n40665, A2 => n40075, B1 => n41049, B2 =>
                           n40068, C1 => n40057, C2 => n30981, ZN => n8215);
   U30289 : OAI222_X1 port map( A1 => n40671, A2 => n40075, B1 => n41055, B2 =>
                           n40068, C1 => n40058, C2 => n30980, ZN => n8214);
   U30290 : OAI222_X1 port map( A1 => n40677, A2 => n40075, B1 => n41061, B2 =>
                           n40068, C1 => n40058, C2 => n30979, ZN => n8213);
   U30291 : OAI222_X1 port map( A1 => n40683, A2 => n40075, B1 => n41067, B2 =>
                           n40068, C1 => n40058, C2 => n30978, ZN => n8212);
   U30292 : OAI222_X1 port map( A1 => n40689, A2 => n40075, B1 => n41073, B2 =>
                           n40068, C1 => n40059, C2 => n30977, ZN => n8211);
   U30293 : OAI222_X1 port map( A1 => n40695, A2 => n40074, B1 => n41079, B2 =>
                           n40067, C1 => n40058, C2 => n30976, ZN => n8210);
   U30294 : OAI222_X1 port map( A1 => n40701, A2 => n40074, B1 => n41085, B2 =>
                           n40067, C1 => n40058, C2 => n30975, ZN => n8209);
   U30295 : OAI222_X1 port map( A1 => n40707, A2 => n40074, B1 => n41091, B2 =>
                           n40067, C1 => n40058, C2 => n30974, ZN => n8208);
   U30296 : OAI222_X1 port map( A1 => n40713, A2 => n40074, B1 => n41097, B2 =>
                           n40067, C1 => n40058, C2 => n30973, ZN => n8207);
   U30297 : OAI222_X1 port map( A1 => n40719, A2 => n40074, B1 => n41103, B2 =>
                           n40067, C1 => n40058, C2 => n30972, ZN => n8206);
   U30298 : OAI222_X1 port map( A1 => n40725, A2 => n40074, B1 => n41109, B2 =>
                           n40067, C1 => n40058, C2 => n30971, ZN => n8205);
   U30299 : OAI222_X1 port map( A1 => n40731, A2 => n40074, B1 => n41115, B2 =>
                           n40067, C1 => n40058, C2 => n30970, ZN => n8204);
   U30300 : OAI222_X1 port map( A1 => n40737, A2 => n40074, B1 => n41121, B2 =>
                           n40067, C1 => n40058, C2 => n30969, ZN => n8203);
   U30301 : OAI222_X1 port map( A1 => n40743, A2 => n40074, B1 => n41127, B2 =>
                           n40067, C1 => n40058, C2 => n30968, ZN => n8202);
   U30302 : OAI222_X1 port map( A1 => n40749, A2 => n40074, B1 => n41133, B2 =>
                           n40067, C1 => n40059, C2 => n30967, ZN => n8201);
   U30303 : OAI222_X1 port map( A1 => n40755, A2 => n40074, B1 => n41139, B2 =>
                           n40067, C1 => n40059, C2 => n30966, ZN => n8200);
   U30304 : OAI222_X1 port map( A1 => n40761, A2 => n40074, B1 => n41145, B2 =>
                           n40067, C1 => n40059, C2 => n30965, ZN => n8199);
   U30305 : OAI222_X1 port map( A1 => n40767, A2 => n40073, B1 => n41151, B2 =>
                           n40066, C1 => n40059, C2 => n30964, ZN => n8198);
   U30306 : OAI222_X1 port map( A1 => n40773, A2 => n40073, B1 => n41157, B2 =>
                           n40066, C1 => n40059, C2 => n30963, ZN => n8197);
   U30307 : OAI222_X1 port map( A1 => n40779, A2 => n40073, B1 => n41163, B2 =>
                           n40066, C1 => n40059, C2 => n30962, ZN => n8196);
   U30308 : OAI222_X1 port map( A1 => n40785, A2 => n40073, B1 => n41169, B2 =>
                           n40066, C1 => n40059, C2 => n30961, ZN => n8195);
   U30309 : OAI222_X1 port map( A1 => n40791, A2 => n40073, B1 => n41175, B2 =>
                           n40066, C1 => n40059, C2 => n30960, ZN => n8194);
   U30310 : OAI222_X1 port map( A1 => n40797, A2 => n40073, B1 => n41181, B2 =>
                           n40066, C1 => n40059, C2 => n30959, ZN => n8193);
   U30311 : OAI222_X1 port map( A1 => n40803, A2 => n40073, B1 => n41187, B2 =>
                           n40066, C1 => n40059, C2 => n30958, ZN => n8192);
   U30312 : OAI222_X1 port map( A1 => n40809, A2 => n40073, B1 => n41193, B2 =>
                           n40066, C1 => n40059, C2 => n30957, ZN => n8191);
   U30313 : OAI222_X1 port map( A1 => n40815, A2 => n40073, B1 => n41199, B2 =>
                           n40066, C1 => n40060, C2 => n30956, ZN => n8190);
   U30314 : OAI222_X1 port map( A1 => n40821, A2 => n40073, B1 => n41205, B2 =>
                           n40066, C1 => n40060, C2 => n30955, ZN => n8189);
   U30315 : OAI222_X1 port map( A1 => n40827, A2 => n40073, B1 => n41211, B2 =>
                           n40066, C1 => n40060, C2 => n30954, ZN => n8188);
   U30316 : OAI222_X1 port map( A1 => n40833, A2 => n40073, B1 => n41217, B2 =>
                           n40066, C1 => n40060, C2 => n30953, ZN => n8187);
   U30317 : OAI222_X1 port map( A1 => n40839, A2 => n40072, B1 => n41223, B2 =>
                           n40065, C1 => n40060, C2 => n30952, ZN => n8186);
   U30318 : OAI222_X1 port map( A1 => n40845, A2 => n40072, B1 => n41229, B2 =>
                           n40065, C1 => n40060, C2 => n30951, ZN => n8185);
   U30319 : OAI222_X1 port map( A1 => n40851, A2 => n40072, B1 => n41235, B2 =>
                           n40065, C1 => n40060, C2 => n30950, ZN => n8184);
   U30320 : OAI222_X1 port map( A1 => n40857, A2 => n40072, B1 => n41241, B2 =>
                           n40065, C1 => n40060, C2 => n30949, ZN => n8183);
   U30321 : OAI222_X1 port map( A1 => n40863, A2 => n40072, B1 => n41247, B2 =>
                           n40065, C1 => n40060, C2 => n30948, ZN => n8182);
   U30322 : OAI222_X1 port map( A1 => n40869, A2 => n40072, B1 => n41253, B2 =>
                           n40065, C1 => n40060, C2 => n30947, ZN => n8181);
   U30323 : OAI222_X1 port map( A1 => n40875, A2 => n40072, B1 => n41259, B2 =>
                           n40065, C1 => n40060, C2 => n30946, ZN => n8180);
   U30324 : OAI222_X1 port map( A1 => n40881, A2 => n40072, B1 => n41265, B2 =>
                           n40065, C1 => n40060, C2 => n30945, ZN => n8179);
   U30325 : OAI222_X1 port map( A1 => n40887, A2 => n40072, B1 => n41271, B2 =>
                           n40065, C1 => n40061, C2 => n30944, ZN => n8178);
   U30326 : OAI222_X1 port map( A1 => n40893, A2 => n40072, B1 => n41277, B2 =>
                           n40065, C1 => n40061, C2 => n30943, ZN => n8177);
   U30327 : OAI222_X1 port map( A1 => n40899, A2 => n40072, B1 => n41283, B2 =>
                           n40065, C1 => n40061, C2 => n30942, ZN => n8176);
   U30328 : OAI222_X1 port map( A1 => n40905, A2 => n40072, B1 => n41289, B2 =>
                           n40065, C1 => n40061, C2 => n30941, ZN => n8175);
   U30329 : OAI222_X1 port map( A1 => n40911, A2 => n40071, B1 => n41295, B2 =>
                           n40064, C1 => n40061, C2 => n30940, ZN => n8174);
   U30330 : OAI222_X1 port map( A1 => n40917, A2 => n40071, B1 => n41301, B2 =>
                           n40064, C1 => n40061, C2 => n30939, ZN => n8173);
   U30331 : OAI222_X1 port map( A1 => n40923, A2 => n40071, B1 => n41307, B2 =>
                           n40064, C1 => n40061, C2 => n30938, ZN => n8172);
   U30332 : OAI222_X1 port map( A1 => n40929, A2 => n40071, B1 => n41313, B2 =>
                           n40064, C1 => n40061, C2 => n30937, ZN => n8171);
   U30333 : OAI222_X1 port map( A1 => n40935, A2 => n40071, B1 => n41319, B2 =>
                           n40064, C1 => n40061, C2 => n30936, ZN => n8170);
   U30334 : OAI222_X1 port map( A1 => n40941, A2 => n40071, B1 => n41325, B2 =>
                           n40064, C1 => n40061, C2 => n30935, ZN => n8169);
   U30335 : OAI222_X1 port map( A1 => n40947, A2 => n40071, B1 => n41331, B2 =>
                           n40064, C1 => n40061, C2 => n30934, ZN => n8168);
   U30336 : OAI222_X1 port map( A1 => n40959, A2 => n40071, B1 => n41343, B2 =>
                           n40064, C1 => n40061, C2 => n30932, ZN => n8166);
   U30337 : OAI222_X1 port map( A1 => n40599, A2 => n40056, B1 => n40983, B2 =>
                           n40049, C1 => n40037, C2 => n30928, ZN => n8162);
   U30338 : OAI222_X1 port map( A1 => n40605, A2 => n40056, B1 => n40989, B2 =>
                           n40049, C1 => n40037, C2 => n30927, ZN => n8161);
   U30339 : OAI222_X1 port map( A1 => n40611, A2 => n40056, B1 => n40995, B2 =>
                           n40049, C1 => n40037, C2 => n30926, ZN => n8160);
   U30340 : OAI222_X1 port map( A1 => n40617, A2 => n40056, B1 => n41001, B2 =>
                           n40049, C1 => n40037, C2 => n30925, ZN => n8159);
   U30341 : OAI222_X1 port map( A1 => n40623, A2 => n40055, B1 => n41007, B2 =>
                           n40048, C1 => n40037, C2 => n30924, ZN => n8158);
   U30342 : OAI222_X1 port map( A1 => n40629, A2 => n40055, B1 => n41013, B2 =>
                           n40048, C1 => n40037, C2 => n30923, ZN => n8157);
   U30343 : OAI222_X1 port map( A1 => n40635, A2 => n40055, B1 => n41019, B2 =>
                           n40048, C1 => n40037, C2 => n30922, ZN => n8156);
   U30344 : OAI222_X1 port map( A1 => n40641, A2 => n40055, B1 => n41025, B2 =>
                           n40048, C1 => n40037, C2 => n30921, ZN => n8155);
   U30345 : OAI222_X1 port map( A1 => n40647, A2 => n40055, B1 => n41031, B2 =>
                           n40048, C1 => n40037, C2 => n30920, ZN => n8154);
   U30346 : OAI222_X1 port map( A1 => n40653, A2 => n40055, B1 => n41037, B2 =>
                           n40048, C1 => n40037, C2 => n30919, ZN => n8153);
   U30347 : OAI222_X1 port map( A1 => n40659, A2 => n40055, B1 => n41043, B2 =>
                           n40048, C1 => n40037, C2 => n30918, ZN => n8152);
   U30348 : OAI222_X1 port map( A1 => n40665, A2 => n40055, B1 => n41049, B2 =>
                           n40048, C1 => n40037, C2 => n30917, ZN => n8151);
   U30349 : OAI222_X1 port map( A1 => n40671, A2 => n40055, B1 => n41055, B2 =>
                           n40048, C1 => n40038, C2 => n30916, ZN => n8150);
   U30350 : OAI222_X1 port map( A1 => n40677, A2 => n40055, B1 => n41061, B2 =>
                           n40048, C1 => n40038, C2 => n30915, ZN => n8149);
   U30351 : OAI222_X1 port map( A1 => n40683, A2 => n40055, B1 => n41067, B2 =>
                           n40048, C1 => n40038, C2 => n30914, ZN => n8148);
   U30352 : OAI222_X1 port map( A1 => n40689, A2 => n40055, B1 => n41073, B2 =>
                           n40048, C1 => n40039, C2 => n30913, ZN => n8147);
   U30353 : OAI222_X1 port map( A1 => n40695, A2 => n40054, B1 => n41079, B2 =>
                           n40047, C1 => n40038, C2 => n30912, ZN => n8146);
   U30354 : OAI222_X1 port map( A1 => n40701, A2 => n40054, B1 => n41085, B2 =>
                           n40047, C1 => n40038, C2 => n30911, ZN => n8145);
   U30355 : OAI222_X1 port map( A1 => n40707, A2 => n40054, B1 => n41091, B2 =>
                           n40047, C1 => n40038, C2 => n30910, ZN => n8144);
   U30356 : OAI222_X1 port map( A1 => n40713, A2 => n40054, B1 => n41097, B2 =>
                           n40047, C1 => n40038, C2 => n30909, ZN => n8143);
   U30357 : OAI222_X1 port map( A1 => n40719, A2 => n40054, B1 => n41103, B2 =>
                           n40047, C1 => n40038, C2 => n30908, ZN => n8142);
   U30358 : OAI222_X1 port map( A1 => n40725, A2 => n40054, B1 => n41109, B2 =>
                           n40047, C1 => n40038, C2 => n30907, ZN => n8141);
   U30359 : OAI222_X1 port map( A1 => n40731, A2 => n40054, B1 => n41115, B2 =>
                           n40047, C1 => n40038, C2 => n30906, ZN => n8140);
   U30360 : OAI222_X1 port map( A1 => n40737, A2 => n40054, B1 => n41121, B2 =>
                           n40047, C1 => n40038, C2 => n30905, ZN => n8139);
   U30361 : OAI222_X1 port map( A1 => n40743, A2 => n40054, B1 => n41127, B2 =>
                           n40047, C1 => n40038, C2 => n30904, ZN => n8138);
   U30362 : OAI222_X1 port map( A1 => n40749, A2 => n40054, B1 => n41133, B2 =>
                           n40047, C1 => n40039, C2 => n30903, ZN => n8137);
   U30363 : OAI222_X1 port map( A1 => n40755, A2 => n40054, B1 => n41139, B2 =>
                           n40047, C1 => n40039, C2 => n30902, ZN => n8136);
   U30364 : OAI222_X1 port map( A1 => n40761, A2 => n40054, B1 => n41145, B2 =>
                           n40047, C1 => n40039, C2 => n30901, ZN => n8135);
   U30365 : OAI222_X1 port map( A1 => n40767, A2 => n40053, B1 => n41151, B2 =>
                           n40046, C1 => n40039, C2 => n30900, ZN => n8134);
   U30366 : OAI222_X1 port map( A1 => n40773, A2 => n40053, B1 => n41157, B2 =>
                           n40046, C1 => n40039, C2 => n30899, ZN => n8133);
   U30367 : OAI222_X1 port map( A1 => n40779, A2 => n40053, B1 => n41163, B2 =>
                           n40046, C1 => n40039, C2 => n30898, ZN => n8132);
   U30368 : OAI222_X1 port map( A1 => n40785, A2 => n40053, B1 => n41169, B2 =>
                           n40046, C1 => n40039, C2 => n30897, ZN => n8131);
   U30369 : OAI222_X1 port map( A1 => n40791, A2 => n40053, B1 => n41175, B2 =>
                           n40046, C1 => n40039, C2 => n30896, ZN => n8130);
   U30370 : OAI222_X1 port map( A1 => n40797, A2 => n40053, B1 => n41181, B2 =>
                           n40046, C1 => n40039, C2 => n30895, ZN => n8129);
   U30371 : OAI222_X1 port map( A1 => n40803, A2 => n40053, B1 => n41187, B2 =>
                           n40046, C1 => n40039, C2 => n30894, ZN => n8128);
   U30372 : OAI222_X1 port map( A1 => n40809, A2 => n40053, B1 => n41193, B2 =>
                           n40046, C1 => n40039, C2 => n30893, ZN => n8127);
   U30373 : OAI222_X1 port map( A1 => n40815, A2 => n40053, B1 => n41199, B2 =>
                           n40046, C1 => n40040, C2 => n30892, ZN => n8126);
   U30374 : OAI222_X1 port map( A1 => n40821, A2 => n40053, B1 => n41205, B2 =>
                           n40046, C1 => n40040, C2 => n30891, ZN => n8125);
   U30375 : OAI222_X1 port map( A1 => n40827, A2 => n40053, B1 => n41211, B2 =>
                           n40046, C1 => n40040, C2 => n30890, ZN => n8124);
   U30376 : OAI222_X1 port map( A1 => n40833, A2 => n40053, B1 => n41217, B2 =>
                           n40046, C1 => n40040, C2 => n30889, ZN => n8123);
   U30377 : OAI222_X1 port map( A1 => n40839, A2 => n40052, B1 => n41223, B2 =>
                           n40045, C1 => n40040, C2 => n30888, ZN => n8122);
   U30378 : OAI222_X1 port map( A1 => n40845, A2 => n40052, B1 => n41229, B2 =>
                           n40045, C1 => n40040, C2 => n30887, ZN => n8121);
   U30379 : OAI222_X1 port map( A1 => n40851, A2 => n40052, B1 => n41235, B2 =>
                           n40045, C1 => n40040, C2 => n30886, ZN => n8120);
   U30380 : OAI222_X1 port map( A1 => n40857, A2 => n40052, B1 => n41241, B2 =>
                           n40045, C1 => n40040, C2 => n30885, ZN => n8119);
   U30381 : OAI222_X1 port map( A1 => n40863, A2 => n40052, B1 => n41247, B2 =>
                           n40045, C1 => n40040, C2 => n30884, ZN => n8118);
   U30382 : OAI222_X1 port map( A1 => n40869, A2 => n40052, B1 => n41253, B2 =>
                           n40045, C1 => n40040, C2 => n30883, ZN => n8117);
   U30383 : OAI222_X1 port map( A1 => n40875, A2 => n40052, B1 => n41259, B2 =>
                           n40045, C1 => n40040, C2 => n30882, ZN => n8116);
   U30384 : OAI222_X1 port map( A1 => n40881, A2 => n40052, B1 => n41265, B2 =>
                           n40045, C1 => n40040, C2 => n30881, ZN => n8115);
   U30385 : OAI222_X1 port map( A1 => n40887, A2 => n40052, B1 => n41271, B2 =>
                           n40045, C1 => n40041, C2 => n30880, ZN => n8114);
   U30386 : OAI222_X1 port map( A1 => n40893, A2 => n40052, B1 => n41277, B2 =>
                           n40045, C1 => n40041, C2 => n30879, ZN => n8113);
   U30387 : OAI222_X1 port map( A1 => n40899, A2 => n40052, B1 => n41283, B2 =>
                           n40045, C1 => n40041, C2 => n30878, ZN => n8112);
   U30388 : OAI222_X1 port map( A1 => n40905, A2 => n40052, B1 => n41289, B2 =>
                           n40045, C1 => n40041, C2 => n30877, ZN => n8111);
   U30389 : OAI222_X1 port map( A1 => n40911, A2 => n40051, B1 => n41295, B2 =>
                           n40044, C1 => n40041, C2 => n30876, ZN => n8110);
   U30390 : OAI222_X1 port map( A1 => n40917, A2 => n40051, B1 => n41301, B2 =>
                           n40044, C1 => n40041, C2 => n30875, ZN => n8109);
   U30391 : OAI222_X1 port map( A1 => n40923, A2 => n40051, B1 => n41307, B2 =>
                           n40044, C1 => n40041, C2 => n30874, ZN => n8108);
   U30392 : OAI222_X1 port map( A1 => n40929, A2 => n40051, B1 => n41313, B2 =>
                           n40044, C1 => n40041, C2 => n30873, ZN => n8107);
   U30393 : OAI222_X1 port map( A1 => n40935, A2 => n40051, B1 => n41319, B2 =>
                           n40044, C1 => n40041, C2 => n30872, ZN => n8106);
   U30394 : OAI222_X1 port map( A1 => n40941, A2 => n40051, B1 => n41325, B2 =>
                           n40044, C1 => n40041, C2 => n30871, ZN => n8105);
   U30395 : OAI222_X1 port map( A1 => n40947, A2 => n40051, B1 => n41331, B2 =>
                           n40044, C1 => n40041, C2 => n30870, ZN => n8104);
   U30396 : OAI222_X1 port map( A1 => n40959, A2 => n40051, B1 => n41343, B2 =>
                           n40044, C1 => n40041, C2 => n30868, ZN => n8102);
   U30397 : OAI222_X1 port map( A1 => n40598, A2 => n39998, B1 => n40982, B2 =>
                           n39991, C1 => n39979, C2 => n30864, ZN => n7970);
   U30398 : OAI222_X1 port map( A1 => n40604, A2 => n39998, B1 => n40988, B2 =>
                           n39991, C1 => n39979, C2 => n30863, ZN => n7969);
   U30399 : OAI222_X1 port map( A1 => n40610, A2 => n39998, B1 => n40994, B2 =>
                           n39991, C1 => n39979, C2 => n30862, ZN => n7968);
   U30400 : OAI222_X1 port map( A1 => n40616, A2 => n39998, B1 => n41000, B2 =>
                           n39991, C1 => n39979, C2 => n30861, ZN => n7967);
   U30401 : OAI222_X1 port map( A1 => n40622, A2 => n39997, B1 => n41006, B2 =>
                           n39990, C1 => n39979, C2 => n30860, ZN => n7966);
   U30402 : OAI222_X1 port map( A1 => n40628, A2 => n39997, B1 => n41012, B2 =>
                           n39990, C1 => n39979, C2 => n30859, ZN => n7965);
   U30403 : OAI222_X1 port map( A1 => n40634, A2 => n39997, B1 => n41018, B2 =>
                           n39990, C1 => n39979, C2 => n30858, ZN => n7964);
   U30404 : OAI222_X1 port map( A1 => n40640, A2 => n39997, B1 => n41024, B2 =>
                           n39990, C1 => n39979, C2 => n30857, ZN => n7963);
   U30405 : OAI222_X1 port map( A1 => n40646, A2 => n39997, B1 => n41030, B2 =>
                           n39990, C1 => n39979, C2 => n30856, ZN => n7962);
   U30406 : OAI222_X1 port map( A1 => n40652, A2 => n39997, B1 => n41036, B2 =>
                           n39990, C1 => n39979, C2 => n30855, ZN => n7961);
   U30407 : OAI222_X1 port map( A1 => n40658, A2 => n39997, B1 => n41042, B2 =>
                           n39990, C1 => n39979, C2 => n30854, ZN => n7960);
   U30408 : OAI222_X1 port map( A1 => n40664, A2 => n39997, B1 => n41048, B2 =>
                           n39990, C1 => n39979, C2 => n30853, ZN => n7959);
   U30409 : OAI222_X1 port map( A1 => n40670, A2 => n39997, B1 => n41054, B2 =>
                           n39990, C1 => n39980, C2 => n30852, ZN => n7958);
   U30410 : OAI222_X1 port map( A1 => n40676, A2 => n39997, B1 => n41060, B2 =>
                           n39990, C1 => n39980, C2 => n30851, ZN => n7957);
   U30411 : OAI222_X1 port map( A1 => n40682, A2 => n39997, B1 => n41066, B2 =>
                           n39990, C1 => n39980, C2 => n30850, ZN => n7956);
   U30412 : OAI222_X1 port map( A1 => n40688, A2 => n39997, B1 => n41072, B2 =>
                           n39990, C1 => n39981, C2 => n30849, ZN => n7955);
   U30413 : OAI222_X1 port map( A1 => n40694, A2 => n39996, B1 => n41078, B2 =>
                           n39989, C1 => n39980, C2 => n30848, ZN => n7954);
   U30414 : OAI222_X1 port map( A1 => n40700, A2 => n39996, B1 => n41084, B2 =>
                           n39989, C1 => n39980, C2 => n30847, ZN => n7953);
   U30415 : OAI222_X1 port map( A1 => n40706, A2 => n39996, B1 => n41090, B2 =>
                           n39989, C1 => n39980, C2 => n30846, ZN => n7952);
   U30416 : OAI222_X1 port map( A1 => n40712, A2 => n39996, B1 => n41096, B2 =>
                           n39989, C1 => n39980, C2 => n30845, ZN => n7951);
   U30417 : OAI222_X1 port map( A1 => n40718, A2 => n39996, B1 => n41102, B2 =>
                           n39989, C1 => n39980, C2 => n30844, ZN => n7950);
   U30418 : OAI222_X1 port map( A1 => n40724, A2 => n39996, B1 => n41108, B2 =>
                           n39989, C1 => n39980, C2 => n30843, ZN => n7949);
   U30419 : OAI222_X1 port map( A1 => n40730, A2 => n39996, B1 => n41114, B2 =>
                           n39989, C1 => n39980, C2 => n30842, ZN => n7948);
   U30420 : OAI222_X1 port map( A1 => n40736, A2 => n39996, B1 => n41120, B2 =>
                           n39989, C1 => n39980, C2 => n30841, ZN => n7947);
   U30421 : OAI222_X1 port map( A1 => n40742, A2 => n39996, B1 => n41126, B2 =>
                           n39989, C1 => n39980, C2 => n30840, ZN => n7946);
   U30422 : OAI222_X1 port map( A1 => n40748, A2 => n39996, B1 => n41132, B2 =>
                           n39989, C1 => n39981, C2 => n30839, ZN => n7945);
   U30423 : OAI222_X1 port map( A1 => n40754, A2 => n39996, B1 => n41138, B2 =>
                           n39989, C1 => n39981, C2 => n30838, ZN => n7944);
   U30424 : OAI222_X1 port map( A1 => n40760, A2 => n39996, B1 => n41144, B2 =>
                           n39989, C1 => n39981, C2 => n30837, ZN => n7943);
   U30425 : OAI222_X1 port map( A1 => n40766, A2 => n39995, B1 => n41150, B2 =>
                           n39988, C1 => n39981, C2 => n30836, ZN => n7942);
   U30426 : OAI222_X1 port map( A1 => n40772, A2 => n39995, B1 => n41156, B2 =>
                           n39988, C1 => n39981, C2 => n30835, ZN => n7941);
   U30427 : OAI222_X1 port map( A1 => n40778, A2 => n39995, B1 => n41162, B2 =>
                           n39988, C1 => n39981, C2 => n30834, ZN => n7940);
   U30428 : OAI222_X1 port map( A1 => n40784, A2 => n39995, B1 => n41168, B2 =>
                           n39988, C1 => n39981, C2 => n30833, ZN => n7939);
   U30429 : OAI222_X1 port map( A1 => n40790, A2 => n39995, B1 => n41174, B2 =>
                           n39988, C1 => n39981, C2 => n30832, ZN => n7938);
   U30430 : OAI222_X1 port map( A1 => n40796, A2 => n39995, B1 => n41180, B2 =>
                           n39988, C1 => n39981, C2 => n30831, ZN => n7937);
   U30431 : OAI222_X1 port map( A1 => n40802, A2 => n39995, B1 => n41186, B2 =>
                           n39988, C1 => n39981, C2 => n30830, ZN => n7936);
   U30432 : OAI222_X1 port map( A1 => n40808, A2 => n39995, B1 => n41192, B2 =>
                           n39988, C1 => n39981, C2 => n30829, ZN => n7935);
   U30433 : OAI222_X1 port map( A1 => n40814, A2 => n39995, B1 => n41198, B2 =>
                           n39988, C1 => n39982, C2 => n30828, ZN => n7934);
   U30434 : OAI222_X1 port map( A1 => n40820, A2 => n39995, B1 => n41204, B2 =>
                           n39988, C1 => n39982, C2 => n30827, ZN => n7933);
   U30435 : OAI222_X1 port map( A1 => n40826, A2 => n39995, B1 => n41210, B2 =>
                           n39988, C1 => n39982, C2 => n30826, ZN => n7932);
   U30436 : OAI222_X1 port map( A1 => n40832, A2 => n39995, B1 => n41216, B2 =>
                           n39988, C1 => n39982, C2 => n30825, ZN => n7931);
   U30437 : OAI222_X1 port map( A1 => n40838, A2 => n39994, B1 => n41222, B2 =>
                           n39987, C1 => n39982, C2 => n30824, ZN => n7930);
   U30438 : OAI222_X1 port map( A1 => n40844, A2 => n39994, B1 => n41228, B2 =>
                           n39987, C1 => n39982, C2 => n30823, ZN => n7929);
   U30439 : OAI222_X1 port map( A1 => n40850, A2 => n39994, B1 => n41234, B2 =>
                           n39987, C1 => n39982, C2 => n30822, ZN => n7928);
   U30440 : OAI222_X1 port map( A1 => n40856, A2 => n39994, B1 => n41240, B2 =>
                           n39987, C1 => n39982, C2 => n30821, ZN => n7927);
   U30441 : OAI222_X1 port map( A1 => n40862, A2 => n39994, B1 => n41246, B2 =>
                           n39987, C1 => n39982, C2 => n30820, ZN => n7926);
   U30442 : OAI222_X1 port map( A1 => n40868, A2 => n39994, B1 => n41252, B2 =>
                           n39987, C1 => n39982, C2 => n30819, ZN => n7925);
   U30443 : OAI222_X1 port map( A1 => n40874, A2 => n39994, B1 => n41258, B2 =>
                           n39987, C1 => n39982, C2 => n30818, ZN => n7924);
   U30444 : OAI222_X1 port map( A1 => n40880, A2 => n39994, B1 => n41264, B2 =>
                           n39987, C1 => n39982, C2 => n30817, ZN => n7923);
   U30445 : OAI222_X1 port map( A1 => n40886, A2 => n39994, B1 => n41270, B2 =>
                           n39987, C1 => n39983, C2 => n30816, ZN => n7922);
   U30446 : OAI222_X1 port map( A1 => n40892, A2 => n39994, B1 => n41276, B2 =>
                           n39987, C1 => n39983, C2 => n30815, ZN => n7921);
   U30447 : OAI222_X1 port map( A1 => n40898, A2 => n39994, B1 => n41282, B2 =>
                           n39987, C1 => n39983, C2 => n30814, ZN => n7920);
   U30448 : OAI222_X1 port map( A1 => n40904, A2 => n39994, B1 => n41288, B2 =>
                           n39987, C1 => n39983, C2 => n30813, ZN => n7919);
   U30449 : OAI222_X1 port map( A1 => n40910, A2 => n39993, B1 => n41294, B2 =>
                           n39986, C1 => n39983, C2 => n30812, ZN => n7918);
   U30450 : OAI222_X1 port map( A1 => n40916, A2 => n39993, B1 => n41300, B2 =>
                           n39986, C1 => n39983, C2 => n30811, ZN => n7917);
   U30451 : OAI222_X1 port map( A1 => n40922, A2 => n39993, B1 => n41306, B2 =>
                           n39986, C1 => n39983, C2 => n30810, ZN => n7916);
   U30452 : OAI222_X1 port map( A1 => n40928, A2 => n39993, B1 => n41312, B2 =>
                           n39986, C1 => n39983, C2 => n30809, ZN => n7915);
   U30453 : OAI222_X1 port map( A1 => n40934, A2 => n39993, B1 => n41318, B2 =>
                           n39986, C1 => n39983, C2 => n30808, ZN => n7914);
   U30454 : OAI222_X1 port map( A1 => n40940, A2 => n39993, B1 => n41324, B2 =>
                           n39986, C1 => n39983, C2 => n30807, ZN => n7913);
   U30455 : OAI222_X1 port map( A1 => n40946, A2 => n39993, B1 => n41330, B2 =>
                           n39986, C1 => n39983, C2 => n30806, ZN => n7912);
   U30456 : OAI222_X1 port map( A1 => n40958, A2 => n39993, B1 => n41342, B2 =>
                           n39986, C1 => n39983, C2 => n30804, ZN => n7910);
   U30457 : OAI222_X1 port map( A1 => n40598, A2 => n39978, B1 => n40982, B2 =>
                           n39971, C1 => n39959, C2 => n30800, ZN => n7906);
   U30458 : OAI222_X1 port map( A1 => n40604, A2 => n39978, B1 => n40988, B2 =>
                           n39971, C1 => n39959, C2 => n30799, ZN => n7905);
   U30459 : OAI222_X1 port map( A1 => n40610, A2 => n39978, B1 => n40994, B2 =>
                           n39971, C1 => n39959, C2 => n30798, ZN => n7904);
   U30460 : OAI222_X1 port map( A1 => n40616, A2 => n39978, B1 => n41000, B2 =>
                           n39971, C1 => n39959, C2 => n30797, ZN => n7903);
   U30461 : OAI222_X1 port map( A1 => n40622, A2 => n39977, B1 => n41006, B2 =>
                           n39970, C1 => n39959, C2 => n30796, ZN => n7902);
   U30462 : OAI222_X1 port map( A1 => n40628, A2 => n39977, B1 => n41012, B2 =>
                           n39970, C1 => n39959, C2 => n30795, ZN => n7901);
   U30463 : OAI222_X1 port map( A1 => n40634, A2 => n39977, B1 => n41018, B2 =>
                           n39970, C1 => n39959, C2 => n30794, ZN => n7900);
   U30464 : OAI222_X1 port map( A1 => n40640, A2 => n39977, B1 => n41024, B2 =>
                           n39970, C1 => n39959, C2 => n30793, ZN => n7899);
   U30465 : OAI222_X1 port map( A1 => n40646, A2 => n39977, B1 => n41030, B2 =>
                           n39970, C1 => n39959, C2 => n30792, ZN => n7898);
   U30466 : OAI222_X1 port map( A1 => n40652, A2 => n39977, B1 => n41036, B2 =>
                           n39970, C1 => n39959, C2 => n30791, ZN => n7897);
   U30467 : OAI222_X1 port map( A1 => n40658, A2 => n39977, B1 => n41042, B2 =>
                           n39970, C1 => n39959, C2 => n30790, ZN => n7896);
   U30468 : OAI222_X1 port map( A1 => n40664, A2 => n39977, B1 => n41048, B2 =>
                           n39970, C1 => n39959, C2 => n30789, ZN => n7895);
   U30469 : OAI222_X1 port map( A1 => n40670, A2 => n39977, B1 => n41054, B2 =>
                           n39970, C1 => n39960, C2 => n30788, ZN => n7894);
   U30470 : OAI222_X1 port map( A1 => n40676, A2 => n39977, B1 => n41060, B2 =>
                           n39970, C1 => n39960, C2 => n30787, ZN => n7893);
   U30471 : OAI222_X1 port map( A1 => n40682, A2 => n39977, B1 => n41066, B2 =>
                           n39970, C1 => n39960, C2 => n30786, ZN => n7892);
   U30472 : OAI222_X1 port map( A1 => n40688, A2 => n39977, B1 => n41072, B2 =>
                           n39970, C1 => n39961, C2 => n30785, ZN => n7891);
   U30473 : OAI222_X1 port map( A1 => n40694, A2 => n39976, B1 => n41078, B2 =>
                           n39969, C1 => n39960, C2 => n30784, ZN => n7890);
   U30474 : OAI222_X1 port map( A1 => n40700, A2 => n39976, B1 => n41084, B2 =>
                           n39969, C1 => n39960, C2 => n30783, ZN => n7889);
   U30475 : OAI222_X1 port map( A1 => n40706, A2 => n39976, B1 => n41090, B2 =>
                           n39969, C1 => n39960, C2 => n30782, ZN => n7888);
   U30476 : OAI222_X1 port map( A1 => n40712, A2 => n39976, B1 => n41096, B2 =>
                           n39969, C1 => n39960, C2 => n30781, ZN => n7887);
   U30477 : OAI222_X1 port map( A1 => n40718, A2 => n39976, B1 => n41102, B2 =>
                           n39969, C1 => n39960, C2 => n30780, ZN => n7886);
   U30478 : OAI222_X1 port map( A1 => n40724, A2 => n39976, B1 => n41108, B2 =>
                           n39969, C1 => n39960, C2 => n30779, ZN => n7885);
   U30479 : OAI222_X1 port map( A1 => n40730, A2 => n39976, B1 => n41114, B2 =>
                           n39969, C1 => n39960, C2 => n30778, ZN => n7884);
   U30480 : OAI222_X1 port map( A1 => n40736, A2 => n39976, B1 => n41120, B2 =>
                           n39969, C1 => n39960, C2 => n30777, ZN => n7883);
   U30481 : OAI222_X1 port map( A1 => n40742, A2 => n39976, B1 => n41126, B2 =>
                           n39969, C1 => n39960, C2 => n30776, ZN => n7882);
   U30482 : OAI222_X1 port map( A1 => n40748, A2 => n39976, B1 => n41132, B2 =>
                           n39969, C1 => n39961, C2 => n30775, ZN => n7881);
   U30483 : OAI222_X1 port map( A1 => n40754, A2 => n39976, B1 => n41138, B2 =>
                           n39969, C1 => n39961, C2 => n30774, ZN => n7880);
   U30484 : OAI222_X1 port map( A1 => n40760, A2 => n39976, B1 => n41144, B2 =>
                           n39969, C1 => n39961, C2 => n30773, ZN => n7879);
   U30485 : OAI222_X1 port map( A1 => n40766, A2 => n39975, B1 => n41150, B2 =>
                           n39968, C1 => n39961, C2 => n30772, ZN => n7878);
   U30486 : OAI222_X1 port map( A1 => n40772, A2 => n39975, B1 => n41156, B2 =>
                           n39968, C1 => n39961, C2 => n30771, ZN => n7877);
   U30487 : OAI222_X1 port map( A1 => n40778, A2 => n39975, B1 => n41162, B2 =>
                           n39968, C1 => n39961, C2 => n30770, ZN => n7876);
   U30488 : OAI222_X1 port map( A1 => n40784, A2 => n39975, B1 => n41168, B2 =>
                           n39968, C1 => n39961, C2 => n30769, ZN => n7875);
   U30489 : OAI222_X1 port map( A1 => n40790, A2 => n39975, B1 => n41174, B2 =>
                           n39968, C1 => n39961, C2 => n30768, ZN => n7874);
   U30490 : OAI222_X1 port map( A1 => n40796, A2 => n39975, B1 => n41180, B2 =>
                           n39968, C1 => n39961, C2 => n30767, ZN => n7873);
   U30491 : OAI222_X1 port map( A1 => n40802, A2 => n39975, B1 => n41186, B2 =>
                           n39968, C1 => n39961, C2 => n30766, ZN => n7872);
   U30492 : OAI222_X1 port map( A1 => n40808, A2 => n39975, B1 => n41192, B2 =>
                           n39968, C1 => n39961, C2 => n30765, ZN => n7871);
   U30493 : OAI222_X1 port map( A1 => n40814, A2 => n39975, B1 => n41198, B2 =>
                           n39968, C1 => n39962, C2 => n30764, ZN => n7870);
   U30494 : OAI222_X1 port map( A1 => n40820, A2 => n39975, B1 => n41204, B2 =>
                           n39968, C1 => n39962, C2 => n30763, ZN => n7869);
   U30495 : OAI222_X1 port map( A1 => n40826, A2 => n39975, B1 => n41210, B2 =>
                           n39968, C1 => n39962, C2 => n30762, ZN => n7868);
   U30496 : OAI222_X1 port map( A1 => n40832, A2 => n39975, B1 => n41216, B2 =>
                           n39968, C1 => n39962, C2 => n30761, ZN => n7867);
   U30497 : OAI222_X1 port map( A1 => n40838, A2 => n39974, B1 => n41222, B2 =>
                           n39967, C1 => n39962, C2 => n30760, ZN => n7866);
   U30498 : OAI222_X1 port map( A1 => n40844, A2 => n39974, B1 => n41228, B2 =>
                           n39967, C1 => n39962, C2 => n30759, ZN => n7865);
   U30499 : OAI222_X1 port map( A1 => n40850, A2 => n39974, B1 => n41234, B2 =>
                           n39967, C1 => n39962, C2 => n30758, ZN => n7864);
   U30500 : OAI222_X1 port map( A1 => n40856, A2 => n39974, B1 => n41240, B2 =>
                           n39967, C1 => n39962, C2 => n30757, ZN => n7863);
   U30501 : OAI222_X1 port map( A1 => n40862, A2 => n39974, B1 => n41246, B2 =>
                           n39967, C1 => n39962, C2 => n30756, ZN => n7862);
   U30502 : OAI222_X1 port map( A1 => n40868, A2 => n39974, B1 => n41252, B2 =>
                           n39967, C1 => n39962, C2 => n30755, ZN => n7861);
   U30503 : OAI222_X1 port map( A1 => n40874, A2 => n39974, B1 => n41258, B2 =>
                           n39967, C1 => n39962, C2 => n30754, ZN => n7860);
   U30504 : OAI222_X1 port map( A1 => n40880, A2 => n39974, B1 => n41264, B2 =>
                           n39967, C1 => n39962, C2 => n30753, ZN => n7859);
   U30505 : OAI222_X1 port map( A1 => n40886, A2 => n39974, B1 => n41270, B2 =>
                           n39967, C1 => n39963, C2 => n30752, ZN => n7858);
   U30506 : OAI222_X1 port map( A1 => n40892, A2 => n39974, B1 => n41276, B2 =>
                           n39967, C1 => n39963, C2 => n30751, ZN => n7857);
   U30507 : OAI222_X1 port map( A1 => n40898, A2 => n39974, B1 => n41282, B2 =>
                           n39967, C1 => n39963, C2 => n30750, ZN => n7856);
   U30508 : OAI222_X1 port map( A1 => n40904, A2 => n39974, B1 => n41288, B2 =>
                           n39967, C1 => n39963, C2 => n30749, ZN => n7855);
   U30509 : OAI222_X1 port map( A1 => n40910, A2 => n39973, B1 => n41294, B2 =>
                           n39966, C1 => n39963, C2 => n30748, ZN => n7854);
   U30510 : OAI222_X1 port map( A1 => n40916, A2 => n39973, B1 => n41300, B2 =>
                           n39966, C1 => n39963, C2 => n30747, ZN => n7853);
   U30511 : OAI222_X1 port map( A1 => n40922, A2 => n39973, B1 => n41306, B2 =>
                           n39966, C1 => n39963, C2 => n30746, ZN => n7852);
   U30512 : OAI222_X1 port map( A1 => n40928, A2 => n39973, B1 => n41312, B2 =>
                           n39966, C1 => n39963, C2 => n30745, ZN => n7851);
   U30513 : OAI222_X1 port map( A1 => n40934, A2 => n39973, B1 => n41318, B2 =>
                           n39966, C1 => n39963, C2 => n30744, ZN => n7850);
   U30514 : OAI222_X1 port map( A1 => n40940, A2 => n39973, B1 => n41324, B2 =>
                           n39966, C1 => n39963, C2 => n30743, ZN => n7849);
   U30515 : OAI222_X1 port map( A1 => n40946, A2 => n39973, B1 => n41330, B2 =>
                           n39966, C1 => n39963, C2 => n30742, ZN => n7848);
   U30516 : OAI222_X1 port map( A1 => n40958, A2 => n39973, B1 => n41342, B2 =>
                           n39966, C1 => n39963, C2 => n30740, ZN => n7846);
   U30517 : OAI222_X1 port map( A1 => n40598, A2 => n39958, B1 => n40982, B2 =>
                           n39951, C1 => n39939, C2 => n30736, ZN => n7842);
   U30518 : OAI222_X1 port map( A1 => n40604, A2 => n39958, B1 => n40988, B2 =>
                           n39951, C1 => n39939, C2 => n30735, ZN => n7841);
   U30519 : OAI222_X1 port map( A1 => n40610, A2 => n39958, B1 => n40994, B2 =>
                           n39951, C1 => n39939, C2 => n30734, ZN => n7840);
   U30520 : OAI222_X1 port map( A1 => n40616, A2 => n39958, B1 => n41000, B2 =>
                           n39951, C1 => n39939, C2 => n30733, ZN => n7839);
   U30521 : OAI222_X1 port map( A1 => n40622, A2 => n39957, B1 => n41006, B2 =>
                           n39950, C1 => n39939, C2 => n30732, ZN => n7838);
   U30522 : OAI222_X1 port map( A1 => n40628, A2 => n39957, B1 => n41012, B2 =>
                           n39950, C1 => n39939, C2 => n30731, ZN => n7837);
   U30523 : OAI222_X1 port map( A1 => n40634, A2 => n39957, B1 => n41018, B2 =>
                           n39950, C1 => n39939, C2 => n30730, ZN => n7836);
   U30524 : OAI222_X1 port map( A1 => n40640, A2 => n39957, B1 => n41024, B2 =>
                           n39950, C1 => n39939, C2 => n30729, ZN => n7835);
   U30525 : OAI222_X1 port map( A1 => n40646, A2 => n39957, B1 => n41030, B2 =>
                           n39950, C1 => n39939, C2 => n30728, ZN => n7834);
   U30526 : OAI222_X1 port map( A1 => n40652, A2 => n39957, B1 => n41036, B2 =>
                           n39950, C1 => n39939, C2 => n30727, ZN => n7833);
   U30527 : OAI222_X1 port map( A1 => n40658, A2 => n39957, B1 => n41042, B2 =>
                           n39950, C1 => n39939, C2 => n30726, ZN => n7832);
   U30528 : OAI222_X1 port map( A1 => n40664, A2 => n39957, B1 => n41048, B2 =>
                           n39950, C1 => n39939, C2 => n30725, ZN => n7831);
   U30529 : OAI222_X1 port map( A1 => n40670, A2 => n39957, B1 => n41054, B2 =>
                           n39950, C1 => n39940, C2 => n30724, ZN => n7830);
   U30530 : OAI222_X1 port map( A1 => n40676, A2 => n39957, B1 => n41060, B2 =>
                           n39950, C1 => n39940, C2 => n30723, ZN => n7829);
   U30531 : OAI222_X1 port map( A1 => n40682, A2 => n39957, B1 => n41066, B2 =>
                           n39950, C1 => n39940, C2 => n30722, ZN => n7828);
   U30532 : OAI222_X1 port map( A1 => n40688, A2 => n39957, B1 => n41072, B2 =>
                           n39950, C1 => n39941, C2 => n30721, ZN => n7827);
   U30533 : OAI222_X1 port map( A1 => n40694, A2 => n39956, B1 => n41078, B2 =>
                           n39949, C1 => n39940, C2 => n30720, ZN => n7826);
   U30534 : OAI222_X1 port map( A1 => n40700, A2 => n39956, B1 => n41084, B2 =>
                           n39949, C1 => n39940, C2 => n30719, ZN => n7825);
   U30535 : OAI222_X1 port map( A1 => n40706, A2 => n39956, B1 => n41090, B2 =>
                           n39949, C1 => n39940, C2 => n30718, ZN => n7824);
   U30536 : OAI222_X1 port map( A1 => n40712, A2 => n39956, B1 => n41096, B2 =>
                           n39949, C1 => n39940, C2 => n30717, ZN => n7823);
   U30537 : OAI222_X1 port map( A1 => n40718, A2 => n39956, B1 => n41102, B2 =>
                           n39949, C1 => n39940, C2 => n30716, ZN => n7822);
   U30538 : OAI222_X1 port map( A1 => n40724, A2 => n39956, B1 => n41108, B2 =>
                           n39949, C1 => n39940, C2 => n30715, ZN => n7821);
   U30539 : OAI222_X1 port map( A1 => n40730, A2 => n39956, B1 => n41114, B2 =>
                           n39949, C1 => n39940, C2 => n30714, ZN => n7820);
   U30540 : OAI222_X1 port map( A1 => n40736, A2 => n39956, B1 => n41120, B2 =>
                           n39949, C1 => n39940, C2 => n30713, ZN => n7819);
   U30541 : OAI222_X1 port map( A1 => n40742, A2 => n39956, B1 => n41126, B2 =>
                           n39949, C1 => n39940, C2 => n30712, ZN => n7818);
   U30542 : OAI222_X1 port map( A1 => n40748, A2 => n39956, B1 => n41132, B2 =>
                           n39949, C1 => n39941, C2 => n30711, ZN => n7817);
   U30543 : OAI222_X1 port map( A1 => n40754, A2 => n39956, B1 => n41138, B2 =>
                           n39949, C1 => n39941, C2 => n30710, ZN => n7816);
   U30544 : OAI222_X1 port map( A1 => n40760, A2 => n39956, B1 => n41144, B2 =>
                           n39949, C1 => n39941, C2 => n30709, ZN => n7815);
   U30545 : OAI222_X1 port map( A1 => n40766, A2 => n39955, B1 => n41150, B2 =>
                           n39948, C1 => n39941, C2 => n30708, ZN => n7814);
   U30546 : OAI222_X1 port map( A1 => n40772, A2 => n39955, B1 => n41156, B2 =>
                           n39948, C1 => n39941, C2 => n30707, ZN => n7813);
   U30547 : OAI222_X1 port map( A1 => n40778, A2 => n39955, B1 => n41162, B2 =>
                           n39948, C1 => n39941, C2 => n30706, ZN => n7812);
   U30548 : OAI222_X1 port map( A1 => n40784, A2 => n39955, B1 => n41168, B2 =>
                           n39948, C1 => n39941, C2 => n30705, ZN => n7811);
   U30549 : OAI222_X1 port map( A1 => n40790, A2 => n39955, B1 => n41174, B2 =>
                           n39948, C1 => n39941, C2 => n30704, ZN => n7810);
   U30550 : OAI222_X1 port map( A1 => n40796, A2 => n39955, B1 => n41180, B2 =>
                           n39948, C1 => n39941, C2 => n30703, ZN => n7809);
   U30551 : OAI222_X1 port map( A1 => n40802, A2 => n39955, B1 => n41186, B2 =>
                           n39948, C1 => n39941, C2 => n30702, ZN => n7808);
   U30552 : OAI222_X1 port map( A1 => n40808, A2 => n39955, B1 => n41192, B2 =>
                           n39948, C1 => n39941, C2 => n30701, ZN => n7807);
   U30553 : OAI222_X1 port map( A1 => n40814, A2 => n39955, B1 => n41198, B2 =>
                           n39948, C1 => n39942, C2 => n30700, ZN => n7806);
   U30554 : OAI222_X1 port map( A1 => n40820, A2 => n39955, B1 => n41204, B2 =>
                           n39948, C1 => n39942, C2 => n30699, ZN => n7805);
   U30555 : OAI222_X1 port map( A1 => n40826, A2 => n39955, B1 => n41210, B2 =>
                           n39948, C1 => n39942, C2 => n30698, ZN => n7804);
   U30556 : OAI222_X1 port map( A1 => n40832, A2 => n39955, B1 => n41216, B2 =>
                           n39948, C1 => n39942, C2 => n30697, ZN => n7803);
   U30557 : OAI222_X1 port map( A1 => n40838, A2 => n39954, B1 => n41222, B2 =>
                           n39947, C1 => n39942, C2 => n30696, ZN => n7802);
   U30558 : OAI222_X1 port map( A1 => n40844, A2 => n39954, B1 => n41228, B2 =>
                           n39947, C1 => n39942, C2 => n30695, ZN => n7801);
   U30559 : OAI222_X1 port map( A1 => n40850, A2 => n39954, B1 => n41234, B2 =>
                           n39947, C1 => n39942, C2 => n30694, ZN => n7800);
   U30560 : OAI222_X1 port map( A1 => n40856, A2 => n39954, B1 => n41240, B2 =>
                           n39947, C1 => n39942, C2 => n30693, ZN => n7799);
   U30561 : OAI222_X1 port map( A1 => n40862, A2 => n39954, B1 => n41246, B2 =>
                           n39947, C1 => n39942, C2 => n30692, ZN => n7798);
   U30562 : OAI222_X1 port map( A1 => n40868, A2 => n39954, B1 => n41252, B2 =>
                           n39947, C1 => n39942, C2 => n30691, ZN => n7797);
   U30563 : OAI222_X1 port map( A1 => n40874, A2 => n39954, B1 => n41258, B2 =>
                           n39947, C1 => n39942, C2 => n30690, ZN => n7796);
   U30564 : OAI222_X1 port map( A1 => n40880, A2 => n39954, B1 => n41264, B2 =>
                           n39947, C1 => n39942, C2 => n30689, ZN => n7795);
   U30565 : OAI222_X1 port map( A1 => n40886, A2 => n39954, B1 => n41270, B2 =>
                           n39947, C1 => n39943, C2 => n30688, ZN => n7794);
   U30566 : OAI222_X1 port map( A1 => n40892, A2 => n39954, B1 => n41276, B2 =>
                           n39947, C1 => n39943, C2 => n30687, ZN => n7793);
   U30567 : OAI222_X1 port map( A1 => n40898, A2 => n39954, B1 => n41282, B2 =>
                           n39947, C1 => n39943, C2 => n30686, ZN => n7792);
   U30568 : OAI222_X1 port map( A1 => n40904, A2 => n39954, B1 => n41288, B2 =>
                           n39947, C1 => n39943, C2 => n30685, ZN => n7791);
   U30569 : OAI222_X1 port map( A1 => n40910, A2 => n39953, B1 => n41294, B2 =>
                           n39946, C1 => n39943, C2 => n30684, ZN => n7790);
   U30570 : OAI222_X1 port map( A1 => n40916, A2 => n39953, B1 => n41300, B2 =>
                           n39946, C1 => n39943, C2 => n30683, ZN => n7789);
   U30571 : OAI222_X1 port map( A1 => n40922, A2 => n39953, B1 => n41306, B2 =>
                           n39946, C1 => n39943, C2 => n30682, ZN => n7788);
   U30572 : OAI222_X1 port map( A1 => n40928, A2 => n39953, B1 => n41312, B2 =>
                           n39946, C1 => n39943, C2 => n30681, ZN => n7787);
   U30573 : OAI222_X1 port map( A1 => n40934, A2 => n39953, B1 => n41318, B2 =>
                           n39946, C1 => n39943, C2 => n30680, ZN => n7786);
   U30574 : OAI222_X1 port map( A1 => n40940, A2 => n39953, B1 => n41324, B2 =>
                           n39946, C1 => n39943, C2 => n30679, ZN => n7785);
   U30575 : OAI222_X1 port map( A1 => n40946, A2 => n39953, B1 => n41330, B2 =>
                           n39946, C1 => n39943, C2 => n30678, ZN => n7784);
   U30576 : OAI222_X1 port map( A1 => n40958, A2 => n39953, B1 => n41342, B2 =>
                           n39946, C1 => n39943, C2 => n30676, ZN => n7782);
   U30577 : OAI222_X1 port map( A1 => n40598, A2 => n39900, B1 => n40982, B2 =>
                           n39893, C1 => n39881, C2 => n30672, ZN => n7650);
   U30578 : OAI222_X1 port map( A1 => n40604, A2 => n39900, B1 => n40988, B2 =>
                           n39893, C1 => n39881, C2 => n30671, ZN => n7649);
   U30579 : OAI222_X1 port map( A1 => n40610, A2 => n39900, B1 => n40994, B2 =>
                           n39893, C1 => n39881, C2 => n30670, ZN => n7648);
   U30580 : OAI222_X1 port map( A1 => n40616, A2 => n39900, B1 => n41000, B2 =>
                           n39893, C1 => n39881, C2 => n30669, ZN => n7647);
   U30581 : OAI222_X1 port map( A1 => n40622, A2 => n39899, B1 => n41006, B2 =>
                           n39892, C1 => n39881, C2 => n30668, ZN => n7646);
   U30582 : OAI222_X1 port map( A1 => n40628, A2 => n39899, B1 => n41012, B2 =>
                           n39892, C1 => n39881, C2 => n30667, ZN => n7645);
   U30583 : OAI222_X1 port map( A1 => n40634, A2 => n39899, B1 => n41018, B2 =>
                           n39892, C1 => n39881, C2 => n30666, ZN => n7644);
   U30584 : OAI222_X1 port map( A1 => n40640, A2 => n39899, B1 => n41024, B2 =>
                           n39892, C1 => n39881, C2 => n30665, ZN => n7643);
   U30585 : OAI222_X1 port map( A1 => n40646, A2 => n39899, B1 => n41030, B2 =>
                           n39892, C1 => n39881, C2 => n30664, ZN => n7642);
   U30586 : OAI222_X1 port map( A1 => n40652, A2 => n39899, B1 => n41036, B2 =>
                           n39892, C1 => n39881, C2 => n30663, ZN => n7641);
   U30587 : OAI222_X1 port map( A1 => n40658, A2 => n39899, B1 => n41042, B2 =>
                           n39892, C1 => n39881, C2 => n30662, ZN => n7640);
   U30588 : OAI222_X1 port map( A1 => n40664, A2 => n39899, B1 => n41048, B2 =>
                           n39892, C1 => n39881, C2 => n30661, ZN => n7639);
   U30589 : OAI222_X1 port map( A1 => n40670, A2 => n39899, B1 => n41054, B2 =>
                           n39892, C1 => n39882, C2 => n30660, ZN => n7638);
   U30590 : OAI222_X1 port map( A1 => n40676, A2 => n39899, B1 => n41060, B2 =>
                           n39892, C1 => n39882, C2 => n30659, ZN => n7637);
   U30591 : OAI222_X1 port map( A1 => n40682, A2 => n39899, B1 => n41066, B2 =>
                           n39892, C1 => n39882, C2 => n30658, ZN => n7636);
   U30592 : OAI222_X1 port map( A1 => n40688, A2 => n39899, B1 => n41072, B2 =>
                           n39892, C1 => n39883, C2 => n30657, ZN => n7635);
   U30593 : OAI222_X1 port map( A1 => n40694, A2 => n39898, B1 => n41078, B2 =>
                           n39891, C1 => n39882, C2 => n30656, ZN => n7634);
   U30594 : OAI222_X1 port map( A1 => n40700, A2 => n39898, B1 => n41084, B2 =>
                           n39891, C1 => n39882, C2 => n30655, ZN => n7633);
   U30595 : OAI222_X1 port map( A1 => n40706, A2 => n39898, B1 => n41090, B2 =>
                           n39891, C1 => n39882, C2 => n30654, ZN => n7632);
   U30596 : OAI222_X1 port map( A1 => n40712, A2 => n39898, B1 => n41096, B2 =>
                           n39891, C1 => n39882, C2 => n30653, ZN => n7631);
   U30597 : OAI222_X1 port map( A1 => n40718, A2 => n39898, B1 => n41102, B2 =>
                           n39891, C1 => n39882, C2 => n30652, ZN => n7630);
   U30598 : OAI222_X1 port map( A1 => n40724, A2 => n39898, B1 => n41108, B2 =>
                           n39891, C1 => n39882, C2 => n30651, ZN => n7629);
   U30599 : OAI222_X1 port map( A1 => n40730, A2 => n39898, B1 => n41114, B2 =>
                           n39891, C1 => n39882, C2 => n30650, ZN => n7628);
   U30600 : OAI222_X1 port map( A1 => n40736, A2 => n39898, B1 => n41120, B2 =>
                           n39891, C1 => n39882, C2 => n30649, ZN => n7627);
   U30601 : OAI222_X1 port map( A1 => n40742, A2 => n39898, B1 => n41126, B2 =>
                           n39891, C1 => n39882, C2 => n30648, ZN => n7626);
   U30602 : OAI222_X1 port map( A1 => n40748, A2 => n39898, B1 => n41132, B2 =>
                           n39891, C1 => n39883, C2 => n30647, ZN => n7625);
   U30603 : OAI222_X1 port map( A1 => n40754, A2 => n39898, B1 => n41138, B2 =>
                           n39891, C1 => n39883, C2 => n30646, ZN => n7624);
   U30604 : OAI222_X1 port map( A1 => n40760, A2 => n39898, B1 => n41144, B2 =>
                           n39891, C1 => n39883, C2 => n30645, ZN => n7623);
   U30605 : OAI222_X1 port map( A1 => n40766, A2 => n39897, B1 => n41150, B2 =>
                           n39890, C1 => n39883, C2 => n30644, ZN => n7622);
   U30606 : OAI222_X1 port map( A1 => n40772, A2 => n39897, B1 => n41156, B2 =>
                           n39890, C1 => n39883, C2 => n30643, ZN => n7621);
   U30607 : OAI222_X1 port map( A1 => n40778, A2 => n39897, B1 => n41162, B2 =>
                           n39890, C1 => n39883, C2 => n30642, ZN => n7620);
   U30608 : OAI222_X1 port map( A1 => n40784, A2 => n39897, B1 => n41168, B2 =>
                           n39890, C1 => n39883, C2 => n30641, ZN => n7619);
   U30609 : OAI222_X1 port map( A1 => n40790, A2 => n39897, B1 => n41174, B2 =>
                           n39890, C1 => n39883, C2 => n30640, ZN => n7618);
   U30610 : OAI222_X1 port map( A1 => n40796, A2 => n39897, B1 => n41180, B2 =>
                           n39890, C1 => n39883, C2 => n30639, ZN => n7617);
   U30611 : OAI222_X1 port map( A1 => n40802, A2 => n39897, B1 => n41186, B2 =>
                           n39890, C1 => n39883, C2 => n30638, ZN => n7616);
   U30612 : OAI222_X1 port map( A1 => n40808, A2 => n39897, B1 => n41192, B2 =>
                           n39890, C1 => n39883, C2 => n30637, ZN => n7615);
   U30613 : OAI222_X1 port map( A1 => n40814, A2 => n39897, B1 => n41198, B2 =>
                           n39890, C1 => n39884, C2 => n30636, ZN => n7614);
   U30614 : OAI222_X1 port map( A1 => n40820, A2 => n39897, B1 => n41204, B2 =>
                           n39890, C1 => n39884, C2 => n30635, ZN => n7613);
   U30615 : OAI222_X1 port map( A1 => n40826, A2 => n39897, B1 => n41210, B2 =>
                           n39890, C1 => n39884, C2 => n30634, ZN => n7612);
   U30616 : OAI222_X1 port map( A1 => n40832, A2 => n39897, B1 => n41216, B2 =>
                           n39890, C1 => n39884, C2 => n30633, ZN => n7611);
   U30617 : OAI222_X1 port map( A1 => n40838, A2 => n39896, B1 => n41222, B2 =>
                           n39889, C1 => n39884, C2 => n30632, ZN => n7610);
   U30618 : OAI222_X1 port map( A1 => n40844, A2 => n39896, B1 => n41228, B2 =>
                           n39889, C1 => n39884, C2 => n30631, ZN => n7609);
   U30619 : OAI222_X1 port map( A1 => n40850, A2 => n39896, B1 => n41234, B2 =>
                           n39889, C1 => n39884, C2 => n30630, ZN => n7608);
   U30620 : OAI222_X1 port map( A1 => n40856, A2 => n39896, B1 => n41240, B2 =>
                           n39889, C1 => n39884, C2 => n30629, ZN => n7607);
   U30621 : OAI222_X1 port map( A1 => n40862, A2 => n39896, B1 => n41246, B2 =>
                           n39889, C1 => n39884, C2 => n30628, ZN => n7606);
   U30622 : OAI222_X1 port map( A1 => n40868, A2 => n39896, B1 => n41252, B2 =>
                           n39889, C1 => n39884, C2 => n30627, ZN => n7605);
   U30623 : OAI222_X1 port map( A1 => n40874, A2 => n39896, B1 => n41258, B2 =>
                           n39889, C1 => n39884, C2 => n30626, ZN => n7604);
   U30624 : OAI222_X1 port map( A1 => n40880, A2 => n39896, B1 => n41264, B2 =>
                           n39889, C1 => n39884, C2 => n30625, ZN => n7603);
   U30625 : OAI222_X1 port map( A1 => n40886, A2 => n39896, B1 => n41270, B2 =>
                           n39889, C1 => n39885, C2 => n30624, ZN => n7602);
   U30626 : OAI222_X1 port map( A1 => n40892, A2 => n39896, B1 => n41276, B2 =>
                           n39889, C1 => n39885, C2 => n30623, ZN => n7601);
   U30627 : OAI222_X1 port map( A1 => n40898, A2 => n39896, B1 => n41282, B2 =>
                           n39889, C1 => n39885, C2 => n30622, ZN => n7600);
   U30628 : OAI222_X1 port map( A1 => n40904, A2 => n39896, B1 => n41288, B2 =>
                           n39889, C1 => n39885, C2 => n30621, ZN => n7599);
   U30629 : OAI222_X1 port map( A1 => n40910, A2 => n39895, B1 => n41294, B2 =>
                           n39888, C1 => n39885, C2 => n30620, ZN => n7598);
   U30630 : OAI222_X1 port map( A1 => n40916, A2 => n39895, B1 => n41300, B2 =>
                           n39888, C1 => n39885, C2 => n30619, ZN => n7597);
   U30631 : OAI222_X1 port map( A1 => n40922, A2 => n39895, B1 => n41306, B2 =>
                           n39888, C1 => n39885, C2 => n30618, ZN => n7596);
   U30632 : OAI222_X1 port map( A1 => n40928, A2 => n39895, B1 => n41312, B2 =>
                           n39888, C1 => n39885, C2 => n30617, ZN => n7595);
   U30633 : OAI222_X1 port map( A1 => n40934, A2 => n39895, B1 => n41318, B2 =>
                           n39888, C1 => n39885, C2 => n30616, ZN => n7594);
   U30634 : OAI222_X1 port map( A1 => n40940, A2 => n39895, B1 => n41324, B2 =>
                           n39888, C1 => n39885, C2 => n30615, ZN => n7593);
   U30635 : OAI222_X1 port map( A1 => n40946, A2 => n39895, B1 => n41330, B2 =>
                           n39888, C1 => n39885, C2 => n30614, ZN => n7592);
   U30636 : OAI222_X1 port map( A1 => n40958, A2 => n39895, B1 => n41342, B2 =>
                           n39888, C1 => n39885, C2 => n30612, ZN => n7590);
   U30637 : OAI222_X1 port map( A1 => n40598, A2 => n39880, B1 => n40982, B2 =>
                           n39873, C1 => n39861, C2 => n30608, ZN => n7586);
   U30638 : OAI222_X1 port map( A1 => n40604, A2 => n39880, B1 => n40988, B2 =>
                           n39873, C1 => n39861, C2 => n30607, ZN => n7585);
   U30639 : OAI222_X1 port map( A1 => n40610, A2 => n39880, B1 => n40994, B2 =>
                           n39873, C1 => n39861, C2 => n30606, ZN => n7584);
   U30640 : OAI222_X1 port map( A1 => n40616, A2 => n39880, B1 => n41000, B2 =>
                           n39873, C1 => n39861, C2 => n30605, ZN => n7583);
   U30641 : OAI222_X1 port map( A1 => n40622, A2 => n39879, B1 => n41006, B2 =>
                           n39872, C1 => n39861, C2 => n30604, ZN => n7582);
   U30642 : OAI222_X1 port map( A1 => n40628, A2 => n39879, B1 => n41012, B2 =>
                           n39872, C1 => n39861, C2 => n30603, ZN => n7581);
   U30643 : OAI222_X1 port map( A1 => n40634, A2 => n39879, B1 => n41018, B2 =>
                           n39872, C1 => n39861, C2 => n30602, ZN => n7580);
   U30644 : OAI222_X1 port map( A1 => n40640, A2 => n39879, B1 => n41024, B2 =>
                           n39872, C1 => n39861, C2 => n30601, ZN => n7579);
   U30645 : OAI222_X1 port map( A1 => n40646, A2 => n39879, B1 => n41030, B2 =>
                           n39872, C1 => n39861, C2 => n30600, ZN => n7578);
   U30646 : OAI222_X1 port map( A1 => n40652, A2 => n39879, B1 => n41036, B2 =>
                           n39872, C1 => n39861, C2 => n30599, ZN => n7577);
   U30647 : OAI222_X1 port map( A1 => n40658, A2 => n39879, B1 => n41042, B2 =>
                           n39872, C1 => n39861, C2 => n30598, ZN => n7576);
   U30648 : OAI222_X1 port map( A1 => n40664, A2 => n39879, B1 => n41048, B2 =>
                           n39872, C1 => n39861, C2 => n30597, ZN => n7575);
   U30649 : OAI222_X1 port map( A1 => n40670, A2 => n39879, B1 => n41054, B2 =>
                           n39872, C1 => n39862, C2 => n30596, ZN => n7574);
   U30650 : OAI222_X1 port map( A1 => n40676, A2 => n39879, B1 => n41060, B2 =>
                           n39872, C1 => n39862, C2 => n30595, ZN => n7573);
   U30651 : OAI222_X1 port map( A1 => n40682, A2 => n39879, B1 => n41066, B2 =>
                           n39872, C1 => n39862, C2 => n30594, ZN => n7572);
   U30652 : OAI222_X1 port map( A1 => n40688, A2 => n39879, B1 => n41072, B2 =>
                           n39872, C1 => n39863, C2 => n30593, ZN => n7571);
   U30653 : OAI222_X1 port map( A1 => n40694, A2 => n39878, B1 => n41078, B2 =>
                           n39871, C1 => n39862, C2 => n30592, ZN => n7570);
   U30654 : OAI222_X1 port map( A1 => n40700, A2 => n39878, B1 => n41084, B2 =>
                           n39871, C1 => n39862, C2 => n30591, ZN => n7569);
   U30655 : OAI222_X1 port map( A1 => n40706, A2 => n39878, B1 => n41090, B2 =>
                           n39871, C1 => n39862, C2 => n30590, ZN => n7568);
   U30656 : OAI222_X1 port map( A1 => n40712, A2 => n39878, B1 => n41096, B2 =>
                           n39871, C1 => n39862, C2 => n30589, ZN => n7567);
   U30657 : OAI222_X1 port map( A1 => n40718, A2 => n39878, B1 => n41102, B2 =>
                           n39871, C1 => n39862, C2 => n30588, ZN => n7566);
   U30658 : OAI222_X1 port map( A1 => n40724, A2 => n39878, B1 => n41108, B2 =>
                           n39871, C1 => n39862, C2 => n30587, ZN => n7565);
   U30659 : OAI222_X1 port map( A1 => n40730, A2 => n39878, B1 => n41114, B2 =>
                           n39871, C1 => n39862, C2 => n30586, ZN => n7564);
   U30660 : OAI222_X1 port map( A1 => n40736, A2 => n39878, B1 => n41120, B2 =>
                           n39871, C1 => n39862, C2 => n30585, ZN => n7563);
   U30661 : OAI222_X1 port map( A1 => n40742, A2 => n39878, B1 => n41126, B2 =>
                           n39871, C1 => n39862, C2 => n30584, ZN => n7562);
   U30662 : OAI222_X1 port map( A1 => n40748, A2 => n39878, B1 => n41132, B2 =>
                           n39871, C1 => n39863, C2 => n30583, ZN => n7561);
   U30663 : OAI222_X1 port map( A1 => n40754, A2 => n39878, B1 => n41138, B2 =>
                           n39871, C1 => n39863, C2 => n30582, ZN => n7560);
   U30664 : OAI222_X1 port map( A1 => n40760, A2 => n39878, B1 => n41144, B2 =>
                           n39871, C1 => n39863, C2 => n30581, ZN => n7559);
   U30665 : OAI222_X1 port map( A1 => n40766, A2 => n39877, B1 => n41150, B2 =>
                           n39870, C1 => n39863, C2 => n30580, ZN => n7558);
   U30666 : OAI222_X1 port map( A1 => n40772, A2 => n39877, B1 => n41156, B2 =>
                           n39870, C1 => n39863, C2 => n30579, ZN => n7557);
   U30667 : OAI222_X1 port map( A1 => n40778, A2 => n39877, B1 => n41162, B2 =>
                           n39870, C1 => n39863, C2 => n30578, ZN => n7556);
   U30668 : OAI222_X1 port map( A1 => n40784, A2 => n39877, B1 => n41168, B2 =>
                           n39870, C1 => n39863, C2 => n30577, ZN => n7555);
   U30669 : OAI222_X1 port map( A1 => n40790, A2 => n39877, B1 => n41174, B2 =>
                           n39870, C1 => n39863, C2 => n30576, ZN => n7554);
   U30670 : OAI222_X1 port map( A1 => n40796, A2 => n39877, B1 => n41180, B2 =>
                           n39870, C1 => n39863, C2 => n30575, ZN => n7553);
   U30671 : OAI222_X1 port map( A1 => n40802, A2 => n39877, B1 => n41186, B2 =>
                           n39870, C1 => n39863, C2 => n30574, ZN => n7552);
   U30672 : OAI222_X1 port map( A1 => n40808, A2 => n39877, B1 => n41192, B2 =>
                           n39870, C1 => n39863, C2 => n30573, ZN => n7551);
   U30673 : OAI222_X1 port map( A1 => n40814, A2 => n39877, B1 => n41198, B2 =>
                           n39870, C1 => n39864, C2 => n30572, ZN => n7550);
   U30674 : OAI222_X1 port map( A1 => n40820, A2 => n39877, B1 => n41204, B2 =>
                           n39870, C1 => n39864, C2 => n30571, ZN => n7549);
   U30675 : OAI222_X1 port map( A1 => n40826, A2 => n39877, B1 => n41210, B2 =>
                           n39870, C1 => n39864, C2 => n30570, ZN => n7548);
   U30676 : OAI222_X1 port map( A1 => n40832, A2 => n39877, B1 => n41216, B2 =>
                           n39870, C1 => n39864, C2 => n30569, ZN => n7547);
   U30677 : OAI222_X1 port map( A1 => n40838, A2 => n39876, B1 => n41222, B2 =>
                           n39869, C1 => n39864, C2 => n30568, ZN => n7546);
   U30678 : OAI222_X1 port map( A1 => n40844, A2 => n39876, B1 => n41228, B2 =>
                           n39869, C1 => n39864, C2 => n30567, ZN => n7545);
   U30679 : OAI222_X1 port map( A1 => n40850, A2 => n39876, B1 => n41234, B2 =>
                           n39869, C1 => n39864, C2 => n30566, ZN => n7544);
   U30680 : OAI222_X1 port map( A1 => n40856, A2 => n39876, B1 => n41240, B2 =>
                           n39869, C1 => n39864, C2 => n30565, ZN => n7543);
   U30681 : OAI222_X1 port map( A1 => n40862, A2 => n39876, B1 => n41246, B2 =>
                           n39869, C1 => n39864, C2 => n30564, ZN => n7542);
   U30682 : OAI222_X1 port map( A1 => n40868, A2 => n39876, B1 => n41252, B2 =>
                           n39869, C1 => n39864, C2 => n30563, ZN => n7541);
   U30683 : OAI222_X1 port map( A1 => n40874, A2 => n39876, B1 => n41258, B2 =>
                           n39869, C1 => n39864, C2 => n30562, ZN => n7540);
   U30684 : OAI222_X1 port map( A1 => n40880, A2 => n39876, B1 => n41264, B2 =>
                           n39869, C1 => n39864, C2 => n30561, ZN => n7539);
   U30685 : OAI222_X1 port map( A1 => n40886, A2 => n39876, B1 => n41270, B2 =>
                           n39869, C1 => n39865, C2 => n30560, ZN => n7538);
   U30686 : OAI222_X1 port map( A1 => n40892, A2 => n39876, B1 => n41276, B2 =>
                           n39869, C1 => n39865, C2 => n30559, ZN => n7537);
   U30687 : OAI222_X1 port map( A1 => n40898, A2 => n39876, B1 => n41282, B2 =>
                           n39869, C1 => n39865, C2 => n30558, ZN => n7536);
   U30688 : OAI222_X1 port map( A1 => n40904, A2 => n39876, B1 => n41288, B2 =>
                           n39869, C1 => n39865, C2 => n30557, ZN => n7535);
   U30689 : OAI222_X1 port map( A1 => n40910, A2 => n39875, B1 => n41294, B2 =>
                           n39868, C1 => n39865, C2 => n30556, ZN => n7534);
   U30690 : OAI222_X1 port map( A1 => n40916, A2 => n39875, B1 => n41300, B2 =>
                           n39868, C1 => n39865, C2 => n30555, ZN => n7533);
   U30691 : OAI222_X1 port map( A1 => n40922, A2 => n39875, B1 => n41306, B2 =>
                           n39868, C1 => n39865, C2 => n30554, ZN => n7532);
   U30692 : OAI222_X1 port map( A1 => n40928, A2 => n39875, B1 => n41312, B2 =>
                           n39868, C1 => n39865, C2 => n30553, ZN => n7531);
   U30693 : OAI222_X1 port map( A1 => n40934, A2 => n39875, B1 => n41318, B2 =>
                           n39868, C1 => n39865, C2 => n30552, ZN => n7530);
   U30694 : OAI222_X1 port map( A1 => n40940, A2 => n39875, B1 => n41324, B2 =>
                           n39868, C1 => n39865, C2 => n30551, ZN => n7529);
   U30695 : OAI222_X1 port map( A1 => n40946, A2 => n39875, B1 => n41330, B2 =>
                           n39868, C1 => n39865, C2 => n30550, ZN => n7528);
   U30696 : OAI222_X1 port map( A1 => n40958, A2 => n39875, B1 => n41342, B2 =>
                           n39868, C1 => n39865, C2 => n30548, ZN => n7526);
   U30697 : OAI222_X1 port map( A1 => n40598, A2 => n39860, B1 => n40982, B2 =>
                           n39853, C1 => n39841, C2 => n30544, ZN => n7522);
   U30698 : OAI222_X1 port map( A1 => n40604, A2 => n39860, B1 => n40988, B2 =>
                           n39853, C1 => n39841, C2 => n30543, ZN => n7521);
   U30699 : OAI222_X1 port map( A1 => n40610, A2 => n39860, B1 => n40994, B2 =>
                           n39853, C1 => n39841, C2 => n30542, ZN => n7520);
   U30700 : OAI222_X1 port map( A1 => n40616, A2 => n39860, B1 => n41000, B2 =>
                           n39853, C1 => n39841, C2 => n30541, ZN => n7519);
   U30701 : OAI222_X1 port map( A1 => n40622, A2 => n39859, B1 => n41006, B2 =>
                           n39852, C1 => n39841, C2 => n30540, ZN => n7518);
   U30702 : OAI222_X1 port map( A1 => n40628, A2 => n39859, B1 => n41012, B2 =>
                           n39852, C1 => n39841, C2 => n30539, ZN => n7517);
   U30703 : OAI222_X1 port map( A1 => n40634, A2 => n39859, B1 => n41018, B2 =>
                           n39852, C1 => n39841, C2 => n30538, ZN => n7516);
   U30704 : OAI222_X1 port map( A1 => n40640, A2 => n39859, B1 => n41024, B2 =>
                           n39852, C1 => n39841, C2 => n30537, ZN => n7515);
   U30705 : OAI222_X1 port map( A1 => n40646, A2 => n39859, B1 => n41030, B2 =>
                           n39852, C1 => n39841, C2 => n30536, ZN => n7514);
   U30706 : OAI222_X1 port map( A1 => n40652, A2 => n39859, B1 => n41036, B2 =>
                           n39852, C1 => n39841, C2 => n30535, ZN => n7513);
   U30707 : OAI222_X1 port map( A1 => n40658, A2 => n39859, B1 => n41042, B2 =>
                           n39852, C1 => n39841, C2 => n30534, ZN => n7512);
   U30708 : OAI222_X1 port map( A1 => n40664, A2 => n39859, B1 => n41048, B2 =>
                           n39852, C1 => n39841, C2 => n30533, ZN => n7511);
   U30709 : OAI222_X1 port map( A1 => n40670, A2 => n39859, B1 => n41054, B2 =>
                           n39852, C1 => n39842, C2 => n30532, ZN => n7510);
   U30710 : OAI222_X1 port map( A1 => n40676, A2 => n39859, B1 => n41060, B2 =>
                           n39852, C1 => n39842, C2 => n30531, ZN => n7509);
   U30711 : OAI222_X1 port map( A1 => n40682, A2 => n39859, B1 => n41066, B2 =>
                           n39852, C1 => n39842, C2 => n30530, ZN => n7508);
   U30712 : OAI222_X1 port map( A1 => n40688, A2 => n39859, B1 => n41072, B2 =>
                           n39852, C1 => n39843, C2 => n30529, ZN => n7507);
   U30713 : OAI222_X1 port map( A1 => n40694, A2 => n39858, B1 => n41078, B2 =>
                           n39851, C1 => n39842, C2 => n30528, ZN => n7506);
   U30714 : OAI222_X1 port map( A1 => n40700, A2 => n39858, B1 => n41084, B2 =>
                           n39851, C1 => n39842, C2 => n30527, ZN => n7505);
   U30715 : OAI222_X1 port map( A1 => n40706, A2 => n39858, B1 => n41090, B2 =>
                           n39851, C1 => n39842, C2 => n30526, ZN => n7504);
   U30716 : OAI222_X1 port map( A1 => n40712, A2 => n39858, B1 => n41096, B2 =>
                           n39851, C1 => n39842, C2 => n30525, ZN => n7503);
   U30717 : OAI222_X1 port map( A1 => n40718, A2 => n39858, B1 => n41102, B2 =>
                           n39851, C1 => n39842, C2 => n30524, ZN => n7502);
   U30718 : OAI222_X1 port map( A1 => n40724, A2 => n39858, B1 => n41108, B2 =>
                           n39851, C1 => n39842, C2 => n30523, ZN => n7501);
   U30719 : OAI222_X1 port map( A1 => n40730, A2 => n39858, B1 => n41114, B2 =>
                           n39851, C1 => n39842, C2 => n30522, ZN => n7500);
   U30720 : OAI222_X1 port map( A1 => n40736, A2 => n39858, B1 => n41120, B2 =>
                           n39851, C1 => n39842, C2 => n30521, ZN => n7499);
   U30721 : OAI222_X1 port map( A1 => n40742, A2 => n39858, B1 => n41126, B2 =>
                           n39851, C1 => n39842, C2 => n30520, ZN => n7498);
   U30722 : OAI222_X1 port map( A1 => n40748, A2 => n39858, B1 => n41132, B2 =>
                           n39851, C1 => n39843, C2 => n30519, ZN => n7497);
   U30723 : OAI222_X1 port map( A1 => n40754, A2 => n39858, B1 => n41138, B2 =>
                           n39851, C1 => n39843, C2 => n30518, ZN => n7496);
   U30724 : OAI222_X1 port map( A1 => n40760, A2 => n39858, B1 => n41144, B2 =>
                           n39851, C1 => n39843, C2 => n30517, ZN => n7495);
   U30725 : OAI222_X1 port map( A1 => n40766, A2 => n39857, B1 => n41150, B2 =>
                           n39850, C1 => n39843, C2 => n30516, ZN => n7494);
   U30726 : OAI222_X1 port map( A1 => n40772, A2 => n39857, B1 => n41156, B2 =>
                           n39850, C1 => n39843, C2 => n30515, ZN => n7493);
   U30727 : OAI222_X1 port map( A1 => n40778, A2 => n39857, B1 => n41162, B2 =>
                           n39850, C1 => n39843, C2 => n30514, ZN => n7492);
   U30728 : OAI222_X1 port map( A1 => n40784, A2 => n39857, B1 => n41168, B2 =>
                           n39850, C1 => n39843, C2 => n30513, ZN => n7491);
   U30729 : OAI222_X1 port map( A1 => n40790, A2 => n39857, B1 => n41174, B2 =>
                           n39850, C1 => n39843, C2 => n30512, ZN => n7490);
   U30730 : OAI222_X1 port map( A1 => n40796, A2 => n39857, B1 => n41180, B2 =>
                           n39850, C1 => n39843, C2 => n30511, ZN => n7489);
   U30731 : OAI222_X1 port map( A1 => n40802, A2 => n39857, B1 => n41186, B2 =>
                           n39850, C1 => n39843, C2 => n30510, ZN => n7488);
   U30732 : OAI222_X1 port map( A1 => n40808, A2 => n39857, B1 => n41192, B2 =>
                           n39850, C1 => n39843, C2 => n30509, ZN => n7487);
   U30733 : OAI222_X1 port map( A1 => n40814, A2 => n39857, B1 => n41198, B2 =>
                           n39850, C1 => n39844, C2 => n30508, ZN => n7486);
   U30734 : OAI222_X1 port map( A1 => n40820, A2 => n39857, B1 => n41204, B2 =>
                           n39850, C1 => n39844, C2 => n30507, ZN => n7485);
   U30735 : OAI222_X1 port map( A1 => n40826, A2 => n39857, B1 => n41210, B2 =>
                           n39850, C1 => n39844, C2 => n30506, ZN => n7484);
   U30736 : OAI222_X1 port map( A1 => n40832, A2 => n39857, B1 => n41216, B2 =>
                           n39850, C1 => n39844, C2 => n30505, ZN => n7483);
   U30737 : OAI222_X1 port map( A1 => n40838, A2 => n39856, B1 => n41222, B2 =>
                           n39849, C1 => n39844, C2 => n30504, ZN => n7482);
   U30738 : OAI222_X1 port map( A1 => n40844, A2 => n39856, B1 => n41228, B2 =>
                           n39849, C1 => n39844, C2 => n30503, ZN => n7481);
   U30739 : OAI222_X1 port map( A1 => n40850, A2 => n39856, B1 => n41234, B2 =>
                           n39849, C1 => n39844, C2 => n30502, ZN => n7480);
   U30740 : OAI222_X1 port map( A1 => n40856, A2 => n39856, B1 => n41240, B2 =>
                           n39849, C1 => n39844, C2 => n30501, ZN => n7479);
   U30741 : OAI222_X1 port map( A1 => n40862, A2 => n39856, B1 => n41246, B2 =>
                           n39849, C1 => n39844, C2 => n30500, ZN => n7478);
   U30742 : OAI222_X1 port map( A1 => n40868, A2 => n39856, B1 => n41252, B2 =>
                           n39849, C1 => n39844, C2 => n30499, ZN => n7477);
   U30743 : OAI222_X1 port map( A1 => n40874, A2 => n39856, B1 => n41258, B2 =>
                           n39849, C1 => n39844, C2 => n30498, ZN => n7476);
   U30744 : OAI222_X1 port map( A1 => n40880, A2 => n39856, B1 => n41264, B2 =>
                           n39849, C1 => n39844, C2 => n30497, ZN => n7475);
   U30745 : OAI222_X1 port map( A1 => n40886, A2 => n39856, B1 => n41270, B2 =>
                           n39849, C1 => n39845, C2 => n30496, ZN => n7474);
   U30746 : OAI222_X1 port map( A1 => n40892, A2 => n39856, B1 => n41276, B2 =>
                           n39849, C1 => n39845, C2 => n30495, ZN => n7473);
   U30747 : OAI222_X1 port map( A1 => n40898, A2 => n39856, B1 => n41282, B2 =>
                           n39849, C1 => n39845, C2 => n30494, ZN => n7472);
   U30748 : OAI222_X1 port map( A1 => n40904, A2 => n39856, B1 => n41288, B2 =>
                           n39849, C1 => n39845, C2 => n30493, ZN => n7471);
   U30749 : OAI222_X1 port map( A1 => n40910, A2 => n39855, B1 => n41294, B2 =>
                           n39848, C1 => n39845, C2 => n30492, ZN => n7470);
   U30750 : OAI222_X1 port map( A1 => n40916, A2 => n39855, B1 => n41300, B2 =>
                           n39848, C1 => n39845, C2 => n30491, ZN => n7469);
   U30751 : OAI222_X1 port map( A1 => n40922, A2 => n39855, B1 => n41306, B2 =>
                           n39848, C1 => n39845, C2 => n30490, ZN => n7468);
   U30752 : OAI222_X1 port map( A1 => n40928, A2 => n39855, B1 => n41312, B2 =>
                           n39848, C1 => n39845, C2 => n30489, ZN => n7467);
   U30753 : OAI222_X1 port map( A1 => n40934, A2 => n39855, B1 => n41318, B2 =>
                           n39848, C1 => n39845, C2 => n30488, ZN => n7466);
   U30754 : OAI222_X1 port map( A1 => n40940, A2 => n39855, B1 => n41324, B2 =>
                           n39848, C1 => n39845, C2 => n30487, ZN => n7465);
   U30755 : OAI222_X1 port map( A1 => n40946, A2 => n39855, B1 => n41330, B2 =>
                           n39848, C1 => n39845, C2 => n30486, ZN => n7464);
   U30756 : OAI222_X1 port map( A1 => n40958, A2 => n39855, B1 => n41342, B2 =>
                           n39848, C1 => n39845, C2 => n30484, ZN => n7462);
   U30757 : AOI221_X1 port map( B1 => n39102, B2 => n33031, C1 => n39096, C2 =>
                           n32983, A => n37026, ZN => n37021);
   U30758 : OAI222_X1 port map( A1 => n30789, A2 => n39090, B1 => n30853, B2 =>
                           n39084, C1 => n30725, C2 => n39078, ZN => n37026);
   U30759 : AOI221_X1 port map( B1 => n39103, B2 => n33030, C1 => n39097, C2 =>
                           n32982, A => n37007, ZN => n37002);
   U30760 : OAI222_X1 port map( A1 => n30788, A2 => n39091, B1 => n30852, B2 =>
                           n39085, C1 => n30724, C2 => n39079, ZN => n37007);
   U30761 : AOI221_X1 port map( B1 => n39103, B2 => n33029, C1 => n39097, C2 =>
                           n32981, A => n36988, ZN => n36983);
   U30762 : OAI222_X1 port map( A1 => n30787, A2 => n39091, B1 => n30851, B2 =>
                           n39085, C1 => n30723, C2 => n39079, ZN => n36988);
   U30763 : AOI221_X1 port map( B1 => n39103, B2 => n33028, C1 => n39097, C2 =>
                           n32980, A => n36969, ZN => n36964);
   U30764 : OAI222_X1 port map( A1 => n30786, A2 => n39091, B1 => n30850, B2 =>
                           n39085, C1 => n30722, C2 => n39079, ZN => n36969);
   U30765 : AOI221_X1 port map( B1 => n39103, B2 => n33027, C1 => n39097, C2 =>
                           n32979, A => n36950, ZN => n36945);
   U30766 : OAI222_X1 port map( A1 => n30785, A2 => n39091, B1 => n30849, B2 =>
                           n39085, C1 => n30721, C2 => n39079, ZN => n36950);
   U30767 : AOI221_X1 port map( B1 => n39103, B2 => n33026, C1 => n39097, C2 =>
                           n32978, A => n36931, ZN => n36926);
   U30768 : OAI222_X1 port map( A1 => n30784, A2 => n39091, B1 => n30848, B2 =>
                           n39085, C1 => n30720, C2 => n39079, ZN => n36931);
   U30769 : AOI221_X1 port map( B1 => n39103, B2 => n33025, C1 => n39097, C2 =>
                           n32977, A => n36912, ZN => n36907);
   U30770 : OAI222_X1 port map( A1 => n30783, A2 => n39091, B1 => n30847, B2 =>
                           n39085, C1 => n30719, C2 => n39079, ZN => n36912);
   U30771 : AOI221_X1 port map( B1 => n39103, B2 => n33024, C1 => n39097, C2 =>
                           n32976, A => n36893, ZN => n36888);
   U30772 : OAI222_X1 port map( A1 => n30782, A2 => n39091, B1 => n30846, B2 =>
                           n39085, C1 => n30718, C2 => n39079, ZN => n36893);
   U30773 : AOI221_X1 port map( B1 => n39103, B2 => n33023, C1 => n39097, C2 =>
                           n32975, A => n36874, ZN => n36869);
   U30774 : OAI222_X1 port map( A1 => n30781, A2 => n39091, B1 => n30845, B2 =>
                           n39085, C1 => n30717, C2 => n39079, ZN => n36874);
   U30775 : AOI221_X1 port map( B1 => n39103, B2 => n33022, C1 => n39097, C2 =>
                           n32974, A => n36855, ZN => n36850);
   U30776 : OAI222_X1 port map( A1 => n30780, A2 => n39091, B1 => n30844, B2 =>
                           n39085, C1 => n30716, C2 => n39079, ZN => n36855);
   U30777 : AOI221_X1 port map( B1 => n39103, B2 => n33021, C1 => n39097, C2 =>
                           n32973, A => n36836, ZN => n36831);
   U30778 : OAI222_X1 port map( A1 => n30779, A2 => n39091, B1 => n30843, B2 =>
                           n39085, C1 => n30715, C2 => n39079, ZN => n36836);
   U30779 : AOI221_X1 port map( B1 => n39103, B2 => n33020, C1 => n39097, C2 =>
                           n32972, A => n36817, ZN => n36812);
   U30780 : OAI222_X1 port map( A1 => n30778, A2 => n39091, B1 => n30842, B2 =>
                           n39085, C1 => n30714, C2 => n39079, ZN => n36817);
   U30781 : AOI221_X1 port map( B1 => n39103, B2 => n33019, C1 => n39097, C2 =>
                           n32971, A => n36798, ZN => n36793);
   U30782 : OAI222_X1 port map( A1 => n30777, A2 => n39091, B1 => n30841, B2 =>
                           n39085, C1 => n30713, C2 => n39079, ZN => n36798);
   U30783 : AOI221_X1 port map( B1 => n39104, B2 => n33018, C1 => n39098, C2 =>
                           n32970, A => n36779, ZN => n36774);
   U30784 : OAI222_X1 port map( A1 => n30776, A2 => n39092, B1 => n30840, B2 =>
                           n39086, C1 => n30712, C2 => n39080, ZN => n36779);
   U30785 : AOI221_X1 port map( B1 => n39104, B2 => n33017, C1 => n39098, C2 =>
                           n32969, A => n36760, ZN => n36755);
   U30786 : OAI222_X1 port map( A1 => n30775, A2 => n39092, B1 => n30839, B2 =>
                           n39086, C1 => n30711, C2 => n39080, ZN => n36760);
   U30787 : AOI221_X1 port map( B1 => n39104, B2 => n33016, C1 => n39098, C2 =>
                           n32968, A => n36741, ZN => n36736);
   U30788 : OAI222_X1 port map( A1 => n30774, A2 => n39092, B1 => n30838, B2 =>
                           n39086, C1 => n30710, C2 => n39080, ZN => n36741);
   U30789 : AOI221_X1 port map( B1 => n39104, B2 => n33015, C1 => n39098, C2 =>
                           n32967, A => n36722, ZN => n36717);
   U30790 : OAI222_X1 port map( A1 => n30773, A2 => n39092, B1 => n30837, B2 =>
                           n39086, C1 => n30709, C2 => n39080, ZN => n36722);
   U30791 : AOI221_X1 port map( B1 => n39104, B2 => n33014, C1 => n39098, C2 =>
                           n32966, A => n36703, ZN => n36698);
   U30792 : OAI222_X1 port map( A1 => n30772, A2 => n39092, B1 => n30836, B2 =>
                           n39086, C1 => n30708, C2 => n39080, ZN => n36703);
   U30793 : AOI221_X1 port map( B1 => n39104, B2 => n33013, C1 => n39098, C2 =>
                           n32965, A => n36684, ZN => n36679);
   U30794 : OAI222_X1 port map( A1 => n30771, A2 => n39092, B1 => n30835, B2 =>
                           n39086, C1 => n30707, C2 => n39080, ZN => n36684);
   U30795 : AOI221_X1 port map( B1 => n39104, B2 => n33012, C1 => n39098, C2 =>
                           n32964, A => n36665, ZN => n36660);
   U30796 : OAI222_X1 port map( A1 => n30770, A2 => n39092, B1 => n30834, B2 =>
                           n39086, C1 => n30706, C2 => n39080, ZN => n36665);
   U30797 : AOI221_X1 port map( B1 => n39104, B2 => n33011, C1 => n39098, C2 =>
                           n32963, A => n36646, ZN => n36641);
   U30798 : OAI222_X1 port map( A1 => n30769, A2 => n39092, B1 => n30833, B2 =>
                           n39086, C1 => n30705, C2 => n39080, ZN => n36646);
   U30799 : AOI221_X1 port map( B1 => n39104, B2 => n33010, C1 => n39098, C2 =>
                           n32962, A => n36627, ZN => n36622);
   U30800 : OAI222_X1 port map( A1 => n30768, A2 => n39092, B1 => n30832, B2 =>
                           n39086, C1 => n30704, C2 => n39080, ZN => n36627);
   U30801 : AOI221_X1 port map( B1 => n39104, B2 => n33009, C1 => n39098, C2 =>
                           n32961, A => n36608, ZN => n36603);
   U30802 : OAI222_X1 port map( A1 => n30767, A2 => n39092, B1 => n30831, B2 =>
                           n39086, C1 => n30703, C2 => n39080, ZN => n36608);
   U30803 : AOI221_X1 port map( B1 => n39104, B2 => n33008, C1 => n39098, C2 =>
                           n32960, A => n36589, ZN => n36584);
   U30804 : OAI222_X1 port map( A1 => n30766, A2 => n39092, B1 => n30830, B2 =>
                           n39086, C1 => n30702, C2 => n39080, ZN => n36589);
   U30805 : AOI221_X1 port map( B1 => n39104, B2 => n33007, C1 => n39098, C2 =>
                           n32959, A => n36570, ZN => n36565);
   U30806 : OAI222_X1 port map( A1 => n30765, A2 => n39092, B1 => n30829, B2 =>
                           n39086, C1 => n30701, C2 => n39080, ZN => n36570);
   U30807 : AOI221_X1 port map( B1 => n39105, B2 => n33006, C1 => n39099, C2 =>
                           n32958, A => n36551, ZN => n36546);
   U30808 : OAI222_X1 port map( A1 => n30764, A2 => n39093, B1 => n30828, B2 =>
                           n39087, C1 => n30700, C2 => n39081, ZN => n36551);
   U30809 : AOI221_X1 port map( B1 => n39105, B2 => n33005, C1 => n39099, C2 =>
                           n32957, A => n36532, ZN => n36527);
   U30810 : OAI222_X1 port map( A1 => n30763, A2 => n39093, B1 => n30827, B2 =>
                           n39087, C1 => n30699, C2 => n39081, ZN => n36532);
   U30811 : AOI221_X1 port map( B1 => n39105, B2 => n33004, C1 => n39099, C2 =>
                           n32956, A => n36513, ZN => n36508);
   U30812 : OAI222_X1 port map( A1 => n30762, A2 => n39093, B1 => n30826, B2 =>
                           n39087, C1 => n30698, C2 => n39081, ZN => n36513);
   U30813 : AOI221_X1 port map( B1 => n39105, B2 => n33003, C1 => n39099, C2 =>
                           n32955, A => n36494, ZN => n36489);
   U30814 : OAI222_X1 port map( A1 => n30761, A2 => n39093, B1 => n30825, B2 =>
                           n39087, C1 => n30697, C2 => n39081, ZN => n36494);
   U30815 : AOI221_X1 port map( B1 => n39105, B2 => n33002, C1 => n39099, C2 =>
                           n32954, A => n36475, ZN => n36470);
   U30816 : OAI222_X1 port map( A1 => n30760, A2 => n39093, B1 => n30824, B2 =>
                           n39087, C1 => n30696, C2 => n39081, ZN => n36475);
   U30817 : AOI221_X1 port map( B1 => n39105, B2 => n33001, C1 => n39099, C2 =>
                           n32953, A => n36456, ZN => n36451);
   U30818 : OAI222_X1 port map( A1 => n30759, A2 => n39093, B1 => n30823, B2 =>
                           n39087, C1 => n30695, C2 => n39081, ZN => n36456);
   U30819 : AOI221_X1 port map( B1 => n39105, B2 => n33000, C1 => n39099, C2 =>
                           n32952, A => n36437, ZN => n36432);
   U30820 : OAI222_X1 port map( A1 => n30758, A2 => n39093, B1 => n30822, B2 =>
                           n39087, C1 => n30694, C2 => n39081, ZN => n36437);
   U30821 : AOI221_X1 port map( B1 => n39105, B2 => n32999, C1 => n39099, C2 =>
                           n32951, A => n36418, ZN => n36413);
   U30822 : OAI222_X1 port map( A1 => n30757, A2 => n39093, B1 => n30821, B2 =>
                           n39087, C1 => n30693, C2 => n39081, ZN => n36418);
   U30823 : AOI221_X1 port map( B1 => n39105, B2 => n32998, C1 => n39099, C2 =>
                           n32950, A => n36399, ZN => n36394);
   U30824 : OAI222_X1 port map( A1 => n30756, A2 => n39093, B1 => n30820, B2 =>
                           n39087, C1 => n30692, C2 => n39081, ZN => n36399);
   U30825 : AOI221_X1 port map( B1 => n39105, B2 => n32997, C1 => n39099, C2 =>
                           n32949, A => n36380, ZN => n36375);
   U30826 : OAI222_X1 port map( A1 => n30755, A2 => n39093, B1 => n30819, B2 =>
                           n39087, C1 => n30691, C2 => n39081, ZN => n36380);
   U30827 : AOI221_X1 port map( B1 => n39105, B2 => n32996, C1 => n39099, C2 =>
                           n32948, A => n36361, ZN => n36356);
   U30828 : OAI222_X1 port map( A1 => n30754, A2 => n39093, B1 => n30818, B2 =>
                           n39087, C1 => n30690, C2 => n39081, ZN => n36361);
   U30829 : AOI221_X1 port map( B1 => n39105, B2 => n32995, C1 => n39099, C2 =>
                           n32947, A => n36342, ZN => n36337);
   U30830 : OAI222_X1 port map( A1 => n30753, A2 => n39093, B1 => n30817, B2 =>
                           n39087, C1 => n30689, C2 => n39081, ZN => n36342);
   U30831 : AOI221_X1 port map( B1 => n39106, B2 => n32994, C1 => n39100, C2 =>
                           n32946, A => n36323, ZN => n36318);
   U30832 : OAI222_X1 port map( A1 => n30752, A2 => n39094, B1 => n30816, B2 =>
                           n39088, C1 => n30688, C2 => n39082, ZN => n36323);
   U30833 : AOI221_X1 port map( B1 => n39106, B2 => n32993, C1 => n39100, C2 =>
                           n32945, A => n36304, ZN => n36299);
   U30834 : OAI222_X1 port map( A1 => n30751, A2 => n39094, B1 => n30815, B2 =>
                           n39088, C1 => n30687, C2 => n39082, ZN => n36304);
   U30835 : AOI221_X1 port map( B1 => n39106, B2 => n32992, C1 => n39100, C2 =>
                           n32944, A => n36285, ZN => n36280);
   U30836 : OAI222_X1 port map( A1 => n30750, A2 => n39094, B1 => n30814, B2 =>
                           n39088, C1 => n30686, C2 => n39082, ZN => n36285);
   U30837 : AOI221_X1 port map( B1 => n39106, B2 => n32991, C1 => n39100, C2 =>
                           n32943, A => n36266, ZN => n36261);
   U30838 : OAI222_X1 port map( A1 => n30749, A2 => n39094, B1 => n30813, B2 =>
                           n39088, C1 => n30685, C2 => n39082, ZN => n36266);
   U30839 : AOI221_X1 port map( B1 => n39106, B2 => n33134, C1 => n39100, C2 =>
                           n33122, A => n36247, ZN => n36242);
   U30840 : OAI222_X1 port map( A1 => n30748, A2 => n39094, B1 => n30812, B2 =>
                           n39088, C1 => n30684, C2 => n39082, ZN => n36247);
   U30841 : AOI221_X1 port map( B1 => n39106, B2 => n33133, C1 => n39100, C2 =>
                           n33121, A => n36228, ZN => n36223);
   U30842 : OAI222_X1 port map( A1 => n30747, A2 => n39094, B1 => n30811, B2 =>
                           n39088, C1 => n30683, C2 => n39082, ZN => n36228);
   U30843 : AOI221_X1 port map( B1 => n39102, B2 => n32490, C1 => n39096, C2 =>
                           n32486, A => n37216, ZN => n37211);
   U30844 : OAI222_X1 port map( A1 => n30799, A2 => n39090, B1 => n30863, B2 =>
                           n39084, C1 => n30735, C2 => n39078, ZN => n37216);
   U30845 : AOI221_X1 port map( B1 => n39102, B2 => n32489, C1 => n39096, C2 =>
                           n32485, A => n37197, ZN => n37192);
   U30846 : OAI222_X1 port map( A1 => n30798, A2 => n39090, B1 => n30862, B2 =>
                           n39084, C1 => n30734, C2 => n39078, ZN => n37197);
   U30847 : AOI221_X1 port map( B1 => n39102, B2 => n32488, C1 => n39096, C2 =>
                           n32484, A => n37178, ZN => n37173);
   U30848 : OAI222_X1 port map( A1 => n30797, A2 => n39090, B1 => n30861, B2 =>
                           n39084, C1 => n30733, C2 => n39078, ZN => n37178);
   U30849 : AOI221_X1 port map( B1 => n39102, B2 => n33038, C1 => n39096, C2 =>
                           n32990, A => n37159, ZN => n37154);
   U30850 : OAI222_X1 port map( A1 => n30796, A2 => n39090, B1 => n30860, B2 =>
                           n39084, C1 => n30732, C2 => n39078, ZN => n37159);
   U30851 : AOI221_X1 port map( B1 => n39102, B2 => n33037, C1 => n39096, C2 =>
                           n32989, A => n37140, ZN => n37135);
   U30852 : OAI222_X1 port map( A1 => n30795, A2 => n39090, B1 => n30859, B2 =>
                           n39084, C1 => n30731, C2 => n39078, ZN => n37140);
   U30853 : AOI221_X1 port map( B1 => n39107, B2 => n33126, C1 => n39101, C2 =>
                           n33114, A => n36095, ZN => n36090);
   U30854 : OAI222_X1 port map( A1 => n30740, A2 => n39095, B1 => n30804, B2 =>
                           n39089, C1 => n30676, C2 => n39083, ZN => n36095);
   U30855 : AOI221_X1 port map( B1 => n39107, B2 => n33125, C1 => n39101, C2 =>
                           n33113, A => n36076, ZN => n36071);
   U30856 : OAI222_X1 port map( A1 => n30739, A2 => n39095, B1 => n30803, B2 =>
                           n39089, C1 => n30675, C2 => n39083, ZN => n36076);
   U30857 : AOI221_X1 port map( B1 => n39107, B2 => n33124, C1 => n39101, C2 =>
                           n33112, A => n36057, ZN => n36052);
   U30858 : OAI222_X1 port map( A1 => n30738, A2 => n39095, B1 => n30802, B2 =>
                           n39089, C1 => n30674, C2 => n39083, ZN => n36057);
   U30859 : AOI221_X1 port map( B1 => n39107, B2 => n33123, C1 => n39101, C2 =>
                           n33111, A => n36030, ZN => n36013);
   U30860 : OAI222_X1 port map( A1 => n30737, A2 => n39095, B1 => n30801, B2 =>
                           n39089, C1 => n30673, C2 => n39083, ZN => n36030);
   U30861 : AOI221_X1 port map( B1 => n39102, B2 => n32491, C1 => n39096, C2 =>
                           n32487, A => n37248, ZN => n37242);
   U30862 : OAI222_X1 port map( A1 => n30800, A2 => n39090, B1 => n30864, B2 =>
                           n39084, C1 => n30736, C2 => n39078, ZN => n37248);
   U30863 : AOI221_X1 port map( B1 => n39102, B2 => n33036, C1 => n39096, C2 =>
                           n32988, A => n37121, ZN => n37116);
   U30864 : OAI222_X1 port map( A1 => n30794, A2 => n39090, B1 => n30858, B2 =>
                           n39084, C1 => n30730, C2 => n39078, ZN => n37121);
   U30865 : AOI221_X1 port map( B1 => n39102, B2 => n33035, C1 => n39096, C2 =>
                           n32987, A => n37102, ZN => n37097);
   U30866 : OAI222_X1 port map( A1 => n30793, A2 => n39090, B1 => n30857, B2 =>
                           n39084, C1 => n30729, C2 => n39078, ZN => n37102);
   U30867 : AOI221_X1 port map( B1 => n39102, B2 => n33034, C1 => n39096, C2 =>
                           n32986, A => n37083, ZN => n37078);
   U30868 : OAI222_X1 port map( A1 => n30792, A2 => n39090, B1 => n30856, B2 =>
                           n39084, C1 => n30728, C2 => n39078, ZN => n37083);
   U30869 : AOI221_X1 port map( B1 => n39102, B2 => n33033, C1 => n39096, C2 =>
                           n32985, A => n37064, ZN => n37059);
   U30870 : OAI222_X1 port map( A1 => n30791, A2 => n39090, B1 => n30855, B2 =>
                           n39084, C1 => n30727, C2 => n39078, ZN => n37064);
   U30871 : AOI221_X1 port map( B1 => n39102, B2 => n33032, C1 => n39096, C2 =>
                           n32984, A => n37045, ZN => n37040);
   U30872 : OAI222_X1 port map( A1 => n30790, A2 => n39090, B1 => n30854, B2 =>
                           n39084, C1 => n30726, C2 => n39078, ZN => n37045);
   U30873 : AOI221_X1 port map( B1 => n39106, B2 => n33132, C1 => n39100, C2 =>
                           n33120, A => n36209, ZN => n36204);
   U30874 : OAI222_X1 port map( A1 => n30746, A2 => n39094, B1 => n30810, B2 =>
                           n39088, C1 => n30682, C2 => n39082, ZN => n36209);
   U30875 : AOI221_X1 port map( B1 => n39106, B2 => n33131, C1 => n39100, C2 =>
                           n33119, A => n36190, ZN => n36185);
   U30876 : OAI222_X1 port map( A1 => n30745, A2 => n39094, B1 => n30809, B2 =>
                           n39088, C1 => n30681, C2 => n39082, ZN => n36190);
   U30877 : AOI221_X1 port map( B1 => n39106, B2 => n33130, C1 => n39100, C2 =>
                           n33118, A => n36171, ZN => n36166);
   U30878 : OAI222_X1 port map( A1 => n30744, A2 => n39094, B1 => n30808, B2 =>
                           n39088, C1 => n30680, C2 => n39082, ZN => n36171);
   U30879 : AOI221_X1 port map( B1 => n39106, B2 => n33129, C1 => n39100, C2 =>
                           n33117, A => n36152, ZN => n36147);
   U30880 : OAI222_X1 port map( A1 => n30743, A2 => n39094, B1 => n30807, B2 =>
                           n39088, C1 => n30679, C2 => n39082, ZN => n36152);
   U30881 : AOI221_X1 port map( B1 => n39106, B2 => n33128, C1 => n39100, C2 =>
                           n33116, A => n36133, ZN => n36128);
   U30882 : OAI222_X1 port map( A1 => n30742, A2 => n39094, B1 => n30806, B2 =>
                           n39088, C1 => n30678, C2 => n39082, ZN => n36133);
   U30883 : AOI221_X1 port map( B1 => n39106, B2 => n33127, C1 => n39100, C2 =>
                           n33115, A => n36114, ZN => n36109);
   U30884 : OAI222_X1 port map( A1 => n30741, A2 => n39094, B1 => n30805, B2 =>
                           n39088, C1 => n30677, C2 => n39082, ZN => n36114);
   U30885 : AOI221_X1 port map( B1 => n39609, B2 => n32491, C1 => n39603, C2 =>
                           n32487, A => n33475, ZN => n33458);
   U30886 : OAI222_X1 port map( A1 => n30800, A2 => n39597, B1 => n30864, B2 =>
                           n39591, C1 => n30736, C2 => n39585, ZN => n33475);
   U30887 : AOI221_X1 port map( B1 => n39357, B2 => n32491, C1 => n39351, C2 =>
                           n32487, A => n34749, ZN => n34732);
   U30888 : OAI222_X1 port map( A1 => n30800, A2 => n39345, B1 => n30864, B2 =>
                           n39339, C1 => n30736, C2 => n39333, ZN => n34749);
   U30889 : AOI221_X1 port map( B1 => n39609, B2 => n32490, C1 => n39603, C2 =>
                           n32486, A => n33502, ZN => n33497);
   U30890 : OAI222_X1 port map( A1 => n30799, A2 => n39597, B1 => n30863, B2 =>
                           n39591, C1 => n30735, C2 => n39585, ZN => n33502);
   U30891 : AOI221_X1 port map( B1 => n39357, B2 => n32490, C1 => n39351, C2 =>
                           n32486, A => n34776, ZN => n34771);
   U30892 : OAI222_X1 port map( A1 => n30799, A2 => n39345, B1 => n30863, B2 =>
                           n39339, C1 => n30735, C2 => n39333, ZN => n34776);
   U30893 : AOI221_X1 port map( B1 => n39609, B2 => n32489, C1 => n39603, C2 =>
                           n32485, A => n33521, ZN => n33516);
   U30894 : OAI222_X1 port map( A1 => n30798, A2 => n39597, B1 => n30862, B2 =>
                           n39591, C1 => n30734, C2 => n39585, ZN => n33521);
   U30895 : AOI221_X1 port map( B1 => n39357, B2 => n32489, C1 => n39351, C2 =>
                           n32485, A => n34795, ZN => n34790);
   U30896 : OAI222_X1 port map( A1 => n30798, A2 => n39345, B1 => n30862, B2 =>
                           n39339, C1 => n30734, C2 => n39333, ZN => n34795);
   U30897 : AOI221_X1 port map( B1 => n39609, B2 => n32488, C1 => n39603, C2 =>
                           n32484, A => n33540, ZN => n33535);
   U30898 : OAI222_X1 port map( A1 => n30797, A2 => n39597, B1 => n30861, B2 =>
                           n39591, C1 => n30733, C2 => n39585, ZN => n33540);
   U30899 : AOI221_X1 port map( B1 => n39357, B2 => n32488, C1 => n39351, C2 =>
                           n32484, A => n34814, ZN => n34809);
   U30900 : OAI222_X1 port map( A1 => n30797, A2 => n39345, B1 => n30861, B2 =>
                           n39339, C1 => n30733, C2 => n39333, ZN => n34814);
   U30901 : AOI221_X1 port map( B1 => n39608, B2 => n33038, C1 => n39602, C2 =>
                           n32990, A => n33559, ZN => n33554);
   U30902 : OAI222_X1 port map( A1 => n30796, A2 => n39596, B1 => n30860, B2 =>
                           n39590, C1 => n30732, C2 => n39584, ZN => n33559);
   U30903 : AOI221_X1 port map( B1 => n39356, B2 => n33038, C1 => n39350, C2 =>
                           n32990, A => n34833, ZN => n34828);
   U30904 : OAI222_X1 port map( A1 => n30796, A2 => n39344, B1 => n30860, B2 =>
                           n39338, C1 => n30732, C2 => n39332, ZN => n34833);
   U30905 : AOI221_X1 port map( B1 => n39608, B2 => n33037, C1 => n39602, C2 =>
                           n32989, A => n33578, ZN => n33573);
   U30906 : OAI222_X1 port map( A1 => n30795, A2 => n39596, B1 => n30859, B2 =>
                           n39590, C1 => n30731, C2 => n39584, ZN => n33578);
   U30907 : AOI221_X1 port map( B1 => n39356, B2 => n33037, C1 => n39350, C2 =>
                           n32989, A => n34852, ZN => n34847);
   U30908 : OAI222_X1 port map( A1 => n30795, A2 => n39344, B1 => n30859, B2 =>
                           n39338, C1 => n30731, C2 => n39332, ZN => n34852);
   U30909 : AOI221_X1 port map( B1 => n39608, B2 => n33036, C1 => n39602, C2 =>
                           n32988, A => n33597, ZN => n33592);
   U30910 : OAI222_X1 port map( A1 => n30794, A2 => n39596, B1 => n30858, B2 =>
                           n39590, C1 => n30730, C2 => n39584, ZN => n33597);
   U30911 : AOI221_X1 port map( B1 => n39356, B2 => n33036, C1 => n39350, C2 =>
                           n32988, A => n34871, ZN => n34866);
   U30912 : OAI222_X1 port map( A1 => n30794, A2 => n39344, B1 => n30858, B2 =>
                           n39338, C1 => n30730, C2 => n39332, ZN => n34871);
   U30913 : AOI221_X1 port map( B1 => n39608, B2 => n33035, C1 => n39602, C2 =>
                           n32987, A => n33616, ZN => n33611);
   U30914 : OAI222_X1 port map( A1 => n30793, A2 => n39596, B1 => n30857, B2 =>
                           n39590, C1 => n30729, C2 => n39584, ZN => n33616);
   U30915 : AOI221_X1 port map( B1 => n39356, B2 => n33035, C1 => n39350, C2 =>
                           n32987, A => n34890, ZN => n34885);
   U30916 : OAI222_X1 port map( A1 => n30793, A2 => n39344, B1 => n30857, B2 =>
                           n39338, C1 => n30729, C2 => n39332, ZN => n34890);
   U30917 : AOI221_X1 port map( B1 => n39608, B2 => n33034, C1 => n39602, C2 =>
                           n32986, A => n33635, ZN => n33630);
   U30918 : OAI222_X1 port map( A1 => n30792, A2 => n39596, B1 => n30856, B2 =>
                           n39590, C1 => n30728, C2 => n39584, ZN => n33635);
   U30919 : AOI221_X1 port map( B1 => n39356, B2 => n33034, C1 => n39350, C2 =>
                           n32986, A => n34909, ZN => n34904);
   U30920 : OAI222_X1 port map( A1 => n30792, A2 => n39344, B1 => n30856, B2 =>
                           n39338, C1 => n30728, C2 => n39332, ZN => n34909);
   U30921 : AOI221_X1 port map( B1 => n39608, B2 => n33033, C1 => n39602, C2 =>
                           n32985, A => n33654, ZN => n33649);
   U30922 : OAI222_X1 port map( A1 => n30791, A2 => n39596, B1 => n30855, B2 =>
                           n39590, C1 => n30727, C2 => n39584, ZN => n33654);
   U30923 : AOI221_X1 port map( B1 => n39356, B2 => n33033, C1 => n39350, C2 =>
                           n32985, A => n34928, ZN => n34923);
   U30924 : OAI222_X1 port map( A1 => n30791, A2 => n39344, B1 => n30855, B2 =>
                           n39338, C1 => n30727, C2 => n39332, ZN => n34928);
   U30925 : AOI221_X1 port map( B1 => n39608, B2 => n33032, C1 => n39602, C2 =>
                           n32984, A => n33673, ZN => n33668);
   U30926 : OAI222_X1 port map( A1 => n30790, A2 => n39596, B1 => n30854, B2 =>
                           n39590, C1 => n30726, C2 => n39584, ZN => n33673);
   U30927 : AOI221_X1 port map( B1 => n39356, B2 => n33032, C1 => n39350, C2 =>
                           n32984, A => n34947, ZN => n34942);
   U30928 : OAI222_X1 port map( A1 => n30790, A2 => n39344, B1 => n30854, B2 =>
                           n39338, C1 => n30726, C2 => n39332, ZN => n34947);
   U30929 : AOI221_X1 port map( B1 => n39608, B2 => n33031, C1 => n39602, C2 =>
                           n32983, A => n33692, ZN => n33687);
   U30930 : OAI222_X1 port map( A1 => n30789, A2 => n39596, B1 => n30853, B2 =>
                           n39590, C1 => n30725, C2 => n39584, ZN => n33692);
   U30931 : AOI221_X1 port map( B1 => n39356, B2 => n33031, C1 => n39350, C2 =>
                           n32983, A => n34966, ZN => n34961);
   U30932 : OAI222_X1 port map( A1 => n30789, A2 => n39344, B1 => n30853, B2 =>
                           n39338, C1 => n30725, C2 => n39332, ZN => n34966);
   U30933 : AOI221_X1 port map( B1 => n39608, B2 => n33030, C1 => n39602, C2 =>
                           n32982, A => n33711, ZN => n33706);
   U30934 : OAI222_X1 port map( A1 => n30788, A2 => n39596, B1 => n30852, B2 =>
                           n39590, C1 => n30724, C2 => n39584, ZN => n33711);
   U30935 : AOI221_X1 port map( B1 => n39356, B2 => n33030, C1 => n39350, C2 =>
                           n32982, A => n34985, ZN => n34980);
   U30936 : OAI222_X1 port map( A1 => n30788, A2 => n39344, B1 => n30852, B2 =>
                           n39338, C1 => n30724, C2 => n39332, ZN => n34985);
   U30937 : AOI221_X1 port map( B1 => n39608, B2 => n33029, C1 => n39602, C2 =>
                           n32981, A => n33730, ZN => n33725);
   U30938 : OAI222_X1 port map( A1 => n30787, A2 => n39596, B1 => n30851, B2 =>
                           n39590, C1 => n30723, C2 => n39584, ZN => n33730);
   U30939 : AOI221_X1 port map( B1 => n39356, B2 => n33029, C1 => n39350, C2 =>
                           n32981, A => n35004, ZN => n34999);
   U30940 : OAI222_X1 port map( A1 => n30787, A2 => n39344, B1 => n30851, B2 =>
                           n39338, C1 => n30723, C2 => n39332, ZN => n35004);
   U30941 : AOI221_X1 port map( B1 => n39608, B2 => n33028, C1 => n39602, C2 =>
                           n32980, A => n33749, ZN => n33744);
   U30942 : OAI222_X1 port map( A1 => n30786, A2 => n39596, B1 => n30850, B2 =>
                           n39590, C1 => n30722, C2 => n39584, ZN => n33749);
   U30943 : AOI221_X1 port map( B1 => n39356, B2 => n33028, C1 => n39350, C2 =>
                           n32980, A => n35023, ZN => n35018);
   U30944 : OAI222_X1 port map( A1 => n30786, A2 => n39344, B1 => n30850, B2 =>
                           n39338, C1 => n30722, C2 => n39332, ZN => n35023);
   U30945 : AOI221_X1 port map( B1 => n39608, B2 => n33027, C1 => n39602, C2 =>
                           n32979, A => n33768, ZN => n33763);
   U30946 : OAI222_X1 port map( A1 => n30785, A2 => n39596, B1 => n30849, B2 =>
                           n39590, C1 => n30721, C2 => n39584, ZN => n33768);
   U30947 : AOI221_X1 port map( B1 => n39356, B2 => n33027, C1 => n39350, C2 =>
                           n32979, A => n35042, ZN => n35037);
   U30948 : OAI222_X1 port map( A1 => n30785, A2 => n39344, B1 => n30849, B2 =>
                           n39338, C1 => n30721, C2 => n39332, ZN => n35042);
   U30949 : AOI221_X1 port map( B1 => n39607, B2 => n33026, C1 => n39601, C2 =>
                           n32978, A => n33787, ZN => n33782);
   U30950 : OAI222_X1 port map( A1 => n30784, A2 => n39595, B1 => n30848, B2 =>
                           n39589, C1 => n30720, C2 => n39583, ZN => n33787);
   U30951 : AOI221_X1 port map( B1 => n39355, B2 => n33026, C1 => n39349, C2 =>
                           n32978, A => n35061, ZN => n35056);
   U30952 : OAI222_X1 port map( A1 => n30784, A2 => n39343, B1 => n30848, B2 =>
                           n39337, C1 => n30720, C2 => n39331, ZN => n35061);
   U30953 : AOI221_X1 port map( B1 => n39607, B2 => n33025, C1 => n39601, C2 =>
                           n32977, A => n33806, ZN => n33801);
   U30954 : OAI222_X1 port map( A1 => n30783, A2 => n39595, B1 => n30847, B2 =>
                           n39589, C1 => n30719, C2 => n39583, ZN => n33806);
   U30955 : AOI221_X1 port map( B1 => n39355, B2 => n33025, C1 => n39349, C2 =>
                           n32977, A => n35080, ZN => n35075);
   U30956 : OAI222_X1 port map( A1 => n30783, A2 => n39343, B1 => n30847, B2 =>
                           n39337, C1 => n30719, C2 => n39331, ZN => n35080);
   U30957 : AOI221_X1 port map( B1 => n39607, B2 => n33024, C1 => n39601, C2 =>
                           n32976, A => n33825, ZN => n33820);
   U30958 : OAI222_X1 port map( A1 => n30782, A2 => n39595, B1 => n30846, B2 =>
                           n39589, C1 => n30718, C2 => n39583, ZN => n33825);
   U30959 : AOI221_X1 port map( B1 => n39355, B2 => n33024, C1 => n39349, C2 =>
                           n32976, A => n35099, ZN => n35094);
   U30960 : OAI222_X1 port map( A1 => n30782, A2 => n39343, B1 => n30846, B2 =>
                           n39337, C1 => n30718, C2 => n39331, ZN => n35099);
   U30961 : AOI221_X1 port map( B1 => n39607, B2 => n33023, C1 => n39601, C2 =>
                           n32975, A => n33844, ZN => n33839);
   U30962 : OAI222_X1 port map( A1 => n30781, A2 => n39595, B1 => n30845, B2 =>
                           n39589, C1 => n30717, C2 => n39583, ZN => n33844);
   U30963 : AOI221_X1 port map( B1 => n39355, B2 => n33023, C1 => n39349, C2 =>
                           n32975, A => n35118, ZN => n35113);
   U30964 : OAI222_X1 port map( A1 => n30781, A2 => n39343, B1 => n30845, B2 =>
                           n39337, C1 => n30717, C2 => n39331, ZN => n35118);
   U30965 : AOI221_X1 port map( B1 => n39607, B2 => n33022, C1 => n39601, C2 =>
                           n32974, A => n33863, ZN => n33858);
   U30966 : OAI222_X1 port map( A1 => n30780, A2 => n39595, B1 => n30844, B2 =>
                           n39589, C1 => n30716, C2 => n39583, ZN => n33863);
   U30967 : AOI221_X1 port map( B1 => n39355, B2 => n33022, C1 => n39349, C2 =>
                           n32974, A => n35137, ZN => n35132);
   U30968 : OAI222_X1 port map( A1 => n30780, A2 => n39343, B1 => n30844, B2 =>
                           n39337, C1 => n30716, C2 => n39331, ZN => n35137);
   U30969 : AOI221_X1 port map( B1 => n39607, B2 => n33021, C1 => n39601, C2 =>
                           n32973, A => n33882, ZN => n33877);
   U30970 : OAI222_X1 port map( A1 => n30779, A2 => n39595, B1 => n30843, B2 =>
                           n39589, C1 => n30715, C2 => n39583, ZN => n33882);
   U30971 : AOI221_X1 port map( B1 => n39355, B2 => n33021, C1 => n39349, C2 =>
                           n32973, A => n35156, ZN => n35151);
   U30972 : OAI222_X1 port map( A1 => n30779, A2 => n39343, B1 => n30843, B2 =>
                           n39337, C1 => n30715, C2 => n39331, ZN => n35156);
   U30973 : AOI221_X1 port map( B1 => n39607, B2 => n33020, C1 => n39601, C2 =>
                           n32972, A => n33901, ZN => n33896);
   U30974 : OAI222_X1 port map( A1 => n30778, A2 => n39595, B1 => n30842, B2 =>
                           n39589, C1 => n30714, C2 => n39583, ZN => n33901);
   U30975 : AOI221_X1 port map( B1 => n39355, B2 => n33020, C1 => n39349, C2 =>
                           n32972, A => n35175, ZN => n35170);
   U30976 : OAI222_X1 port map( A1 => n30778, A2 => n39343, B1 => n30842, B2 =>
                           n39337, C1 => n30714, C2 => n39331, ZN => n35175);
   U30977 : AOI221_X1 port map( B1 => n39607, B2 => n33019, C1 => n39601, C2 =>
                           n32971, A => n33920, ZN => n33915);
   U30978 : OAI222_X1 port map( A1 => n30777, A2 => n39595, B1 => n30841, B2 =>
                           n39589, C1 => n30713, C2 => n39583, ZN => n33920);
   U30979 : AOI221_X1 port map( B1 => n39355, B2 => n33019, C1 => n39349, C2 =>
                           n32971, A => n35194, ZN => n35189);
   U30980 : OAI222_X1 port map( A1 => n30777, A2 => n39343, B1 => n30841, B2 =>
                           n39337, C1 => n30713, C2 => n39331, ZN => n35194);
   U30981 : AOI221_X1 port map( B1 => n39607, B2 => n33018, C1 => n39601, C2 =>
                           n32970, A => n33939, ZN => n33934);
   U30982 : OAI222_X1 port map( A1 => n30776, A2 => n39595, B1 => n30840, B2 =>
                           n39589, C1 => n30712, C2 => n39583, ZN => n33939);
   U30983 : AOI221_X1 port map( B1 => n39355, B2 => n33018, C1 => n39349, C2 =>
                           n32970, A => n35213, ZN => n35208);
   U30984 : OAI222_X1 port map( A1 => n30776, A2 => n39343, B1 => n30840, B2 =>
                           n39337, C1 => n30712, C2 => n39331, ZN => n35213);
   U30985 : AOI221_X1 port map( B1 => n39607, B2 => n33017, C1 => n39601, C2 =>
                           n32969, A => n33958, ZN => n33953);
   U30986 : OAI222_X1 port map( A1 => n30775, A2 => n39595, B1 => n30839, B2 =>
                           n39589, C1 => n30711, C2 => n39583, ZN => n33958);
   U30987 : AOI221_X1 port map( B1 => n39355, B2 => n33017, C1 => n39349, C2 =>
                           n32969, A => n35232, ZN => n35227);
   U30988 : OAI222_X1 port map( A1 => n30775, A2 => n39343, B1 => n30839, B2 =>
                           n39337, C1 => n30711, C2 => n39331, ZN => n35232);
   U30989 : AOI221_X1 port map( B1 => n39607, B2 => n33016, C1 => n39601, C2 =>
                           n32968, A => n33977, ZN => n33972);
   U30990 : OAI222_X1 port map( A1 => n30774, A2 => n39595, B1 => n30838, B2 =>
                           n39589, C1 => n30710, C2 => n39583, ZN => n33977);
   U30991 : AOI221_X1 port map( B1 => n39355, B2 => n33016, C1 => n39349, C2 =>
                           n32968, A => n35251, ZN => n35246);
   U30992 : OAI222_X1 port map( A1 => n30774, A2 => n39343, B1 => n30838, B2 =>
                           n39337, C1 => n30710, C2 => n39331, ZN => n35251);
   U30993 : AOI221_X1 port map( B1 => n39607, B2 => n33015, C1 => n39601, C2 =>
                           n32967, A => n33996, ZN => n33991);
   U30994 : OAI222_X1 port map( A1 => n30773, A2 => n39595, B1 => n30837, B2 =>
                           n39589, C1 => n30709, C2 => n39583, ZN => n33996);
   U30995 : AOI221_X1 port map( B1 => n39355, B2 => n33015, C1 => n39349, C2 =>
                           n32967, A => n35270, ZN => n35265);
   U30996 : OAI222_X1 port map( A1 => n30773, A2 => n39343, B1 => n30837, B2 =>
                           n39337, C1 => n30709, C2 => n39331, ZN => n35270);
   U30997 : AOI221_X1 port map( B1 => n39606, B2 => n33014, C1 => n39600, C2 =>
                           n32966, A => n34015, ZN => n34010);
   U30998 : OAI222_X1 port map( A1 => n30772, A2 => n39594, B1 => n30836, B2 =>
                           n39588, C1 => n30708, C2 => n39582, ZN => n34015);
   U30999 : AOI221_X1 port map( B1 => n39354, B2 => n33014, C1 => n39348, C2 =>
                           n32966, A => n35289, ZN => n35284);
   U31000 : OAI222_X1 port map( A1 => n30772, A2 => n39342, B1 => n30836, B2 =>
                           n39336, C1 => n30708, C2 => n39330, ZN => n35289);
   U31001 : AOI221_X1 port map( B1 => n39606, B2 => n33013, C1 => n39600, C2 =>
                           n32965, A => n34034, ZN => n34029);
   U31002 : OAI222_X1 port map( A1 => n30771, A2 => n39594, B1 => n30835, B2 =>
                           n39588, C1 => n30707, C2 => n39582, ZN => n34034);
   U31003 : AOI221_X1 port map( B1 => n39354, B2 => n33013, C1 => n39348, C2 =>
                           n32965, A => n35308, ZN => n35303);
   U31004 : OAI222_X1 port map( A1 => n30771, A2 => n39342, B1 => n30835, B2 =>
                           n39336, C1 => n30707, C2 => n39330, ZN => n35308);
   U31005 : AOI221_X1 port map( B1 => n39606, B2 => n33012, C1 => n39600, C2 =>
                           n32964, A => n34053, ZN => n34048);
   U31006 : OAI222_X1 port map( A1 => n30770, A2 => n39594, B1 => n30834, B2 =>
                           n39588, C1 => n30706, C2 => n39582, ZN => n34053);
   U31007 : AOI221_X1 port map( B1 => n39354, B2 => n33012, C1 => n39348, C2 =>
                           n32964, A => n35327, ZN => n35322);
   U31008 : OAI222_X1 port map( A1 => n30770, A2 => n39342, B1 => n30834, B2 =>
                           n39336, C1 => n30706, C2 => n39330, ZN => n35327);
   U31009 : AOI221_X1 port map( B1 => n39606, B2 => n33011, C1 => n39600, C2 =>
                           n32963, A => n34072, ZN => n34067);
   U31010 : OAI222_X1 port map( A1 => n30769, A2 => n39594, B1 => n30833, B2 =>
                           n39588, C1 => n30705, C2 => n39582, ZN => n34072);
   U31011 : AOI221_X1 port map( B1 => n39354, B2 => n33011, C1 => n39348, C2 =>
                           n32963, A => n35346, ZN => n35341);
   U31012 : OAI222_X1 port map( A1 => n30769, A2 => n39342, B1 => n30833, B2 =>
                           n39336, C1 => n30705, C2 => n39330, ZN => n35346);
   U31013 : AOI221_X1 port map( B1 => n39606, B2 => n33010, C1 => n39600, C2 =>
                           n32962, A => n34091, ZN => n34086);
   U31014 : OAI222_X1 port map( A1 => n30768, A2 => n39594, B1 => n30832, B2 =>
                           n39588, C1 => n30704, C2 => n39582, ZN => n34091);
   U31015 : AOI221_X1 port map( B1 => n39354, B2 => n33010, C1 => n39348, C2 =>
                           n32962, A => n35365, ZN => n35360);
   U31016 : OAI222_X1 port map( A1 => n30768, A2 => n39342, B1 => n30832, B2 =>
                           n39336, C1 => n30704, C2 => n39330, ZN => n35365);
   U31017 : AOI221_X1 port map( B1 => n39606, B2 => n33009, C1 => n39600, C2 =>
                           n32961, A => n34110, ZN => n34105);
   U31018 : OAI222_X1 port map( A1 => n30767, A2 => n39594, B1 => n30831, B2 =>
                           n39588, C1 => n30703, C2 => n39582, ZN => n34110);
   U31019 : AOI221_X1 port map( B1 => n39354, B2 => n33009, C1 => n39348, C2 =>
                           n32961, A => n35384, ZN => n35379);
   U31020 : OAI222_X1 port map( A1 => n30767, A2 => n39342, B1 => n30831, B2 =>
                           n39336, C1 => n30703, C2 => n39330, ZN => n35384);
   U31021 : AOI221_X1 port map( B1 => n39606, B2 => n33008, C1 => n39600, C2 =>
                           n32960, A => n34129, ZN => n34124);
   U31022 : OAI222_X1 port map( A1 => n30766, A2 => n39594, B1 => n30830, B2 =>
                           n39588, C1 => n30702, C2 => n39582, ZN => n34129);
   U31023 : AOI221_X1 port map( B1 => n39354, B2 => n33008, C1 => n39348, C2 =>
                           n32960, A => n35403, ZN => n35398);
   U31024 : OAI222_X1 port map( A1 => n30766, A2 => n39342, B1 => n30830, B2 =>
                           n39336, C1 => n30702, C2 => n39330, ZN => n35403);
   U31025 : AOI221_X1 port map( B1 => n39606, B2 => n33007, C1 => n39600, C2 =>
                           n32959, A => n34148, ZN => n34143);
   U31026 : OAI222_X1 port map( A1 => n30765, A2 => n39594, B1 => n30829, B2 =>
                           n39588, C1 => n30701, C2 => n39582, ZN => n34148);
   U31027 : AOI221_X1 port map( B1 => n39354, B2 => n33007, C1 => n39348, C2 =>
                           n32959, A => n35422, ZN => n35417);
   U31028 : OAI222_X1 port map( A1 => n30765, A2 => n39342, B1 => n30829, B2 =>
                           n39336, C1 => n30701, C2 => n39330, ZN => n35422);
   U31029 : AOI221_X1 port map( B1 => n39606, B2 => n33006, C1 => n39600, C2 =>
                           n32958, A => n34167, ZN => n34162);
   U31030 : OAI222_X1 port map( A1 => n30764, A2 => n39594, B1 => n30828, B2 =>
                           n39588, C1 => n30700, C2 => n39582, ZN => n34167);
   U31031 : AOI221_X1 port map( B1 => n39354, B2 => n33006, C1 => n39348, C2 =>
                           n32958, A => n35441, ZN => n35436);
   U31032 : OAI222_X1 port map( A1 => n30764, A2 => n39342, B1 => n30828, B2 =>
                           n39336, C1 => n30700, C2 => n39330, ZN => n35441);
   U31033 : AOI221_X1 port map( B1 => n39606, B2 => n33005, C1 => n39600, C2 =>
                           n32957, A => n34186, ZN => n34181);
   U31034 : OAI222_X1 port map( A1 => n30763, A2 => n39594, B1 => n30827, B2 =>
                           n39588, C1 => n30699, C2 => n39582, ZN => n34186);
   U31035 : AOI221_X1 port map( B1 => n39354, B2 => n33005, C1 => n39348, C2 =>
                           n32957, A => n35460, ZN => n35455);
   U31036 : OAI222_X1 port map( A1 => n30763, A2 => n39342, B1 => n30827, B2 =>
                           n39336, C1 => n30699, C2 => n39330, ZN => n35460);
   U31037 : AOI221_X1 port map( B1 => n39606, B2 => n33004, C1 => n39600, C2 =>
                           n32956, A => n34205, ZN => n34200);
   U31038 : OAI222_X1 port map( A1 => n30762, A2 => n39594, B1 => n30826, B2 =>
                           n39588, C1 => n30698, C2 => n39582, ZN => n34205);
   U31039 : AOI221_X1 port map( B1 => n39354, B2 => n33004, C1 => n39348, C2 =>
                           n32956, A => n35479, ZN => n35474);
   U31040 : OAI222_X1 port map( A1 => n30762, A2 => n39342, B1 => n30826, B2 =>
                           n39336, C1 => n30698, C2 => n39330, ZN => n35479);
   U31041 : AOI221_X1 port map( B1 => n39606, B2 => n33003, C1 => n39600, C2 =>
                           n32955, A => n34224, ZN => n34219);
   U31042 : OAI222_X1 port map( A1 => n30761, A2 => n39594, B1 => n30825, B2 =>
                           n39588, C1 => n30697, C2 => n39582, ZN => n34224);
   U31043 : AOI221_X1 port map( B1 => n39354, B2 => n33003, C1 => n39348, C2 =>
                           n32955, A => n35498, ZN => n35493);
   U31044 : OAI222_X1 port map( A1 => n30761, A2 => n39342, B1 => n30825, B2 =>
                           n39336, C1 => n30697, C2 => n39330, ZN => n35498);
   U31045 : AOI221_X1 port map( B1 => n39605, B2 => n33002, C1 => n39599, C2 =>
                           n32954, A => n34243, ZN => n34238);
   U31046 : OAI222_X1 port map( A1 => n30760, A2 => n39593, B1 => n30824, B2 =>
                           n39587, C1 => n30696, C2 => n39581, ZN => n34243);
   U31047 : AOI221_X1 port map( B1 => n39353, B2 => n33002, C1 => n39347, C2 =>
                           n32954, A => n35517, ZN => n35512);
   U31048 : OAI222_X1 port map( A1 => n30760, A2 => n39341, B1 => n30824, B2 =>
                           n39335, C1 => n30696, C2 => n39329, ZN => n35517);
   U31049 : AOI221_X1 port map( B1 => n39605, B2 => n33001, C1 => n39599, C2 =>
                           n32953, A => n34262, ZN => n34257);
   U31050 : OAI222_X1 port map( A1 => n30759, A2 => n39593, B1 => n30823, B2 =>
                           n39587, C1 => n30695, C2 => n39581, ZN => n34262);
   U31051 : AOI221_X1 port map( B1 => n39353, B2 => n33001, C1 => n39347, C2 =>
                           n32953, A => n35536, ZN => n35531);
   U31052 : OAI222_X1 port map( A1 => n30759, A2 => n39341, B1 => n30823, B2 =>
                           n39335, C1 => n30695, C2 => n39329, ZN => n35536);
   U31053 : AOI221_X1 port map( B1 => n39605, B2 => n33000, C1 => n39599, C2 =>
                           n32952, A => n34281, ZN => n34276);
   U31054 : OAI222_X1 port map( A1 => n30758, A2 => n39593, B1 => n30822, B2 =>
                           n39587, C1 => n30694, C2 => n39581, ZN => n34281);
   U31055 : AOI221_X1 port map( B1 => n39353, B2 => n33000, C1 => n39347, C2 =>
                           n32952, A => n35555, ZN => n35550);
   U31056 : OAI222_X1 port map( A1 => n30758, A2 => n39341, B1 => n30822, B2 =>
                           n39335, C1 => n30694, C2 => n39329, ZN => n35555);
   U31057 : AOI221_X1 port map( B1 => n39605, B2 => n32999, C1 => n39599, C2 =>
                           n32951, A => n34300, ZN => n34295);
   U31058 : OAI222_X1 port map( A1 => n30757, A2 => n39593, B1 => n30821, B2 =>
                           n39587, C1 => n30693, C2 => n39581, ZN => n34300);
   U31059 : AOI221_X1 port map( B1 => n39353, B2 => n32999, C1 => n39347, C2 =>
                           n32951, A => n35574, ZN => n35569);
   U31060 : OAI222_X1 port map( A1 => n30757, A2 => n39341, B1 => n30821, B2 =>
                           n39335, C1 => n30693, C2 => n39329, ZN => n35574);
   U31061 : AOI221_X1 port map( B1 => n39605, B2 => n32998, C1 => n39599, C2 =>
                           n32950, A => n34319, ZN => n34314);
   U31062 : OAI222_X1 port map( A1 => n30756, A2 => n39593, B1 => n30820, B2 =>
                           n39587, C1 => n30692, C2 => n39581, ZN => n34319);
   U31063 : AOI221_X1 port map( B1 => n39353, B2 => n32998, C1 => n39347, C2 =>
                           n32950, A => n35593, ZN => n35588);
   U31064 : OAI222_X1 port map( A1 => n30756, A2 => n39341, B1 => n30820, B2 =>
                           n39335, C1 => n30692, C2 => n39329, ZN => n35593);
   U31065 : AOI221_X1 port map( B1 => n39605, B2 => n32997, C1 => n39599, C2 =>
                           n32949, A => n34338, ZN => n34333);
   U31066 : OAI222_X1 port map( A1 => n30755, A2 => n39593, B1 => n30819, B2 =>
                           n39587, C1 => n30691, C2 => n39581, ZN => n34338);
   U31067 : AOI221_X1 port map( B1 => n39353, B2 => n32997, C1 => n39347, C2 =>
                           n32949, A => n35612, ZN => n35607);
   U31068 : OAI222_X1 port map( A1 => n30755, A2 => n39341, B1 => n30819, B2 =>
                           n39335, C1 => n30691, C2 => n39329, ZN => n35612);
   U31069 : AOI221_X1 port map( B1 => n39605, B2 => n32996, C1 => n39599, C2 =>
                           n32948, A => n34357, ZN => n34352);
   U31070 : OAI222_X1 port map( A1 => n30754, A2 => n39593, B1 => n30818, B2 =>
                           n39587, C1 => n30690, C2 => n39581, ZN => n34357);
   U31071 : AOI221_X1 port map( B1 => n39353, B2 => n32996, C1 => n39347, C2 =>
                           n32948, A => n35631, ZN => n35626);
   U31072 : OAI222_X1 port map( A1 => n30754, A2 => n39341, B1 => n30818, B2 =>
                           n39335, C1 => n30690, C2 => n39329, ZN => n35631);
   U31073 : AOI221_X1 port map( B1 => n39605, B2 => n32995, C1 => n39599, C2 =>
                           n32947, A => n34376, ZN => n34371);
   U31074 : OAI222_X1 port map( A1 => n30753, A2 => n39593, B1 => n30817, B2 =>
                           n39587, C1 => n30689, C2 => n39581, ZN => n34376);
   U31075 : AOI221_X1 port map( B1 => n39353, B2 => n32995, C1 => n39347, C2 =>
                           n32947, A => n35650, ZN => n35645);
   U31076 : OAI222_X1 port map( A1 => n30753, A2 => n39341, B1 => n30817, B2 =>
                           n39335, C1 => n30689, C2 => n39329, ZN => n35650);
   U31077 : AOI221_X1 port map( B1 => n39605, B2 => n32994, C1 => n39599, C2 =>
                           n32946, A => n34395, ZN => n34390);
   U31078 : OAI222_X1 port map( A1 => n30752, A2 => n39593, B1 => n30816, B2 =>
                           n39587, C1 => n30688, C2 => n39581, ZN => n34395);
   U31079 : AOI221_X1 port map( B1 => n39353, B2 => n32994, C1 => n39347, C2 =>
                           n32946, A => n35669, ZN => n35664);
   U31080 : OAI222_X1 port map( A1 => n30752, A2 => n39341, B1 => n30816, B2 =>
                           n39335, C1 => n30688, C2 => n39329, ZN => n35669);
   U31081 : AOI221_X1 port map( B1 => n39605, B2 => n32993, C1 => n39599, C2 =>
                           n32945, A => n34414, ZN => n34409);
   U31082 : OAI222_X1 port map( A1 => n30751, A2 => n39593, B1 => n30815, B2 =>
                           n39587, C1 => n30687, C2 => n39581, ZN => n34414);
   U31083 : AOI221_X1 port map( B1 => n39353, B2 => n32993, C1 => n39347, C2 =>
                           n32945, A => n35688, ZN => n35683);
   U31084 : OAI222_X1 port map( A1 => n30751, A2 => n39341, B1 => n30815, B2 =>
                           n39335, C1 => n30687, C2 => n39329, ZN => n35688);
   U31085 : AOI221_X1 port map( B1 => n39605, B2 => n32992, C1 => n39599, C2 =>
                           n32944, A => n34433, ZN => n34428);
   U31086 : OAI222_X1 port map( A1 => n30750, A2 => n39593, B1 => n30814, B2 =>
                           n39587, C1 => n30686, C2 => n39581, ZN => n34433);
   U31087 : AOI221_X1 port map( B1 => n39353, B2 => n32992, C1 => n39347, C2 =>
                           n32944, A => n35707, ZN => n35702);
   U31088 : OAI222_X1 port map( A1 => n30750, A2 => n39341, B1 => n30814, B2 =>
                           n39335, C1 => n30686, C2 => n39329, ZN => n35707);
   U31089 : AOI221_X1 port map( B1 => n39605, B2 => n32991, C1 => n39599, C2 =>
                           n32943, A => n34452, ZN => n34447);
   U31090 : OAI222_X1 port map( A1 => n30749, A2 => n39593, B1 => n30813, B2 =>
                           n39587, C1 => n30685, C2 => n39581, ZN => n34452);
   U31091 : AOI221_X1 port map( B1 => n39353, B2 => n32991, C1 => n39347, C2 =>
                           n32943, A => n35726, ZN => n35721);
   U31092 : OAI222_X1 port map( A1 => n30749, A2 => n39341, B1 => n30813, B2 =>
                           n39335, C1 => n30685, C2 => n39329, ZN => n35726);
   U31093 : AOI221_X1 port map( B1 => n39604, B2 => n33134, C1 => n39598, C2 =>
                           n33122, A => n34471, ZN => n34466);
   U31094 : OAI222_X1 port map( A1 => n30748, A2 => n39592, B1 => n30812, B2 =>
                           n39586, C1 => n30684, C2 => n39580, ZN => n34471);
   U31095 : AOI221_X1 port map( B1 => n39352, B2 => n33134, C1 => n39346, C2 =>
                           n33122, A => n35745, ZN => n35740);
   U31096 : OAI222_X1 port map( A1 => n30748, A2 => n39340, B1 => n30812, B2 =>
                           n39334, C1 => n30684, C2 => n39328, ZN => n35745);
   U31097 : AOI221_X1 port map( B1 => n39604, B2 => n33133, C1 => n39598, C2 =>
                           n33121, A => n34490, ZN => n34485);
   U31098 : OAI222_X1 port map( A1 => n30747, A2 => n39592, B1 => n30811, B2 =>
                           n39586, C1 => n30683, C2 => n39580, ZN => n34490);
   U31099 : AOI221_X1 port map( B1 => n39352, B2 => n33133, C1 => n39346, C2 =>
                           n33121, A => n35764, ZN => n35759);
   U31100 : OAI222_X1 port map( A1 => n30747, A2 => n39340, B1 => n30811, B2 =>
                           n39334, C1 => n30683, C2 => n39328, ZN => n35764);
   U31101 : AOI221_X1 port map( B1 => n39604, B2 => n33132, C1 => n39598, C2 =>
                           n33120, A => n34509, ZN => n34504);
   U31102 : OAI222_X1 port map( A1 => n30746, A2 => n39592, B1 => n30810, B2 =>
                           n39586, C1 => n30682, C2 => n39580, ZN => n34509);
   U31103 : AOI221_X1 port map( B1 => n39352, B2 => n33132, C1 => n39346, C2 =>
                           n33120, A => n35783, ZN => n35778);
   U31104 : OAI222_X1 port map( A1 => n30746, A2 => n39340, B1 => n30810, B2 =>
                           n39334, C1 => n30682, C2 => n39328, ZN => n35783);
   U31105 : AOI221_X1 port map( B1 => n39604, B2 => n33131, C1 => n39598, C2 =>
                           n33119, A => n34528, ZN => n34523);
   U31106 : OAI222_X1 port map( A1 => n30745, A2 => n39592, B1 => n30809, B2 =>
                           n39586, C1 => n30681, C2 => n39580, ZN => n34528);
   U31107 : AOI221_X1 port map( B1 => n39352, B2 => n33131, C1 => n39346, C2 =>
                           n33119, A => n35802, ZN => n35797);
   U31108 : OAI222_X1 port map( A1 => n30745, A2 => n39340, B1 => n30809, B2 =>
                           n39334, C1 => n30681, C2 => n39328, ZN => n35802);
   U31109 : AOI221_X1 port map( B1 => n39604, B2 => n33130, C1 => n39598, C2 =>
                           n33118, A => n34547, ZN => n34542);
   U31110 : OAI222_X1 port map( A1 => n30744, A2 => n39592, B1 => n30808, B2 =>
                           n39586, C1 => n30680, C2 => n39580, ZN => n34547);
   U31111 : AOI221_X1 port map( B1 => n39352, B2 => n33130, C1 => n39346, C2 =>
                           n33118, A => n35821, ZN => n35816);
   U31112 : OAI222_X1 port map( A1 => n30744, A2 => n39340, B1 => n30808, B2 =>
                           n39334, C1 => n30680, C2 => n39328, ZN => n35821);
   U31113 : AOI221_X1 port map( B1 => n39604, B2 => n33129, C1 => n39598, C2 =>
                           n33117, A => n34566, ZN => n34561);
   U31114 : OAI222_X1 port map( A1 => n30743, A2 => n39592, B1 => n30807, B2 =>
                           n39586, C1 => n30679, C2 => n39580, ZN => n34566);
   U31115 : AOI221_X1 port map( B1 => n39352, B2 => n33129, C1 => n39346, C2 =>
                           n33117, A => n35840, ZN => n35835);
   U31116 : OAI222_X1 port map( A1 => n30743, A2 => n39340, B1 => n30807, B2 =>
                           n39334, C1 => n30679, C2 => n39328, ZN => n35840);
   U31117 : AOI221_X1 port map( B1 => n39604, B2 => n33128, C1 => n39598, C2 =>
                           n33116, A => n34585, ZN => n34580);
   U31118 : OAI222_X1 port map( A1 => n30742, A2 => n39592, B1 => n30806, B2 =>
                           n39586, C1 => n30678, C2 => n39580, ZN => n34585);
   U31119 : AOI221_X1 port map( B1 => n39352, B2 => n33128, C1 => n39346, C2 =>
                           n33116, A => n35859, ZN => n35854);
   U31120 : OAI222_X1 port map( A1 => n30742, A2 => n39340, B1 => n30806, B2 =>
                           n39334, C1 => n30678, C2 => n39328, ZN => n35859);
   U31121 : AOI221_X1 port map( B1 => n39604, B2 => n33127, C1 => n39598, C2 =>
                           n33115, A => n34604, ZN => n34599);
   U31122 : OAI222_X1 port map( A1 => n30741, A2 => n39592, B1 => n30805, B2 =>
                           n39586, C1 => n30677, C2 => n39580, ZN => n34604);
   U31123 : AOI221_X1 port map( B1 => n39352, B2 => n33127, C1 => n39346, C2 =>
                           n33115, A => n35878, ZN => n35873);
   U31124 : OAI222_X1 port map( A1 => n30741, A2 => n39340, B1 => n30805, B2 =>
                           n39334, C1 => n30677, C2 => n39328, ZN => n35878);
   U31125 : AOI221_X1 port map( B1 => n39604, B2 => n33126, C1 => n39598, C2 =>
                           n33114, A => n34623, ZN => n34618);
   U31126 : OAI222_X1 port map( A1 => n30740, A2 => n39592, B1 => n30804, B2 =>
                           n39586, C1 => n30676, C2 => n39580, ZN => n34623);
   U31127 : AOI221_X1 port map( B1 => n39352, B2 => n33126, C1 => n39346, C2 =>
                           n33114, A => n35897, ZN => n35892);
   U31128 : OAI222_X1 port map( A1 => n30740, A2 => n39340, B1 => n30804, B2 =>
                           n39334, C1 => n30676, C2 => n39328, ZN => n35897);
   U31129 : AOI221_X1 port map( B1 => n39604, B2 => n33125, C1 => n39598, C2 =>
                           n33113, A => n34642, ZN => n34637);
   U31130 : OAI222_X1 port map( A1 => n30739, A2 => n39592, B1 => n30803, B2 =>
                           n39586, C1 => n30675, C2 => n39580, ZN => n34642);
   U31131 : AOI221_X1 port map( B1 => n39352, B2 => n33125, C1 => n39346, C2 =>
                           n33113, A => n35916, ZN => n35911);
   U31132 : OAI222_X1 port map( A1 => n30739, A2 => n39340, B1 => n30803, B2 =>
                           n39334, C1 => n30675, C2 => n39328, ZN => n35916);
   U31133 : AOI221_X1 port map( B1 => n39604, B2 => n33124, C1 => n39598, C2 =>
                           n33112, A => n34661, ZN => n34656);
   U31134 : OAI222_X1 port map( A1 => n30738, A2 => n39592, B1 => n30802, B2 =>
                           n39586, C1 => n30674, C2 => n39580, ZN => n34661);
   U31135 : AOI221_X1 port map( B1 => n39352, B2 => n33124, C1 => n39346, C2 =>
                           n33112, A => n35935, ZN => n35930);
   U31136 : OAI222_X1 port map( A1 => n30738, A2 => n39340, B1 => n30802, B2 =>
                           n39334, C1 => n30674, C2 => n39328, ZN => n35935);
   U31137 : AOI221_X1 port map( B1 => n39604, B2 => n33123, C1 => n39598, C2 =>
                           n33111, A => n34692, ZN => n34686);
   U31138 : OAI222_X1 port map( A1 => n30737, A2 => n39592, B1 => n30801, B2 =>
                           n39586, C1 => n30673, C2 => n39580, ZN => n34692);
   U31139 : AOI221_X1 port map( B1 => n39352, B2 => n33123, C1 => n39346, C2 =>
                           n33111, A => n35966, ZN => n35960);
   U31140 : OAI222_X1 port map( A1 => n30737, A2 => n39340, B1 => n30801, B2 =>
                           n39334, C1 => n30673, C2 => n39328, ZN => n35966);
   U31141 : NAND2_X1 port map( A1 => n33330, A2 => n33294, ZN => n33394);
   U31142 : AND2_X1 port map( A1 => N6273, A2 => n32164, ZN => n34684);
   U31143 : AND2_X1 port map( A1 => N6398, A2 => n32169, ZN => n35958);
   U31144 : INV_X1 port map( A => n33398, ZN => n32254);
   U31145 : AND2_X1 port map( A1 => N6272, A2 => N6273, ZN => n34681);
   U31146 : AND2_X1 port map( A1 => N6397, A2 => N6398, ZN => n35955);
   U31147 : INV_X1 port map( A => n34694, ZN => n32168);
   U31148 : INV_X1 port map( A => n35968, ZN => n32173);
   U31149 : AND3_X1 port map( A1 => N931, A2 => n32151, A3 => n33331, ZN => 
                           n33367);
   U31150 : AND3_X1 port map( A1 => N932, A2 => N931, A3 => n33331, ZN => 
                           n33306);
   U31151 : AND3_X1 port map( A1 => N932, A2 => n32152, A3 => n33331, ZN => 
                           n33338);
   U31152 : AND3_X1 port map( A1 => n33294, A2 => n32150, A3 => n33300, ZN => 
                           n33257);
   U31153 : INV_X1 port map( A => n33402, ZN => n32163);
   U31154 : INV_X1 port map( A => N689, ZN => n32248);
   U31155 : INV_X1 port map( A => N6271, ZN => n32165);
   U31156 : INV_X1 port map( A => N6396, ZN => n32170);
   U31157 : INV_X1 port map( A => N688, ZN => n32251);
   U31158 : INV_X1 port map( A => N6270, ZN => n32166);
   U31159 : INV_X1 port map( A => N6395, ZN => n32171);
   U31160 : BUF_X1 port map( A => n33272, Z => n40522);
   U31161 : OAI211_X1 port map( C1 => n33256, C2 => n33274, A => n40521, B => 
                           n41368, ZN => n33272);
   U31162 : BUF_X1 port map( A => n33277, Z => n40502);
   U31163 : OAI211_X1 port map( C1 => n33256, C2 => n32157, A => n40501, B => 
                           n41367, ZN => n33277);
   U31164 : BUF_X1 port map( A => n33262, Z => n40562);
   U31165 : OAI211_X1 port map( C1 => n33256, C2 => n33264, A => n40561, B => 
                           n41367, ZN => n33262);
   U31166 : BUF_X1 port map( A => n33267, Z => n40542);
   U31167 : OAI211_X1 port map( C1 => n33256, C2 => n33269, A => n40541, B => 
                           n41368, ZN => n33267);
   U31168 : BUF_X1 port map( A => n33282, Z => n40482);
   U31169 : OAI211_X1 port map( C1 => n33256, C2 => n32158, A => n40481, B => 
                           n41367, ZN => n33282);
   U31170 : BUF_X1 port map( A => n33287, Z => n40462);
   U31171 : OAI211_X1 port map( C1 => n33256, C2 => n32159, A => n40461, B => 
                           n41367, ZN => n33287);
   U31172 : BUF_X1 port map( A => n33292, Z => n40442);
   U31173 : OAI211_X1 port map( C1 => n33256, C2 => n32160, A => n40441, B => 
                           n41367, ZN => n33292);
   U31174 : BUF_X1 port map( A => n33253, Z => n40582);
   U31175 : OAI211_X1 port map( C1 => n33255, C2 => n33256, A => n40581, B => 
                           n41367, ZN => n33253);
   U31176 : INV_X1 port map( A => N929, ZN => n32161);
   U31177 : INV_X1 port map( A => n37240, ZN => n32243);
   U31178 : AND2_X1 port map( A1 => n33301, A2 => n33299, ZN => n33333);
   U31179 : INV_X1 port map( A => N931, ZN => n32152);
   U31180 : INV_X1 port map( A => N932, ZN => n32151);
   U31181 : INV_X1 port map( A => N812, ZN => n32249);
   U31182 : AND2_X1 port map( A1 => n33301, A2 => n33300, ZN => n33331);
   U31183 : INV_X1 port map( A => n33362, ZN => n32239);
   U31184 : INV_X1 port map( A => N690, ZN => n32246);
   U31185 : INV_X1 port map( A => N6272, ZN => n32164);
   U31186 : INV_X1 port map( A => N6397, ZN => n32169);
   U31187 : INV_X1 port map( A => N813, ZN => n32247);
   U31188 : NAND2_X1 port map( A1 => add_136_carry_4_port, A2 => n32242, ZN => 
                           n37251);
   U31189 : NOR3_X1 port map( A1 => n33223, A2 => n32075, A3 => n33222, ZN => 
                           n33224);
   U31190 : INV_X1 port map( A => n39297, ZN => n39295);
   U31191 : INV_X1 port map( A => n39297, ZN => n39294);
   U31192 : INV_X1 port map( A => n39297, ZN => n39296);
   U31193 : OAI21_X1 port map( B1 => n33230, B2 => n33231, A => n33232, ZN => 
                           n33225);
   U31194 : AND3_X1 port map( A1 => n33233, A2 => n41370, A3 => n33237, ZN => 
                           n33249);
   U31195 : AND3_X1 port map( A1 => n33211, A2 => n33212, A3 => n33213, ZN => 
                           n33210);
   U31196 : NAND4_X1 port map( A1 => n33218, A2 => n33212, A3 => n41367, A4 => 
                           n32083, ZN => n33211);
   U31197 : OAI21_X1 port map( B1 => n33216, B2 => N659, A => n33245, ZN => 
                           n33244);
   U31198 : NAND4_X1 port map( A1 => n32241, A2 => n33239, A3 => n33245, A4 => 
                           n33218, ZN => n35977);
   U31199 : INV_X1 port map( A => n33238, ZN => n32241);
   U31200 : NAND4_X1 port map( A1 => n32323, A2 => n32322, A3 => n32260, A4 => 
                           n32258, ZN => n35976);
   U31201 : INV_X1 port map( A => n33233, ZN => n32077);
   U31202 : OAI21_X1 port map( B1 => n32322, B2 => n33225, A => n33226, ZN => 
                           n9896);
   U31203 : OAI21_X1 port map( B1 => n33222, B2 => n33223, A => n32322, ZN => 
                           n33226);
   U31204 : NOR2_X1 port map( A1 => n33224, A2 => n32260, ZN => n9899);
   U31205 : NOR2_X1 port map( A1 => n33224, A2 => n32258, ZN => n9897);
   U31206 : INV_X1 port map( A => n33234, ZN => n32076);
   U31207 : BUF_X1 port map( A => n32079, Z => n41368);
   U31208 : BUF_X1 port map( A => n32079, Z => n41369);
   U31209 : BUF_X1 port map( A => n32079, Z => n41370);
   U31210 : BUF_X1 port map( A => n32079, Z => n41367);
   U31211 : BUF_X1 port map( A => n32079, Z => n41364);
   U31212 : BUF_X1 port map( A => n32079, Z => n41366);
   U31213 : BUF_X1 port map( A => n32079, Z => n41365);
   U31214 : BUF_X1 port map( A => n33424, Z => n39796);
   U31215 : BUF_X1 port map( A => n34698, Z => n39544);
   U31216 : BUF_X1 port map( A => n33424, Z => n39800);
   U31217 : BUF_X1 port map( A => n34698, Z => n39548);
   U31218 : BUF_X1 port map( A => n33424, Z => n39799);
   U31219 : BUF_X1 port map( A => n34698, Z => n39547);
   U31220 : BUF_X1 port map( A => n33424, Z => n39798);
   U31221 : BUF_X1 port map( A => n34698, Z => n39546);
   U31222 : BUF_X1 port map( A => n33424, Z => n39797);
   U31223 : BUF_X1 port map( A => n34698, Z => n39545);
   U31224 : INV_X1 port map( A => n33208, ZN => n32167);
   U31225 : INV_X1 port map( A => n33207, ZN => n32172);
   U31226 : INV_X1 port map( A => n33209, ZN => n32162);
   U31227 : BUF_X1 port map( A => n32124, Z => n41118);
   U31228 : BUF_X1 port map( A => n32214, Z => n40734);
   U31229 : BUF_X1 port map( A => n32123, Z => n41124);
   U31230 : BUF_X1 port map( A => n32213, Z => n40740);
   U31231 : BUF_X1 port map( A => n32122, Z => n41130);
   U31232 : BUF_X1 port map( A => n32212, Z => n40746);
   U31233 : BUF_X1 port map( A => n32121, Z => n41136);
   U31234 : BUF_X1 port map( A => n32211, Z => n40752);
   U31235 : BUF_X1 port map( A => n32120, Z => n41142);
   U31236 : BUF_X1 port map( A => n32210, Z => n40758);
   U31237 : BUF_X1 port map( A => n32119, Z => n41148);
   U31238 : BUF_X1 port map( A => n32209, Z => n40764);
   U31239 : BUF_X1 port map( A => n32118, Z => n41154);
   U31240 : BUF_X1 port map( A => n32208, Z => n40770);
   U31241 : BUF_X1 port map( A => n32117, Z => n41160);
   U31242 : BUF_X1 port map( A => n32207, Z => n40776);
   U31243 : BUF_X1 port map( A => n32116, Z => n41166);
   U31244 : BUF_X1 port map( A => n32206, Z => n40782);
   U31245 : BUF_X1 port map( A => n32115, Z => n41172);
   U31246 : BUF_X1 port map( A => n32205, Z => n40788);
   U31247 : BUF_X1 port map( A => n32114, Z => n41178);
   U31248 : BUF_X1 port map( A => n32204, Z => n40794);
   U31249 : BUF_X1 port map( A => n32113, Z => n41184);
   U31250 : BUF_X1 port map( A => n32203, Z => n40800);
   U31251 : BUF_X1 port map( A => n32112, Z => n41190);
   U31252 : BUF_X1 port map( A => n32202, Z => n40806);
   U31253 : BUF_X1 port map( A => n32111, Z => n41196);
   U31254 : BUF_X1 port map( A => n32201, Z => n40812);
   U31255 : BUF_X1 port map( A => n32110, Z => n41202);
   U31256 : BUF_X1 port map( A => n32200, Z => n40818);
   U31257 : BUF_X1 port map( A => n32109, Z => n41208);
   U31258 : BUF_X1 port map( A => n32199, Z => n40824);
   U31259 : BUF_X1 port map( A => n32108, Z => n41214);
   U31260 : BUF_X1 port map( A => n32198, Z => n40830);
   U31261 : BUF_X1 port map( A => n32107, Z => n41220);
   U31262 : BUF_X1 port map( A => n32197, Z => n40836);
   U31263 : BUF_X1 port map( A => n32106, Z => n41226);
   U31264 : BUF_X1 port map( A => n32196, Z => n40842);
   U31265 : BUF_X1 port map( A => n32105, Z => n41232);
   U31266 : BUF_X1 port map( A => n32195, Z => n40848);
   U31267 : BUF_X1 port map( A => n32104, Z => n41238);
   U31268 : BUF_X1 port map( A => n32194, Z => n40854);
   U31269 : BUF_X1 port map( A => n32103, Z => n41244);
   U31270 : BUF_X1 port map( A => n32193, Z => n40860);
   U31271 : BUF_X1 port map( A => n32102, Z => n41250);
   U31272 : BUF_X1 port map( A => n32192, Z => n40866);
   U31273 : BUF_X1 port map( A => n32101, Z => n41256);
   U31274 : BUF_X1 port map( A => n32191, Z => n40872);
   U31275 : BUF_X1 port map( A => n32100, Z => n41262);
   U31276 : BUF_X1 port map( A => n32190, Z => n40878);
   U31277 : BUF_X1 port map( A => n32099, Z => n41268);
   U31278 : BUF_X1 port map( A => n32189, Z => n40884);
   U31279 : BUF_X1 port map( A => n32098, Z => n41274);
   U31280 : BUF_X1 port map( A => n32188, Z => n40890);
   U31281 : BUF_X1 port map( A => n32097, Z => n41280);
   U31282 : BUF_X1 port map( A => n32187, Z => n40896);
   U31283 : BUF_X1 port map( A => n32096, Z => n41286);
   U31284 : BUF_X1 port map( A => n32186, Z => n40902);
   U31285 : BUF_X1 port map( A => n32095, Z => n41292);
   U31286 : BUF_X1 port map( A => n32185, Z => n40908);
   U31287 : BUF_X1 port map( A => n32094, Z => n41298);
   U31288 : BUF_X1 port map( A => n32184, Z => n40914);
   U31289 : BUF_X1 port map( A => n32093, Z => n41304);
   U31290 : BUF_X1 port map( A => n32183, Z => n40920);
   U31291 : BUF_X1 port map( A => n32092, Z => n41310);
   U31292 : BUF_X1 port map( A => n32182, Z => n40926);
   U31293 : BUF_X1 port map( A => n32091, Z => n41316);
   U31294 : BUF_X1 port map( A => n32181, Z => n40932);
   U31295 : BUF_X1 port map( A => n32090, Z => n41322);
   U31296 : BUF_X1 port map( A => n32180, Z => n40938);
   U31297 : BUF_X1 port map( A => n32089, Z => n41328);
   U31298 : BUF_X1 port map( A => n32179, Z => n40944);
   U31299 : BUF_X1 port map( A => n32088, Z => n41334);
   U31300 : BUF_X1 port map( A => n32178, Z => n40950);
   U31301 : BUF_X1 port map( A => n32087, Z => n41340);
   U31302 : BUF_X1 port map( A => n32177, Z => n40956);
   U31303 : BUF_X1 port map( A => n32086, Z => n41346);
   U31304 : BUF_X1 port map( A => n32176, Z => n40962);
   U31305 : BUF_X1 port map( A => n32085, Z => n41352);
   U31306 : BUF_X1 port map( A => n32175, Z => n40968);
   U31307 : BUF_X1 port map( A => n32084, Z => n41358);
   U31308 : BUF_X1 port map( A => n32174, Z => n40974);
   U31309 : BUF_X1 port map( A => n32147, Z => n40980);
   U31310 : BUF_X1 port map( A => n32237, Z => n40596);
   U31311 : BUF_X1 port map( A => n32146, Z => n40986);
   U31312 : BUF_X1 port map( A => n32236, Z => n40602);
   U31313 : BUF_X1 port map( A => n32145, Z => n40992);
   U31314 : BUF_X1 port map( A => n32235, Z => n40608);
   U31315 : BUF_X1 port map( A => n32144, Z => n40998);
   U31316 : BUF_X1 port map( A => n32234, Z => n40614);
   U31317 : BUF_X1 port map( A => n32143, Z => n41004);
   U31318 : BUF_X1 port map( A => n32233, Z => n40620);
   U31319 : BUF_X1 port map( A => n32142, Z => n41010);
   U31320 : BUF_X1 port map( A => n32232, Z => n40626);
   U31321 : BUF_X1 port map( A => n32141, Z => n41016);
   U31322 : BUF_X1 port map( A => n32231, Z => n40632);
   U31323 : BUF_X1 port map( A => n32140, Z => n41022);
   U31324 : BUF_X1 port map( A => n32230, Z => n40638);
   U31325 : BUF_X1 port map( A => n32139, Z => n41028);
   U31326 : BUF_X1 port map( A => n32229, Z => n40644);
   U31327 : BUF_X1 port map( A => n32138, Z => n41034);
   U31328 : BUF_X1 port map( A => n32228, Z => n40650);
   U31329 : BUF_X1 port map( A => n32137, Z => n41040);
   U31330 : BUF_X1 port map( A => n32227, Z => n40656);
   U31331 : BUF_X1 port map( A => n32136, Z => n41046);
   U31332 : BUF_X1 port map( A => n32226, Z => n40662);
   U31333 : BUF_X1 port map( A => n32135, Z => n41052);
   U31334 : BUF_X1 port map( A => n32225, Z => n40668);
   U31335 : BUF_X1 port map( A => n32134, Z => n41058);
   U31336 : BUF_X1 port map( A => n32224, Z => n40674);
   U31337 : BUF_X1 port map( A => n32133, Z => n41064);
   U31338 : BUF_X1 port map( A => n32223, Z => n40680);
   U31339 : BUF_X1 port map( A => n32132, Z => n41070);
   U31340 : BUF_X1 port map( A => n32222, Z => n40686);
   U31341 : BUF_X1 port map( A => n32131, Z => n41076);
   U31342 : BUF_X1 port map( A => n32221, Z => n40692);
   U31343 : BUF_X1 port map( A => n32130, Z => n41082);
   U31344 : BUF_X1 port map( A => n32220, Z => n40698);
   U31345 : BUF_X1 port map( A => n32129, Z => n41088);
   U31346 : BUF_X1 port map( A => n32219, Z => n40704);
   U31347 : BUF_X1 port map( A => n32128, Z => n41094);
   U31348 : BUF_X1 port map( A => n32218, Z => n40710);
   U31349 : BUF_X1 port map( A => n32127, Z => n41100);
   U31350 : BUF_X1 port map( A => n32217, Z => n40716);
   U31351 : BUF_X1 port map( A => n32126, Z => n41106);
   U31352 : BUF_X1 port map( A => n32216, Z => n40722);
   U31353 : BUF_X1 port map( A => n32125, Z => n41112);
   U31354 : BUF_X1 port map( A => n32215, Z => n40728);
   U31355 : BUF_X1 port map( A => n32147, Z => n40981);
   U31356 : BUF_X1 port map( A => n32237, Z => n40597);
   U31357 : BUF_X1 port map( A => n32146, Z => n40987);
   U31358 : BUF_X1 port map( A => n32236, Z => n40603);
   U31359 : BUF_X1 port map( A => n32145, Z => n40993);
   U31360 : BUF_X1 port map( A => n32235, Z => n40609);
   U31361 : BUF_X1 port map( A => n32144, Z => n40999);
   U31362 : BUF_X1 port map( A => n32234, Z => n40615);
   U31363 : BUF_X1 port map( A => n32143, Z => n41005);
   U31364 : BUF_X1 port map( A => n32233, Z => n40621);
   U31365 : BUF_X1 port map( A => n32142, Z => n41011);
   U31366 : BUF_X1 port map( A => n32232, Z => n40627);
   U31367 : BUF_X1 port map( A => n32141, Z => n41017);
   U31368 : BUF_X1 port map( A => n32231, Z => n40633);
   U31369 : BUF_X1 port map( A => n32140, Z => n41023);
   U31370 : BUF_X1 port map( A => n32230, Z => n40639);
   U31371 : BUF_X1 port map( A => n32139, Z => n41029);
   U31372 : BUF_X1 port map( A => n32229, Z => n40645);
   U31373 : BUF_X1 port map( A => n32138, Z => n41035);
   U31374 : BUF_X1 port map( A => n32228, Z => n40651);
   U31375 : BUF_X1 port map( A => n32137, Z => n41041);
   U31376 : BUF_X1 port map( A => n32227, Z => n40657);
   U31377 : BUF_X1 port map( A => n32136, Z => n41047);
   U31378 : BUF_X1 port map( A => n32226, Z => n40663);
   U31379 : BUF_X1 port map( A => n32135, Z => n41053);
   U31380 : BUF_X1 port map( A => n32225, Z => n40669);
   U31381 : BUF_X1 port map( A => n32134, Z => n41059);
   U31382 : BUF_X1 port map( A => n32224, Z => n40675);
   U31383 : BUF_X1 port map( A => n32133, Z => n41065);
   U31384 : BUF_X1 port map( A => n32223, Z => n40681);
   U31385 : BUF_X1 port map( A => n32132, Z => n41071);
   U31386 : BUF_X1 port map( A => n32222, Z => n40687);
   U31387 : BUF_X1 port map( A => n32131, Z => n41077);
   U31388 : BUF_X1 port map( A => n32221, Z => n40693);
   U31389 : BUF_X1 port map( A => n32130, Z => n41083);
   U31390 : BUF_X1 port map( A => n32220, Z => n40699);
   U31391 : BUF_X1 port map( A => n32129, Z => n41089);
   U31392 : BUF_X1 port map( A => n32219, Z => n40705);
   U31393 : BUF_X1 port map( A => n32128, Z => n41095);
   U31394 : BUF_X1 port map( A => n32218, Z => n40711);
   U31395 : BUF_X1 port map( A => n32127, Z => n41101);
   U31396 : BUF_X1 port map( A => n32217, Z => n40717);
   U31397 : BUF_X1 port map( A => n32126, Z => n41107);
   U31398 : BUF_X1 port map( A => n32216, Z => n40723);
   U31399 : BUF_X1 port map( A => n32125, Z => n41113);
   U31400 : BUF_X1 port map( A => n32215, Z => n40729);
   U31401 : BUF_X1 port map( A => n32124, Z => n41119);
   U31402 : BUF_X1 port map( A => n32214, Z => n40735);
   U31403 : BUF_X1 port map( A => n32123, Z => n41125);
   U31404 : BUF_X1 port map( A => n32213, Z => n40741);
   U31405 : BUF_X1 port map( A => n32122, Z => n41131);
   U31406 : BUF_X1 port map( A => n32212, Z => n40747);
   U31407 : BUF_X1 port map( A => n32121, Z => n41137);
   U31408 : BUF_X1 port map( A => n32211, Z => n40753);
   U31409 : BUF_X1 port map( A => n32120, Z => n41143);
   U31410 : BUF_X1 port map( A => n32210, Z => n40759);
   U31411 : BUF_X1 port map( A => n32119, Z => n41149);
   U31412 : BUF_X1 port map( A => n32209, Z => n40765);
   U31413 : BUF_X1 port map( A => n32118, Z => n41155);
   U31414 : BUF_X1 port map( A => n32208, Z => n40771);
   U31415 : BUF_X1 port map( A => n32117, Z => n41161);
   U31416 : BUF_X1 port map( A => n32207, Z => n40777);
   U31417 : BUF_X1 port map( A => n32116, Z => n41167);
   U31418 : BUF_X1 port map( A => n32206, Z => n40783);
   U31419 : BUF_X1 port map( A => n32115, Z => n41173);
   U31420 : BUF_X1 port map( A => n32205, Z => n40789);
   U31421 : BUF_X1 port map( A => n32114, Z => n41179);
   U31422 : BUF_X1 port map( A => n32204, Z => n40795);
   U31423 : BUF_X1 port map( A => n32113, Z => n41185);
   U31424 : BUF_X1 port map( A => n32203, Z => n40801);
   U31425 : BUF_X1 port map( A => n32112, Z => n41191);
   U31426 : BUF_X1 port map( A => n32202, Z => n40807);
   U31427 : BUF_X1 port map( A => n32111, Z => n41197);
   U31428 : BUF_X1 port map( A => n32201, Z => n40813);
   U31429 : BUF_X1 port map( A => n32110, Z => n41203);
   U31430 : BUF_X1 port map( A => n32200, Z => n40819);
   U31431 : BUF_X1 port map( A => n32109, Z => n41209);
   U31432 : BUF_X1 port map( A => n32199, Z => n40825);
   U31433 : BUF_X1 port map( A => n32108, Z => n41215);
   U31434 : BUF_X1 port map( A => n32198, Z => n40831);
   U31435 : BUF_X1 port map( A => n32107, Z => n41221);
   U31436 : BUF_X1 port map( A => n32197, Z => n40837);
   U31437 : BUF_X1 port map( A => n32106, Z => n41227);
   U31438 : BUF_X1 port map( A => n32196, Z => n40843);
   U31439 : BUF_X1 port map( A => n32105, Z => n41233);
   U31440 : BUF_X1 port map( A => n32195, Z => n40849);
   U31441 : BUF_X1 port map( A => n32104, Z => n41239);
   U31442 : BUF_X1 port map( A => n32194, Z => n40855);
   U31443 : BUF_X1 port map( A => n32103, Z => n41245);
   U31444 : BUF_X1 port map( A => n32193, Z => n40861);
   U31445 : BUF_X1 port map( A => n32102, Z => n41251);
   U31446 : BUF_X1 port map( A => n32192, Z => n40867);
   U31447 : BUF_X1 port map( A => n32101, Z => n41257);
   U31448 : BUF_X1 port map( A => n32191, Z => n40873);
   U31449 : BUF_X1 port map( A => n32100, Z => n41263);
   U31450 : BUF_X1 port map( A => n32190, Z => n40879);
   U31451 : BUF_X1 port map( A => n32099, Z => n41269);
   U31452 : BUF_X1 port map( A => n32189, Z => n40885);
   U31453 : BUF_X1 port map( A => n32098, Z => n41275);
   U31454 : BUF_X1 port map( A => n32188, Z => n40891);
   U31455 : BUF_X1 port map( A => n32097, Z => n41281);
   U31456 : BUF_X1 port map( A => n32187, Z => n40897);
   U31457 : BUF_X1 port map( A => n32096, Z => n41287);
   U31458 : BUF_X1 port map( A => n32186, Z => n40903);
   U31459 : BUF_X1 port map( A => n32095, Z => n41293);
   U31460 : BUF_X1 port map( A => n32185, Z => n40909);
   U31461 : BUF_X1 port map( A => n32094, Z => n41299);
   U31462 : BUF_X1 port map( A => n32184, Z => n40915);
   U31463 : BUF_X1 port map( A => n32093, Z => n41305);
   U31464 : BUF_X1 port map( A => n32183, Z => n40921);
   U31465 : BUF_X1 port map( A => n32092, Z => n41311);
   U31466 : BUF_X1 port map( A => n32182, Z => n40927);
   U31467 : BUF_X1 port map( A => n32091, Z => n41317);
   U31468 : BUF_X1 port map( A => n32181, Z => n40933);
   U31469 : BUF_X1 port map( A => n32090, Z => n41323);
   U31470 : BUF_X1 port map( A => n32180, Z => n40939);
   U31471 : BUF_X1 port map( A => n32089, Z => n41329);
   U31472 : BUF_X1 port map( A => n32179, Z => n40945);
   U31473 : BUF_X1 port map( A => n32088, Z => n41335);
   U31474 : BUF_X1 port map( A => n32178, Z => n40951);
   U31475 : BUF_X1 port map( A => n32087, Z => n41341);
   U31476 : BUF_X1 port map( A => n32177, Z => n40957);
   U31477 : BUF_X1 port map( A => n32086, Z => n41347);
   U31478 : BUF_X1 port map( A => n32176, Z => n40963);
   U31479 : BUF_X1 port map( A => n32085, Z => n41353);
   U31480 : BUF_X1 port map( A => n32175, Z => n40969);
   U31481 : BUF_X1 port map( A => n32084, Z => n41359);
   U31482 : BUF_X1 port map( A => n32174, Z => n40975);
   U31483 : NAND2_X1 port map( A1 => n32253, A2 => n33208, ZN => n34696);
   U31484 : NAND2_X1 port map( A1 => n32253, A2 => n33207, ZN => n35970);
   U31485 : NAND2_X1 port map( A1 => n32253, A2 => n33209, ZN => n33423);
   U31486 : NOR3_X1 port map( A1 => n32239, A2 => n23853, A3 => N813, ZN => 
                           n33298);
   U31487 : NOR2_X1 port map( A1 => n2695, A2 => n32162, ZN => U3_U193_Z_4);
   U31488 : AOI221_X1 port map( B1 => n39287, B2 => n30006, C1 => n39281, C2 =>
                           n30070, A => n36085, ZN => n36084);
   U31489 : OAI222_X1 port map( A1 => n31994, A2 => n39275, B1 => n32286, B2 =>
                           n39269, C1 => n31934, C2 => n39263, ZN => n36085);
   U31490 : AOI221_X1 port map( B1 => n39287, B2 => n30005, C1 => n39281, C2 =>
                           n30069, A => n36066, ZN => n36065);
   U31491 : OAI222_X1 port map( A1 => n31993, A2 => n39275, B1 => n32053, B2 =>
                           n39269, C1 => n31933, C2 => n39263, ZN => n36066);
   U31492 : AOI221_X1 port map( B1 => n39287, B2 => n30004, C1 => n39281, C2 =>
                           n30068, A => n36047, ZN => n36046);
   U31493 : OAI222_X1 port map( A1 => n31992, A2 => n39275, B1 => n32052, B2 =>
                           n39269, C1 => n31932, C2 => n39263, ZN => n36047);
   U31494 : AOI221_X1 port map( B1 => n39287, B2 => n30003, C1 => n39281, C2 =>
                           n30067, A => n35990, ZN => n35987);
   U31495 : OAI222_X1 port map( A1 => n31991, A2 => n39275, B1 => n32051, B2 =>
                           n39269, C1 => n31931, C2 => n39263, ZN => n35990);
   U31496 : OAI222_X1 port map( A1 => n40954, A2 => n40430, B1 => n41338, B2 =>
                           n40423, C1 => n40421, C2 => n33199, ZN => n9319);
   U31497 : OAI222_X1 port map( A1 => n40966, A2 => n40430, B1 => n41350, B2 =>
                           n40423, C1 => n40421, C2 => n33197, ZN => n9317);
   U31498 : OAI222_X1 port map( A1 => n40972, A2 => n40430, B1 => n41356, B2 =>
                           n40423, C1 => n40421, C2 => n33196, ZN => n9316);
   U31499 : OAI222_X1 port map( A1 => n40978, A2 => n40430, B1 => n41362, B2 =>
                           n40423, C1 => n40421, C2 => n33195, ZN => n9315);
   U31500 : OAI222_X1 port map( A1 => n40954, A2 => n40410, B1 => n41338, B2 =>
                           n40403, C1 => n40401, C2 => n33139, ZN => n9255);
   U31501 : OAI222_X1 port map( A1 => n40966, A2 => n40410, B1 => n41350, B2 =>
                           n40403, C1 => n40401, C2 => n33137, ZN => n9253);
   U31502 : OAI222_X1 port map( A1 => n40972, A2 => n40410, B1 => n41356, B2 =>
                           n40403, C1 => n40401, C2 => n33136, ZN => n9252);
   U31503 : OAI222_X1 port map( A1 => n40978, A2 => n40410, B1 => n41362, B2 =>
                           n40403, C1 => n40401, C2 => n33135, ZN => n9251);
   U31504 : OAI222_X1 port map( A1 => n40953, A2 => n40210, B1 => n41337, B2 =>
                           n40203, C1 => n40201, C2 => n33103, ZN => n8615);
   U31505 : OAI222_X1 port map( A1 => n40965, A2 => n40210, B1 => n41349, B2 =>
                           n40203, C1 => n40201, C2 => n33101, ZN => n8613);
   U31506 : OAI222_X1 port map( A1 => n40971, A2 => n40210, B1 => n41355, B2 =>
                           n40203, C1 => n40201, C2 => n33100, ZN => n8612);
   U31507 : OAI222_X1 port map( A1 => n40977, A2 => n40210, B1 => n41361, B2 =>
                           n40203, C1 => n40201, C2 => n33099, ZN => n8611);
   U31508 : OAI222_X1 port map( A1 => n40953, A2 => n40230, B1 => n41337, B2 =>
                           n40223, C1 => n40221, C2 => n33091, ZN => n8679);
   U31509 : OAI222_X1 port map( A1 => n40965, A2 => n40230, B1 => n41349, B2 =>
                           n40223, C1 => n40221, C2 => n33089, ZN => n8677);
   U31510 : OAI222_X1 port map( A1 => n40971, A2 => n40230, B1 => n41355, B2 =>
                           n40223, C1 => n40221, C2 => n33088, ZN => n8676);
   U31511 : OAI222_X1 port map( A1 => n40977, A2 => n40230, B1 => n41361, B2 =>
                           n40223, C1 => n40221, C2 => n33087, ZN => n8675);
   U31512 : OAI222_X1 port map( A1 => n40954, A2 => n40310, B1 => n41338, B2 =>
                           n40303, C1 => n40301, C2 => n32719, ZN => n8935);
   U31513 : OAI222_X1 port map( A1 => n40966, A2 => n40310, B1 => n41350, B2 =>
                           n40303, C1 => n40301, C2 => n32717, ZN => n8933);
   U31514 : OAI222_X1 port map( A1 => n40972, A2 => n40310, B1 => n41356, B2 =>
                           n40303, C1 => n40301, C2 => n32716, ZN => n8932);
   U31515 : OAI222_X1 port map( A1 => n40978, A2 => n40310, B1 => n41362, B2 =>
                           n40303, C1 => n40301, C2 => n32715, ZN => n8931);
   U31516 : OAI222_X1 port map( A1 => n40954, A2 => n40330, B1 => n41338, B2 =>
                           n40323, C1 => n40321, C2 => n32707, ZN => n8999);
   U31517 : OAI222_X1 port map( A1 => n40966, A2 => n40330, B1 => n41350, B2 =>
                           n40323, C1 => n40321, C2 => n32705, ZN => n8997);
   U31518 : OAI222_X1 port map( A1 => n40972, A2 => n40330, B1 => n41356, B2 =>
                           n40323, C1 => n40321, C2 => n32704, ZN => n8996);
   U31519 : OAI222_X1 port map( A1 => n40978, A2 => n40330, B1 => n41362, B2 =>
                           n40323, C1 => n40321, C2 => n32703, ZN => n8995);
   U31520 : OAI222_X1 port map( A1 => n40955, A2 => n40530, B1 => n41339, B2 =>
                           n40523, C1 => n40521, C2 => n32444, ZN => n9639);
   U31521 : OAI222_X1 port map( A1 => n40967, A2 => n40530, B1 => n41351, B2 =>
                           n40523, C1 => n40521, C2 => n38791, ZN => n9637);
   U31522 : OAI222_X1 port map( A1 => n40973, A2 => n40530, B1 => n41357, B2 =>
                           n40523, C1 => n40521, C2 => n38792, ZN => n9636);
   U31523 : OAI222_X1 port map( A1 => n40979, A2 => n40530, B1 => n41363, B2 =>
                           n40523, C1 => n40521, C2 => n38793, ZN => n9635);
   U31524 : OAI222_X1 port map( A1 => n40954, A2 => n40510, B1 => n41338, B2 =>
                           n40503, C1 => n40501, C2 => n32384, ZN => n9575);
   U31525 : OAI222_X1 port map( A1 => n40966, A2 => n40510, B1 => n41350, B2 =>
                           n40503, C1 => n40501, C2 => n38924, ZN => n9573);
   U31526 : OAI222_X1 port map( A1 => n40972, A2 => n40510, B1 => n41356, B2 =>
                           n40503, C1 => n40501, C2 => n38925, ZN => n9572);
   U31527 : OAI222_X1 port map( A1 => n40978, A2 => n40510, B1 => n41362, B2 =>
                           n40503, C1 => n40501, C2 => n38926, ZN => n9571);
   U31528 : OAI222_X1 port map( A1 => n40952, A2 => n39835, B1 => n41336, B2 =>
                           n39828, C1 => n39826, C2 => n32695, ZN => n7399);
   U31529 : OAI222_X1 port map( A1 => n40964, A2 => n39835, B1 => n41348, B2 =>
                           n39828, C1 => n39826, C2 => n32693, ZN => n7397);
   U31530 : OAI222_X1 port map( A1 => n40970, A2 => n39835, B1 => n41354, B2 =>
                           n39828, C1 => n39826, C2 => n32692, ZN => n7396);
   U31531 : OAI222_X1 port map( A1 => n40976, A2 => n39835, B1 => n41360, B2 =>
                           n39828, C1 => n39826, C2 => n32691, ZN => n7395);
   U31532 : NOR3_X1 port map( A1 => n33297, A2 => n23853, A3 => n32081, ZN => 
                           n33332);
   U31533 : AOI221_X1 port map( B1 => n39282, B2 => n30055, C1 => n39276, C2 =>
                           n30119, A => n37016, ZN => n37015);
   U31534 : OAI222_X1 port map( A1 => n32043, A2 => n39270, B1 => n32067, B2 =>
                           n39264, C1 => n31983, C2 => n39258, ZN => n37016);
   U31535 : AOI221_X1 port map( B1 => n39283, B2 => n30054, C1 => n39277, C2 =>
                           n30118, A => n36997, ZN => n36996);
   U31536 : OAI222_X1 port map( A1 => n32042, A2 => n39271, B1 => n32066, B2 =>
                           n39265, C1 => n31982, C2 => n39259, ZN => n36997);
   U31537 : AOI221_X1 port map( B1 => n39283, B2 => n30053, C1 => n39277, C2 =>
                           n30117, A => n36978, ZN => n36977);
   U31538 : OAI222_X1 port map( A1 => n32041, A2 => n39271, B1 => n32065, B2 =>
                           n39265, C1 => n31981, C2 => n39259, ZN => n36978);
   U31539 : AOI221_X1 port map( B1 => n39283, B2 => n30052, C1 => n39277, C2 =>
                           n30116, A => n36959, ZN => n36958);
   U31540 : OAI222_X1 port map( A1 => n32040, A2 => n39271, B1 => n32064, B2 =>
                           n39265, C1 => n31980, C2 => n39259, ZN => n36959);
   U31541 : AOI221_X1 port map( B1 => n39283, B2 => n30051, C1 => n39277, C2 =>
                           n30115, A => n36940, ZN => n36939);
   U31542 : OAI222_X1 port map( A1 => n32039, A2 => n39271, B1 => n32063, B2 =>
                           n39265, C1 => n31979, C2 => n39259, ZN => n36940);
   U31543 : AOI221_X1 port map( B1 => n39283, B2 => n30050, C1 => n39277, C2 =>
                           n30114, A => n36921, ZN => n36920);
   U31544 : OAI222_X1 port map( A1 => n32038, A2 => n39271, B1 => n32062, B2 =>
                           n39265, C1 => n31978, C2 => n39259, ZN => n36921);
   U31545 : AOI221_X1 port map( B1 => n39283, B2 => n30049, C1 => n39277, C2 =>
                           n30113, A => n36902, ZN => n36901);
   U31546 : OAI222_X1 port map( A1 => n32037, A2 => n39271, B1 => n32061, B2 =>
                           n39265, C1 => n31977, C2 => n39259, ZN => n36902);
   U31547 : AOI221_X1 port map( B1 => n39283, B2 => n30048, C1 => n39277, C2 =>
                           n30112, A => n36883, ZN => n36882);
   U31548 : OAI222_X1 port map( A1 => n32036, A2 => n39271, B1 => n32060, B2 =>
                           n39265, C1 => n31976, C2 => n39259, ZN => n36883);
   U31549 : AOI221_X1 port map( B1 => n39283, B2 => n30047, C1 => n39277, C2 =>
                           n30111, A => n36864, ZN => n36863);
   U31550 : OAI222_X1 port map( A1 => n32035, A2 => n39271, B1 => n32059, B2 =>
                           n39265, C1 => n31975, C2 => n39259, ZN => n36864);
   U31551 : AOI221_X1 port map( B1 => n39283, B2 => n30046, C1 => n39277, C2 =>
                           n30110, A => n36845, ZN => n36844);
   U31552 : OAI222_X1 port map( A1 => n32034, A2 => n39271, B1 => n32058, B2 =>
                           n39265, C1 => n31974, C2 => n39259, ZN => n36845);
   U31553 : AOI221_X1 port map( B1 => n39283, B2 => n30045, C1 => n39277, C2 =>
                           n30109, A => n36826, ZN => n36825);
   U31554 : OAI222_X1 port map( A1 => n32033, A2 => n39271, B1 => n32057, B2 =>
                           n39265, C1 => n31973, C2 => n39259, ZN => n36826);
   U31555 : AOI221_X1 port map( B1 => n39283, B2 => n30044, C1 => n39277, C2 =>
                           n30108, A => n36807, ZN => n36806);
   U31556 : OAI222_X1 port map( A1 => n32032, A2 => n39271, B1 => n32056, B2 =>
                           n39265, C1 => n31972, C2 => n39259, ZN => n36807);
   U31557 : AOI221_X1 port map( B1 => n39283, B2 => n30043, C1 => n39277, C2 =>
                           n30107, A => n36788, ZN => n36787);
   U31558 : OAI222_X1 port map( A1 => n32031, A2 => n39271, B1 => n32055, B2 =>
                           n39265, C1 => n31971, C2 => n39259, ZN => n36788);
   U31559 : AOI221_X1 port map( B1 => n39284, B2 => n30042, C1 => n39278, C2 =>
                           n30106, A => n36769, ZN => n36768);
   U31560 : OAI222_X1 port map( A1 => n32030, A2 => n39272, B1 => n32321, B2 =>
                           n39266, C1 => n31970, C2 => n39260, ZN => n36769);
   U31561 : AOI221_X1 port map( B1 => n39284, B2 => n30041, C1 => n39278, C2 =>
                           n30105, A => n36750, ZN => n36749);
   U31562 : OAI222_X1 port map( A1 => n32029, A2 => n39272, B1 => n32320, B2 =>
                           n39266, C1 => n31969, C2 => n39260, ZN => n36750);
   U31563 : AOI221_X1 port map( B1 => n39284, B2 => n30040, C1 => n39278, C2 =>
                           n30104, A => n36731, ZN => n36730);
   U31564 : OAI222_X1 port map( A1 => n32028, A2 => n39272, B1 => n32319, B2 =>
                           n39266, C1 => n31968, C2 => n39260, ZN => n36731);
   U31565 : AOI221_X1 port map( B1 => n39284, B2 => n30039, C1 => n39278, C2 =>
                           n30103, A => n36712, ZN => n36711);
   U31566 : OAI222_X1 port map( A1 => n32027, A2 => n39272, B1 => n32318, B2 =>
                           n39266, C1 => n31967, C2 => n39260, ZN => n36712);
   U31567 : AOI221_X1 port map( B1 => n39284, B2 => n30038, C1 => n39278, C2 =>
                           n30102, A => n36693, ZN => n36692);
   U31568 : OAI222_X1 port map( A1 => n32026, A2 => n39272, B1 => n32317, B2 =>
                           n39266, C1 => n31966, C2 => n39260, ZN => n36693);
   U31569 : AOI221_X1 port map( B1 => n39284, B2 => n30037, C1 => n39278, C2 =>
                           n30101, A => n36674, ZN => n36673);
   U31570 : OAI222_X1 port map( A1 => n32025, A2 => n39272, B1 => n32316, B2 =>
                           n39266, C1 => n31965, C2 => n39260, ZN => n36674);
   U31571 : AOI221_X1 port map( B1 => n39284, B2 => n30036, C1 => n39278, C2 =>
                           n30100, A => n36655, ZN => n36654);
   U31572 : OAI222_X1 port map( A1 => n32024, A2 => n39272, B1 => n32315, B2 =>
                           n39266, C1 => n31964, C2 => n39260, ZN => n36655);
   U31573 : AOI221_X1 port map( B1 => n39284, B2 => n30035, C1 => n39278, C2 =>
                           n30099, A => n36636, ZN => n36635);
   U31574 : OAI222_X1 port map( A1 => n32023, A2 => n39272, B1 => n32314, B2 =>
                           n39266, C1 => n31963, C2 => n39260, ZN => n36636);
   U31575 : AOI221_X1 port map( B1 => n39284, B2 => n30034, C1 => n39278, C2 =>
                           n30098, A => n36617, ZN => n36616);
   U31576 : OAI222_X1 port map( A1 => n32022, A2 => n39272, B1 => n32313, B2 =>
                           n39266, C1 => n31962, C2 => n39260, ZN => n36617);
   U31577 : AOI221_X1 port map( B1 => n39284, B2 => n30033, C1 => n39278, C2 =>
                           n30097, A => n36598, ZN => n36597);
   U31578 : OAI222_X1 port map( A1 => n32021, A2 => n39272, B1 => n32312, B2 =>
                           n39266, C1 => n31961, C2 => n39260, ZN => n36598);
   U31579 : AOI221_X1 port map( B1 => n39284, B2 => n30032, C1 => n39278, C2 =>
                           n30096, A => n36579, ZN => n36578);
   U31580 : OAI222_X1 port map( A1 => n32020, A2 => n39272, B1 => n32311, B2 =>
                           n39266, C1 => n31960, C2 => n39260, ZN => n36579);
   U31581 : AOI221_X1 port map( B1 => n39284, B2 => n30031, C1 => n39278, C2 =>
                           n30095, A => n36560, ZN => n36559);
   U31582 : OAI222_X1 port map( A1 => n32019, A2 => n39272, B1 => n32310, B2 =>
                           n39266, C1 => n31959, C2 => n39260, ZN => n36560);
   U31583 : AOI221_X1 port map( B1 => n39285, B2 => n30030, C1 => n39279, C2 =>
                           n30094, A => n36541, ZN => n36540);
   U31584 : OAI222_X1 port map( A1 => n32018, A2 => n39273, B1 => n32309, B2 =>
                           n39267, C1 => n31958, C2 => n39261, ZN => n36541);
   U31585 : AOI221_X1 port map( B1 => n39285, B2 => n30029, C1 => n39279, C2 =>
                           n30093, A => n36522, ZN => n36521);
   U31586 : OAI222_X1 port map( A1 => n32017, A2 => n39273, B1 => n32308, B2 =>
                           n39267, C1 => n31957, C2 => n39261, ZN => n36522);
   U31587 : AOI221_X1 port map( B1 => n39285, B2 => n30028, C1 => n39279, C2 =>
                           n30092, A => n36503, ZN => n36502);
   U31588 : OAI222_X1 port map( A1 => n32016, A2 => n39273, B1 => n32307, B2 =>
                           n39267, C1 => n31956, C2 => n39261, ZN => n36503);
   U31589 : AOI221_X1 port map( B1 => n39285, B2 => n30027, C1 => n39279, C2 =>
                           n30091, A => n36484, ZN => n36483);
   U31590 : OAI222_X1 port map( A1 => n32015, A2 => n39273, B1 => n32306, B2 =>
                           n39267, C1 => n31955, C2 => n39261, ZN => n36484);
   U31591 : AOI221_X1 port map( B1 => n39285, B2 => n30026, C1 => n39279, C2 =>
                           n30090, A => n36465, ZN => n36464);
   U31592 : OAI222_X1 port map( A1 => n32014, A2 => n39273, B1 => n32305, B2 =>
                           n39267, C1 => n31954, C2 => n39261, ZN => n36465);
   U31593 : AOI221_X1 port map( B1 => n39285, B2 => n30025, C1 => n39279, C2 =>
                           n30089, A => n36446, ZN => n36445);
   U31594 : OAI222_X1 port map( A1 => n32013, A2 => n39273, B1 => n32304, B2 =>
                           n39267, C1 => n31953, C2 => n39261, ZN => n36446);
   U31595 : AOI221_X1 port map( B1 => n39285, B2 => n30024, C1 => n39279, C2 =>
                           n30088, A => n36427, ZN => n36426);
   U31596 : OAI222_X1 port map( A1 => n32012, A2 => n39273, B1 => n32303, B2 =>
                           n39267, C1 => n31952, C2 => n39261, ZN => n36427);
   U31597 : AOI221_X1 port map( B1 => n39285, B2 => n30023, C1 => n39279, C2 =>
                           n30087, A => n36408, ZN => n36407);
   U31598 : OAI222_X1 port map( A1 => n32011, A2 => n39273, B1 => n32302, B2 =>
                           n39267, C1 => n31951, C2 => n39261, ZN => n36408);
   U31599 : AOI221_X1 port map( B1 => n39285, B2 => n30022, C1 => n39279, C2 =>
                           n30086, A => n36389, ZN => n36388);
   U31600 : OAI222_X1 port map( A1 => n32010, A2 => n39273, B1 => n32301, B2 =>
                           n39267, C1 => n31950, C2 => n39261, ZN => n36389);
   U31601 : AOI221_X1 port map( B1 => n39285, B2 => n30021, C1 => n39279, C2 =>
                           n30085, A => n36370, ZN => n36369);
   U31602 : OAI222_X1 port map( A1 => n32009, A2 => n39273, B1 => n32300, B2 =>
                           n39267, C1 => n31949, C2 => n39261, ZN => n36370);
   U31603 : AOI221_X1 port map( B1 => n39285, B2 => n30020, C1 => n39279, C2 =>
                           n30084, A => n36351, ZN => n36350);
   U31604 : OAI222_X1 port map( A1 => n32008, A2 => n39273, B1 => n32299, B2 =>
                           n39267, C1 => n31948, C2 => n39261, ZN => n36351);
   U31605 : AOI221_X1 port map( B1 => n39285, B2 => n30019, C1 => n39279, C2 =>
                           n30083, A => n36332, ZN => n36331);
   U31606 : OAI222_X1 port map( A1 => n32007, A2 => n39273, B1 => n32298, B2 =>
                           n39267, C1 => n31947, C2 => n39261, ZN => n36332);
   U31607 : AOI221_X1 port map( B1 => n39286, B2 => n30018, C1 => n39280, C2 =>
                           n30082, A => n36313, ZN => n36312);
   U31608 : OAI222_X1 port map( A1 => n32006, A2 => n39274, B1 => n32297, B2 =>
                           n39268, C1 => n31946, C2 => n39262, ZN => n36313);
   U31609 : AOI221_X1 port map( B1 => n39286, B2 => n30017, C1 => n39280, C2 =>
                           n30081, A => n36294, ZN => n36293);
   U31610 : OAI222_X1 port map( A1 => n32005, A2 => n39274, B1 => n32296, B2 =>
                           n39268, C1 => n31945, C2 => n39262, ZN => n36294);
   U31611 : AOI221_X1 port map( B1 => n39286, B2 => n30016, C1 => n39280, C2 =>
                           n30080, A => n36275, ZN => n36274);
   U31612 : OAI222_X1 port map( A1 => n32004, A2 => n39274, B1 => n32295, B2 =>
                           n39268, C1 => n31944, C2 => n39262, ZN => n36275);
   U31613 : AOI221_X1 port map( B1 => n39286, B2 => n30015, C1 => n39280, C2 =>
                           n30079, A => n36256, ZN => n36255);
   U31614 : OAI222_X1 port map( A1 => n32003, A2 => n39274, B1 => n32294, B2 =>
                           n39268, C1 => n31943, C2 => n39262, ZN => n36256);
   U31615 : AOI221_X1 port map( B1 => n39286, B2 => n30014, C1 => n39280, C2 =>
                           n30078, A => n36237, ZN => n36236);
   U31616 : OAI222_X1 port map( A1 => n32002, A2 => n39274, B1 => n32293, B2 =>
                           n39268, C1 => n31942, C2 => n39262, ZN => n36237);
   U31617 : AOI221_X1 port map( B1 => n39286, B2 => n30013, C1 => n39280, C2 =>
                           n30077, A => n36218, ZN => n36217);
   U31618 : OAI222_X1 port map( A1 => n32001, A2 => n39274, B1 => n32292, B2 =>
                           n39268, C1 => n31941, C2 => n39262, ZN => n36218);
   U31619 : AOI221_X1 port map( B1 => n39162, B2 => n31119, C1 => n39156, C2 =>
                           n28849, A => n37214, ZN => n37213);
   U31620 : OAI222_X1 port map( A1 => n31301, A2 => n39150, B1 => n31365, B2 =>
                           n39144, C1 => n31237, C2 => n39138, ZN => n37214);
   U31621 : AOI221_X1 port map( B1 => n39282, B2 => n30065, C1 => n39276, C2 =>
                           n30129, A => n37206, ZN => n37205);
   U31622 : OAI222_X1 port map( A1 => n32280, A2 => n39270, B1 => n32264, B2 =>
                           n39264, C1 => n32284, C2 => n39258, ZN => n37206);
   U31623 : AOI221_X1 port map( B1 => n39162, B2 => n31118, C1 => n39156, C2 =>
                           n28848, A => n37195, ZN => n37194);
   U31624 : OAI222_X1 port map( A1 => n31300, A2 => n39150, B1 => n31364, B2 =>
                           n39144, C1 => n31236, C2 => n39138, ZN => n37195);
   U31625 : AOI221_X1 port map( B1 => n39282, B2 => n30064, C1 => n39276, C2 =>
                           n30128, A => n37187, ZN => n37186);
   U31626 : OAI222_X1 port map( A1 => n32279, A2 => n39270, B1 => n32263, B2 =>
                           n39264, C1 => n32283, C2 => n39258, ZN => n37187);
   U31627 : AOI221_X1 port map( B1 => n39162, B2 => n31117, C1 => n39156, C2 =>
                           n28847, A => n37176, ZN => n37175);
   U31628 : OAI222_X1 port map( A1 => n31299, A2 => n39150, B1 => n31363, B2 =>
                           n39144, C1 => n31235, C2 => n39138, ZN => n37176);
   U31629 : AOI221_X1 port map( B1 => n39282, B2 => n30063, C1 => n39276, C2 =>
                           n30127, A => n37168, ZN => n37167);
   U31630 : OAI222_X1 port map( A1 => n32278, A2 => n39270, B1 => n32262, B2 =>
                           n39264, C1 => n32282, C2 => n39258, ZN => n37168);
   U31631 : AOI221_X1 port map( B1 => n39162, B2 => n31116, C1 => n39156, C2 =>
                           n28846, A => n37157, ZN => n37156);
   U31632 : OAI222_X1 port map( A1 => n31298, A2 => n39150, B1 => n31362, B2 =>
                           n39144, C1 => n31234, C2 => n39138, ZN => n37157);
   U31633 : AOI221_X1 port map( B1 => n39282, B2 => n30062, C1 => n39276, C2 =>
                           n30126, A => n37149, ZN => n37148);
   U31634 : OAI222_X1 port map( A1 => n32050, A2 => n39270, B1 => n32074, B2 =>
                           n39264, C1 => n31990, C2 => n39258, ZN => n37149);
   U31635 : AOI221_X1 port map( B1 => n39162, B2 => n31115, C1 => n39156, C2 =>
                           n28845, A => n37138, ZN => n37137);
   U31636 : OAI222_X1 port map( A1 => n31297, A2 => n39150, B1 => n31361, B2 =>
                           n39144, C1 => n31233, C2 => n39138, ZN => n37138);
   U31637 : AOI221_X1 port map( B1 => n39282, B2 => n30061, C1 => n39276, C2 =>
                           n30125, A => n37130, ZN => n37129);
   U31638 : OAI222_X1 port map( A1 => n32049, A2 => n39270, B1 => n32073, B2 =>
                           n39264, C1 => n31989, C2 => n39258, ZN => n37130);
   U31639 : AOI221_X1 port map( B1 => n39162, B2 => n31120, C1 => n39156, C2 =>
                           n28850, A => n37245, ZN => n37244);
   U31640 : OAI222_X1 port map( A1 => n31302, A2 => n39150, B1 => n31366, B2 =>
                           n39144, C1 => n31238, C2 => n39138, ZN => n37245);
   U31641 : AOI221_X1 port map( B1 => n39282, B2 => n30066, C1 => n39276, C2 =>
                           n30130, A => n37225, ZN => n37224);
   U31642 : OAI222_X1 port map( A1 => n32281, A2 => n39270, B1 => n32265, B2 =>
                           n39264, C1 => n32285, C2 => n39258, ZN => n37225);
   U31643 : AOI221_X1 port map( B1 => n39162, B2 => n31114, C1 => n39156, C2 =>
                           n28844, A => n37119, ZN => n37118);
   U31644 : OAI222_X1 port map( A1 => n31296, A2 => n39150, B1 => n31360, B2 =>
                           n39144, C1 => n31232, C2 => n39138, ZN => n37119);
   U31645 : AOI221_X1 port map( B1 => n39282, B2 => n30060, C1 => n39276, C2 =>
                           n30124, A => n37111, ZN => n37110);
   U31646 : OAI222_X1 port map( A1 => n32048, A2 => n39270, B1 => n32072, B2 =>
                           n39264, C1 => n31988, C2 => n39258, ZN => n37111);
   U31647 : AOI221_X1 port map( B1 => n39162, B2 => n31113, C1 => n39156, C2 =>
                           n28843, A => n37100, ZN => n37099);
   U31648 : OAI222_X1 port map( A1 => n31295, A2 => n39150, B1 => n31359, B2 =>
                           n39144, C1 => n31231, C2 => n39138, ZN => n37100);
   U31649 : AOI221_X1 port map( B1 => n39282, B2 => n30059, C1 => n39276, C2 =>
                           n30123, A => n37092, ZN => n37091);
   U31650 : OAI222_X1 port map( A1 => n32047, A2 => n39270, B1 => n32071, B2 =>
                           n39264, C1 => n31987, C2 => n39258, ZN => n37092);
   U31651 : AOI221_X1 port map( B1 => n39162, B2 => n31112, C1 => n39156, C2 =>
                           n28842, A => n37081, ZN => n37080);
   U31652 : OAI222_X1 port map( A1 => n31294, A2 => n39150, B1 => n31358, B2 =>
                           n39144, C1 => n31230, C2 => n39138, ZN => n37081);
   U31653 : AOI221_X1 port map( B1 => n39282, B2 => n30058, C1 => n39276, C2 =>
                           n30122, A => n37073, ZN => n37072);
   U31654 : OAI222_X1 port map( A1 => n32046, A2 => n39270, B1 => n32070, B2 =>
                           n39264, C1 => n31986, C2 => n39258, ZN => n37073);
   U31655 : AOI221_X1 port map( B1 => n39162, B2 => n31111, C1 => n39156, C2 =>
                           n28841, A => n37062, ZN => n37061);
   U31656 : OAI222_X1 port map( A1 => n31293, A2 => n39150, B1 => n31357, B2 =>
                           n39144, C1 => n31229, C2 => n39138, ZN => n37062);
   U31657 : AOI221_X1 port map( B1 => n39282, B2 => n30057, C1 => n39276, C2 =>
                           n30121, A => n37054, ZN => n37053);
   U31658 : OAI222_X1 port map( A1 => n32045, A2 => n39270, B1 => n32069, B2 =>
                           n39264, C1 => n31985, C2 => n39258, ZN => n37054);
   U31659 : AOI221_X1 port map( B1 => n39282, B2 => n30056, C1 => n39276, C2 =>
                           n30120, A => n37035, ZN => n37034);
   U31660 : OAI222_X1 port map( A1 => n32044, A2 => n39270, B1 => n32068, B2 =>
                           n39264, C1 => n31984, C2 => n39258, ZN => n37035);
   U31661 : AOI221_X1 port map( B1 => n39286, B2 => n30012, C1 => n39280, C2 =>
                           n30076, A => n36199, ZN => n36198);
   U31662 : OAI222_X1 port map( A1 => n32000, A2 => n39274, B1 => n32291, B2 =>
                           n39268, C1 => n31940, C2 => n39262, ZN => n36199);
   U31663 : AOI221_X1 port map( B1 => n39286, B2 => n30011, C1 => n39280, C2 =>
                           n30075, A => n36180, ZN => n36179);
   U31664 : OAI222_X1 port map( A1 => n31999, A2 => n39274, B1 => n32290, B2 =>
                           n39268, C1 => n31939, C2 => n39262, ZN => n36180);
   U31665 : AOI221_X1 port map( B1 => n39286, B2 => n30010, C1 => n39280, C2 =>
                           n30074, A => n36161, ZN => n36160);
   U31666 : OAI222_X1 port map( A1 => n31998, A2 => n39274, B1 => n32289, B2 =>
                           n39268, C1 => n31938, C2 => n39262, ZN => n36161);
   U31667 : AOI221_X1 port map( B1 => n39286, B2 => n30009, C1 => n39280, C2 =>
                           n30073, A => n36142, ZN => n36141);
   U31668 : OAI222_X1 port map( A1 => n31997, A2 => n39274, B1 => n32288, B2 =>
                           n39268, C1 => n31937, C2 => n39262, ZN => n36142);
   U31669 : AOI221_X1 port map( B1 => n39286, B2 => n30008, C1 => n39280, C2 =>
                           n30072, A => n36123, ZN => n36122);
   U31670 : OAI222_X1 port map( A1 => n31996, A2 => n39274, B1 => n32287, B2 =>
                           n39268, C1 => n31936, C2 => n39262, ZN => n36123);
   U31671 : AOI221_X1 port map( B1 => n39286, B2 => n30007, C1 => n39280, C2 =>
                           n30071, A => n36104, ZN => n36103);
   U31672 : OAI222_X1 port map( A1 => n31995, A2 => n39274, B1 => n32054, B2 =>
                           n39268, C1 => n31935, C2 => n39262, ZN => n36104);
   U31673 : AOI221_X1 port map( B1 => n39669, B2 => n31120, C1 => n39663, C2 =>
                           n28850, A => n33463, ZN => n33460);
   U31674 : OAI222_X1 port map( A1 => n31302, A2 => n39657, B1 => n31366, B2 =>
                           n39651, C1 => n31238, C2 => n39645, ZN => n33463);
   U31675 : AOI221_X1 port map( B1 => n39789, B2 => n30066, C1 => n39783, C2 =>
                           n30130, A => n33435, ZN => n33432);
   U31676 : OAI222_X1 port map( A1 => n32281, A2 => n39777, B1 => n32265, B2 =>
                           n39771, C1 => n32285, C2 => n39765, ZN => n33435);
   U31677 : AOI221_X1 port map( B1 => n39417, B2 => n31120, C1 => n39411, C2 =>
                           n28850, A => n34737, ZN => n34734);
   U31678 : OAI222_X1 port map( A1 => n31302, A2 => n39405, B1 => n31366, B2 =>
                           n39399, C1 => n31238, C2 => n39393, ZN => n34737);
   U31679 : AOI221_X1 port map( B1 => n39537, B2 => n30066, C1 => n39531, C2 =>
                           n30130, A => n34709, ZN => n34706);
   U31680 : OAI222_X1 port map( A1 => n32281, A2 => n39525, B1 => n32265, B2 =>
                           n39519, C1 => n32285, C2 => n39513, ZN => n34709);
   U31681 : AOI221_X1 port map( B1 => n39669, B2 => n31119, C1 => n39663, C2 =>
                           n28849, A => n33500, ZN => n33499);
   U31682 : OAI222_X1 port map( A1 => n31301, A2 => n39657, B1 => n31365, B2 =>
                           n39651, C1 => n31237, C2 => n39645, ZN => n33500);
   U31683 : AOI221_X1 port map( B1 => n39789, B2 => n30065, C1 => n39783, C2 =>
                           n30129, A => n33492, ZN => n33491);
   U31684 : OAI222_X1 port map( A1 => n32280, A2 => n39777, B1 => n32264, B2 =>
                           n39771, C1 => n32284, C2 => n39765, ZN => n33492);
   U31685 : AOI221_X1 port map( B1 => n39417, B2 => n31119, C1 => n39411, C2 =>
                           n28849, A => n34774, ZN => n34773);
   U31686 : OAI222_X1 port map( A1 => n31301, A2 => n39405, B1 => n31365, B2 =>
                           n39399, C1 => n31237, C2 => n39393, ZN => n34774);
   U31687 : AOI221_X1 port map( B1 => n39537, B2 => n30065, C1 => n39531, C2 =>
                           n30129, A => n34766, ZN => n34765);
   U31688 : OAI222_X1 port map( A1 => n32280, A2 => n39525, B1 => n32264, B2 =>
                           n39519, C1 => n32284, C2 => n39513, ZN => n34766);
   U31689 : AOI221_X1 port map( B1 => n39669, B2 => n31118, C1 => n39663, C2 =>
                           n28848, A => n33519, ZN => n33518);
   U31690 : OAI222_X1 port map( A1 => n31300, A2 => n39657, B1 => n31364, B2 =>
                           n39651, C1 => n31236, C2 => n39645, ZN => n33519);
   U31691 : AOI221_X1 port map( B1 => n39789, B2 => n30064, C1 => n39783, C2 =>
                           n30128, A => n33511, ZN => n33510);
   U31692 : OAI222_X1 port map( A1 => n32279, A2 => n39777, B1 => n32263, B2 =>
                           n39771, C1 => n32283, C2 => n39765, ZN => n33511);
   U31693 : AOI221_X1 port map( B1 => n39417, B2 => n31118, C1 => n39411, C2 =>
                           n28848, A => n34793, ZN => n34792);
   U31694 : OAI222_X1 port map( A1 => n31300, A2 => n39405, B1 => n31364, B2 =>
                           n39399, C1 => n31236, C2 => n39393, ZN => n34793);
   U31695 : AOI221_X1 port map( B1 => n39537, B2 => n30064, C1 => n39531, C2 =>
                           n30128, A => n34785, ZN => n34784);
   U31696 : OAI222_X1 port map( A1 => n32279, A2 => n39525, B1 => n32263, B2 =>
                           n39519, C1 => n32283, C2 => n39513, ZN => n34785);
   U31697 : AOI221_X1 port map( B1 => n39669, B2 => n31117, C1 => n39663, C2 =>
                           n28847, A => n33538, ZN => n33537);
   U31698 : OAI222_X1 port map( A1 => n31299, A2 => n39657, B1 => n31363, B2 =>
                           n39651, C1 => n31235, C2 => n39645, ZN => n33538);
   U31699 : AOI221_X1 port map( B1 => n39789, B2 => n30063, C1 => n39783, C2 =>
                           n30127, A => n33530, ZN => n33529);
   U31700 : OAI222_X1 port map( A1 => n32278, A2 => n39777, B1 => n32262, B2 =>
                           n39771, C1 => n32282, C2 => n39765, ZN => n33530);
   U31701 : AOI221_X1 port map( B1 => n39417, B2 => n31117, C1 => n39411, C2 =>
                           n28847, A => n34812, ZN => n34811);
   U31702 : OAI222_X1 port map( A1 => n31299, A2 => n39405, B1 => n31363, B2 =>
                           n39399, C1 => n31235, C2 => n39393, ZN => n34812);
   U31703 : AOI221_X1 port map( B1 => n39537, B2 => n30063, C1 => n39531, C2 =>
                           n30127, A => n34804, ZN => n34803);
   U31704 : OAI222_X1 port map( A1 => n32278, A2 => n39525, B1 => n32262, B2 =>
                           n39519, C1 => n32282, C2 => n39513, ZN => n34804);
   U31705 : AOI221_X1 port map( B1 => n39668, B2 => n31116, C1 => n39662, C2 =>
                           n28846, A => n33557, ZN => n33556);
   U31706 : OAI222_X1 port map( A1 => n31298, A2 => n39656, B1 => n31362, B2 =>
                           n39650, C1 => n31234, C2 => n39644, ZN => n33557);
   U31707 : AOI221_X1 port map( B1 => n39788, B2 => n30062, C1 => n39782, C2 =>
                           n30126, A => n33549, ZN => n33548);
   U31708 : OAI222_X1 port map( A1 => n32050, A2 => n39776, B1 => n32074, B2 =>
                           n39770, C1 => n31990, C2 => n39764, ZN => n33549);
   U31709 : AOI221_X1 port map( B1 => n39416, B2 => n31116, C1 => n39410, C2 =>
                           n28846, A => n34831, ZN => n34830);
   U31710 : OAI222_X1 port map( A1 => n31298, A2 => n39404, B1 => n31362, B2 =>
                           n39398, C1 => n31234, C2 => n39392, ZN => n34831);
   U31711 : AOI221_X1 port map( B1 => n39536, B2 => n30062, C1 => n39530, C2 =>
                           n30126, A => n34823, ZN => n34822);
   U31712 : OAI222_X1 port map( A1 => n32050, A2 => n39524, B1 => n32074, B2 =>
                           n39518, C1 => n31990, C2 => n39512, ZN => n34823);
   U31713 : AOI221_X1 port map( B1 => n39668, B2 => n31115, C1 => n39662, C2 =>
                           n28845, A => n33576, ZN => n33575);
   U31714 : OAI222_X1 port map( A1 => n31297, A2 => n39656, B1 => n31361, B2 =>
                           n39650, C1 => n31233, C2 => n39644, ZN => n33576);
   U31715 : AOI221_X1 port map( B1 => n39788, B2 => n30061, C1 => n39782, C2 =>
                           n30125, A => n33568, ZN => n33567);
   U31716 : OAI222_X1 port map( A1 => n32049, A2 => n39776, B1 => n32073, B2 =>
                           n39770, C1 => n31989, C2 => n39764, ZN => n33568);
   U31717 : AOI221_X1 port map( B1 => n39416, B2 => n31115, C1 => n39410, C2 =>
                           n28845, A => n34850, ZN => n34849);
   U31718 : OAI222_X1 port map( A1 => n31297, A2 => n39404, B1 => n31361, B2 =>
                           n39398, C1 => n31233, C2 => n39392, ZN => n34850);
   U31719 : AOI221_X1 port map( B1 => n39536, B2 => n30061, C1 => n39530, C2 =>
                           n30125, A => n34842, ZN => n34841);
   U31720 : OAI222_X1 port map( A1 => n32049, A2 => n39524, B1 => n32073, B2 =>
                           n39518, C1 => n31989, C2 => n39512, ZN => n34842);
   U31721 : AOI221_X1 port map( B1 => n39668, B2 => n31114, C1 => n39662, C2 =>
                           n28844, A => n33595, ZN => n33594);
   U31722 : OAI222_X1 port map( A1 => n31296, A2 => n39656, B1 => n31360, B2 =>
                           n39650, C1 => n31232, C2 => n39644, ZN => n33595);
   U31723 : AOI221_X1 port map( B1 => n39788, B2 => n30060, C1 => n39782, C2 =>
                           n30124, A => n33587, ZN => n33586);
   U31724 : OAI222_X1 port map( A1 => n32048, A2 => n39776, B1 => n32072, B2 =>
                           n39770, C1 => n31988, C2 => n39764, ZN => n33587);
   U31725 : AOI221_X1 port map( B1 => n39416, B2 => n31114, C1 => n39410, C2 =>
                           n28844, A => n34869, ZN => n34868);
   U31726 : OAI222_X1 port map( A1 => n31296, A2 => n39404, B1 => n31360, B2 =>
                           n39398, C1 => n31232, C2 => n39392, ZN => n34869);
   U31727 : AOI221_X1 port map( B1 => n39536, B2 => n30060, C1 => n39530, C2 =>
                           n30124, A => n34861, ZN => n34860);
   U31728 : OAI222_X1 port map( A1 => n32048, A2 => n39524, B1 => n32072, B2 =>
                           n39518, C1 => n31988, C2 => n39512, ZN => n34861);
   U31729 : AOI221_X1 port map( B1 => n39668, B2 => n31113, C1 => n39662, C2 =>
                           n28843, A => n33614, ZN => n33613);
   U31730 : OAI222_X1 port map( A1 => n31295, A2 => n39656, B1 => n31359, B2 =>
                           n39650, C1 => n31231, C2 => n39644, ZN => n33614);
   U31731 : AOI221_X1 port map( B1 => n39788, B2 => n30059, C1 => n39782, C2 =>
                           n30123, A => n33606, ZN => n33605);
   U31732 : OAI222_X1 port map( A1 => n32047, A2 => n39776, B1 => n32071, B2 =>
                           n39770, C1 => n31987, C2 => n39764, ZN => n33606);
   U31733 : AOI221_X1 port map( B1 => n39416, B2 => n31113, C1 => n39410, C2 =>
                           n28843, A => n34888, ZN => n34887);
   U31734 : OAI222_X1 port map( A1 => n31295, A2 => n39404, B1 => n31359, B2 =>
                           n39398, C1 => n31231, C2 => n39392, ZN => n34888);
   U31735 : AOI221_X1 port map( B1 => n39536, B2 => n30059, C1 => n39530, C2 =>
                           n30123, A => n34880, ZN => n34879);
   U31736 : OAI222_X1 port map( A1 => n32047, A2 => n39524, B1 => n32071, B2 =>
                           n39518, C1 => n31987, C2 => n39512, ZN => n34880);
   U31737 : AOI221_X1 port map( B1 => n39668, B2 => n31112, C1 => n39662, C2 =>
                           n28842, A => n33633, ZN => n33632);
   U31738 : OAI222_X1 port map( A1 => n31294, A2 => n39656, B1 => n31358, B2 =>
                           n39650, C1 => n31230, C2 => n39644, ZN => n33633);
   U31739 : AOI221_X1 port map( B1 => n39788, B2 => n30058, C1 => n39782, C2 =>
                           n30122, A => n33625, ZN => n33624);
   U31740 : OAI222_X1 port map( A1 => n32046, A2 => n39776, B1 => n32070, B2 =>
                           n39770, C1 => n31986, C2 => n39764, ZN => n33625);
   U31741 : AOI221_X1 port map( B1 => n39416, B2 => n31112, C1 => n39410, C2 =>
                           n28842, A => n34907, ZN => n34906);
   U31742 : OAI222_X1 port map( A1 => n31294, A2 => n39404, B1 => n31358, B2 =>
                           n39398, C1 => n31230, C2 => n39392, ZN => n34907);
   U31743 : AOI221_X1 port map( B1 => n39536, B2 => n30058, C1 => n39530, C2 =>
                           n30122, A => n34899, ZN => n34898);
   U31744 : OAI222_X1 port map( A1 => n32046, A2 => n39524, B1 => n32070, B2 =>
                           n39518, C1 => n31986, C2 => n39512, ZN => n34899);
   U31745 : AOI221_X1 port map( B1 => n39668, B2 => n31111, C1 => n39662, C2 =>
                           n28841, A => n33652, ZN => n33651);
   U31746 : OAI222_X1 port map( A1 => n31293, A2 => n39656, B1 => n31357, B2 =>
                           n39650, C1 => n31229, C2 => n39644, ZN => n33652);
   U31747 : AOI221_X1 port map( B1 => n39788, B2 => n30057, C1 => n39782, C2 =>
                           n30121, A => n33644, ZN => n33643);
   U31748 : OAI222_X1 port map( A1 => n32045, A2 => n39776, B1 => n32069, B2 =>
                           n39770, C1 => n31985, C2 => n39764, ZN => n33644);
   U31749 : AOI221_X1 port map( B1 => n39416, B2 => n31111, C1 => n39410, C2 =>
                           n28841, A => n34926, ZN => n34925);
   U31750 : OAI222_X1 port map( A1 => n31293, A2 => n39404, B1 => n31357, B2 =>
                           n39398, C1 => n31229, C2 => n39392, ZN => n34926);
   U31751 : AOI221_X1 port map( B1 => n39536, B2 => n30057, C1 => n39530, C2 =>
                           n30121, A => n34918, ZN => n34917);
   U31752 : OAI222_X1 port map( A1 => n32045, A2 => n39524, B1 => n32069, B2 =>
                           n39518, C1 => n31985, C2 => n39512, ZN => n34918);
   U31753 : AOI221_X1 port map( B1 => n39788, B2 => n30056, C1 => n39782, C2 =>
                           n30120, A => n33663, ZN => n33662);
   U31754 : OAI222_X1 port map( A1 => n32044, A2 => n39776, B1 => n32068, B2 =>
                           n39770, C1 => n31984, C2 => n39764, ZN => n33663);
   U31755 : AOI221_X1 port map( B1 => n39536, B2 => n30056, C1 => n39530, C2 =>
                           n30120, A => n34937, ZN => n34936);
   U31756 : OAI222_X1 port map( A1 => n32044, A2 => n39524, B1 => n32068, B2 =>
                           n39518, C1 => n31984, C2 => n39512, ZN => n34937);
   U31757 : AOI221_X1 port map( B1 => n39788, B2 => n30055, C1 => n39782, C2 =>
                           n30119, A => n33682, ZN => n33681);
   U31758 : OAI222_X1 port map( A1 => n32043, A2 => n39776, B1 => n32067, B2 =>
                           n39770, C1 => n31983, C2 => n39764, ZN => n33682);
   U31759 : AOI221_X1 port map( B1 => n39536, B2 => n30055, C1 => n39530, C2 =>
                           n30119, A => n34956, ZN => n34955);
   U31760 : OAI222_X1 port map( A1 => n32043, A2 => n39524, B1 => n32067, B2 =>
                           n39518, C1 => n31983, C2 => n39512, ZN => n34956);
   U31761 : AOI221_X1 port map( B1 => n39788, B2 => n30054, C1 => n39782, C2 =>
                           n30118, A => n33701, ZN => n33700);
   U31762 : OAI222_X1 port map( A1 => n32042, A2 => n39776, B1 => n32066, B2 =>
                           n39770, C1 => n31982, C2 => n39764, ZN => n33701);
   U31763 : AOI221_X1 port map( B1 => n39536, B2 => n30054, C1 => n39530, C2 =>
                           n30118, A => n34975, ZN => n34974);
   U31764 : OAI222_X1 port map( A1 => n32042, A2 => n39524, B1 => n32066, B2 =>
                           n39518, C1 => n31982, C2 => n39512, ZN => n34975);
   U31765 : AOI221_X1 port map( B1 => n39788, B2 => n30053, C1 => n39782, C2 =>
                           n30117, A => n33720, ZN => n33719);
   U31766 : OAI222_X1 port map( A1 => n32041, A2 => n39776, B1 => n32065, B2 =>
                           n39770, C1 => n31981, C2 => n39764, ZN => n33720);
   U31767 : AOI221_X1 port map( B1 => n39536, B2 => n30053, C1 => n39530, C2 =>
                           n30117, A => n34994, ZN => n34993);
   U31768 : OAI222_X1 port map( A1 => n32041, A2 => n39524, B1 => n32065, B2 =>
                           n39518, C1 => n31981, C2 => n39512, ZN => n34994);
   U31769 : AOI221_X1 port map( B1 => n39788, B2 => n30052, C1 => n39782, C2 =>
                           n30116, A => n33739, ZN => n33738);
   U31770 : OAI222_X1 port map( A1 => n32040, A2 => n39776, B1 => n32064, B2 =>
                           n39770, C1 => n31980, C2 => n39764, ZN => n33739);
   U31771 : AOI221_X1 port map( B1 => n39536, B2 => n30052, C1 => n39530, C2 =>
                           n30116, A => n35013, ZN => n35012);
   U31772 : OAI222_X1 port map( A1 => n32040, A2 => n39524, B1 => n32064, B2 =>
                           n39518, C1 => n31980, C2 => n39512, ZN => n35013);
   U31773 : AOI221_X1 port map( B1 => n39788, B2 => n30051, C1 => n39782, C2 =>
                           n30115, A => n33758, ZN => n33757);
   U31774 : OAI222_X1 port map( A1 => n32039, A2 => n39776, B1 => n32063, B2 =>
                           n39770, C1 => n31979, C2 => n39764, ZN => n33758);
   U31775 : AOI221_X1 port map( B1 => n39536, B2 => n30051, C1 => n39530, C2 =>
                           n30115, A => n35032, ZN => n35031);
   U31776 : OAI222_X1 port map( A1 => n32039, A2 => n39524, B1 => n32063, B2 =>
                           n39518, C1 => n31979, C2 => n39512, ZN => n35032);
   U31777 : AOI221_X1 port map( B1 => n39787, B2 => n30050, C1 => n39781, C2 =>
                           n30114, A => n33777, ZN => n33776);
   U31778 : OAI222_X1 port map( A1 => n32038, A2 => n39775, B1 => n32062, B2 =>
                           n39769, C1 => n31978, C2 => n39763, ZN => n33777);
   U31779 : AOI221_X1 port map( B1 => n39535, B2 => n30050, C1 => n39529, C2 =>
                           n30114, A => n35051, ZN => n35050);
   U31780 : OAI222_X1 port map( A1 => n32038, A2 => n39523, B1 => n32062, B2 =>
                           n39517, C1 => n31978, C2 => n39511, ZN => n35051);
   U31781 : AOI221_X1 port map( B1 => n39787, B2 => n30049, C1 => n39781, C2 =>
                           n30113, A => n33796, ZN => n33795);
   U31782 : OAI222_X1 port map( A1 => n32037, A2 => n39775, B1 => n32061, B2 =>
                           n39769, C1 => n31977, C2 => n39763, ZN => n33796);
   U31783 : AOI221_X1 port map( B1 => n39535, B2 => n30049, C1 => n39529, C2 =>
                           n30113, A => n35070, ZN => n35069);
   U31784 : OAI222_X1 port map( A1 => n32037, A2 => n39523, B1 => n32061, B2 =>
                           n39517, C1 => n31977, C2 => n39511, ZN => n35070);
   U31785 : AOI221_X1 port map( B1 => n39787, B2 => n30048, C1 => n39781, C2 =>
                           n30112, A => n33815, ZN => n33814);
   U31786 : OAI222_X1 port map( A1 => n32036, A2 => n39775, B1 => n32060, B2 =>
                           n39769, C1 => n31976, C2 => n39763, ZN => n33815);
   U31787 : AOI221_X1 port map( B1 => n39535, B2 => n30048, C1 => n39529, C2 =>
                           n30112, A => n35089, ZN => n35088);
   U31788 : OAI222_X1 port map( A1 => n32036, A2 => n39523, B1 => n32060, B2 =>
                           n39517, C1 => n31976, C2 => n39511, ZN => n35089);
   U31789 : AOI221_X1 port map( B1 => n39787, B2 => n30047, C1 => n39781, C2 =>
                           n30111, A => n33834, ZN => n33833);
   U31790 : OAI222_X1 port map( A1 => n32035, A2 => n39775, B1 => n32059, B2 =>
                           n39769, C1 => n31975, C2 => n39763, ZN => n33834);
   U31791 : AOI221_X1 port map( B1 => n39535, B2 => n30047, C1 => n39529, C2 =>
                           n30111, A => n35108, ZN => n35107);
   U31792 : OAI222_X1 port map( A1 => n32035, A2 => n39523, B1 => n32059, B2 =>
                           n39517, C1 => n31975, C2 => n39511, ZN => n35108);
   U31793 : AOI221_X1 port map( B1 => n39787, B2 => n30046, C1 => n39781, C2 =>
                           n30110, A => n33853, ZN => n33852);
   U31794 : OAI222_X1 port map( A1 => n32034, A2 => n39775, B1 => n32058, B2 =>
                           n39769, C1 => n31974, C2 => n39763, ZN => n33853);
   U31795 : AOI221_X1 port map( B1 => n39535, B2 => n30046, C1 => n39529, C2 =>
                           n30110, A => n35127, ZN => n35126);
   U31796 : OAI222_X1 port map( A1 => n32034, A2 => n39523, B1 => n32058, B2 =>
                           n39517, C1 => n31974, C2 => n39511, ZN => n35127);
   U31797 : AOI221_X1 port map( B1 => n39787, B2 => n30045, C1 => n39781, C2 =>
                           n30109, A => n33872, ZN => n33871);
   U31798 : OAI222_X1 port map( A1 => n32033, A2 => n39775, B1 => n32057, B2 =>
                           n39769, C1 => n31973, C2 => n39763, ZN => n33872);
   U31799 : AOI221_X1 port map( B1 => n39535, B2 => n30045, C1 => n39529, C2 =>
                           n30109, A => n35146, ZN => n35145);
   U31800 : OAI222_X1 port map( A1 => n32033, A2 => n39523, B1 => n32057, B2 =>
                           n39517, C1 => n31973, C2 => n39511, ZN => n35146);
   U31801 : AOI221_X1 port map( B1 => n39787, B2 => n30044, C1 => n39781, C2 =>
                           n30108, A => n33891, ZN => n33890);
   U31802 : OAI222_X1 port map( A1 => n32032, A2 => n39775, B1 => n32056, B2 =>
                           n39769, C1 => n31972, C2 => n39763, ZN => n33891);
   U31803 : AOI221_X1 port map( B1 => n39535, B2 => n30044, C1 => n39529, C2 =>
                           n30108, A => n35165, ZN => n35164);
   U31804 : OAI222_X1 port map( A1 => n32032, A2 => n39523, B1 => n32056, B2 =>
                           n39517, C1 => n31972, C2 => n39511, ZN => n35165);
   U31805 : AOI221_X1 port map( B1 => n39787, B2 => n30043, C1 => n39781, C2 =>
                           n30107, A => n33910, ZN => n33909);
   U31806 : OAI222_X1 port map( A1 => n32031, A2 => n39775, B1 => n32055, B2 =>
                           n39769, C1 => n31971, C2 => n39763, ZN => n33910);
   U31807 : AOI221_X1 port map( B1 => n39535, B2 => n30043, C1 => n39529, C2 =>
                           n30107, A => n35184, ZN => n35183);
   U31808 : OAI222_X1 port map( A1 => n32031, A2 => n39523, B1 => n32055, B2 =>
                           n39517, C1 => n31971, C2 => n39511, ZN => n35184);
   U31809 : AOI221_X1 port map( B1 => n39787, B2 => n30042, C1 => n39781, C2 =>
                           n30106, A => n33929, ZN => n33928);
   U31810 : OAI222_X1 port map( A1 => n32030, A2 => n39775, B1 => n32321, B2 =>
                           n39769, C1 => n31970, C2 => n39763, ZN => n33929);
   U31811 : AOI221_X1 port map( B1 => n39535, B2 => n30042, C1 => n39529, C2 =>
                           n30106, A => n35203, ZN => n35202);
   U31812 : OAI222_X1 port map( A1 => n32030, A2 => n39523, B1 => n32321, B2 =>
                           n39517, C1 => n31970, C2 => n39511, ZN => n35203);
   U31813 : AOI221_X1 port map( B1 => n39787, B2 => n30041, C1 => n39781, C2 =>
                           n30105, A => n33948, ZN => n33947);
   U31814 : OAI222_X1 port map( A1 => n32029, A2 => n39775, B1 => n32320, B2 =>
                           n39769, C1 => n31969, C2 => n39763, ZN => n33948);
   U31815 : AOI221_X1 port map( B1 => n39535, B2 => n30041, C1 => n39529, C2 =>
                           n30105, A => n35222, ZN => n35221);
   U31816 : OAI222_X1 port map( A1 => n32029, A2 => n39523, B1 => n32320, B2 =>
                           n39517, C1 => n31969, C2 => n39511, ZN => n35222);
   U31817 : AOI221_X1 port map( B1 => n39787, B2 => n30040, C1 => n39781, C2 =>
                           n30104, A => n33967, ZN => n33966);
   U31818 : OAI222_X1 port map( A1 => n32028, A2 => n39775, B1 => n32319, B2 =>
                           n39769, C1 => n31968, C2 => n39763, ZN => n33967);
   U31819 : AOI221_X1 port map( B1 => n39535, B2 => n30040, C1 => n39529, C2 =>
                           n30104, A => n35241, ZN => n35240);
   U31820 : OAI222_X1 port map( A1 => n32028, A2 => n39523, B1 => n32319, B2 =>
                           n39517, C1 => n31968, C2 => n39511, ZN => n35241);
   U31821 : AOI221_X1 port map( B1 => n39787, B2 => n30039, C1 => n39781, C2 =>
                           n30103, A => n33986, ZN => n33985);
   U31822 : OAI222_X1 port map( A1 => n32027, A2 => n39775, B1 => n32318, B2 =>
                           n39769, C1 => n31967, C2 => n39763, ZN => n33986);
   U31823 : AOI221_X1 port map( B1 => n39535, B2 => n30039, C1 => n39529, C2 =>
                           n30103, A => n35260, ZN => n35259);
   U31824 : OAI222_X1 port map( A1 => n32027, A2 => n39523, B1 => n32318, B2 =>
                           n39517, C1 => n31967, C2 => n39511, ZN => n35260);
   U31825 : AOI221_X1 port map( B1 => n39786, B2 => n30038, C1 => n39780, C2 =>
                           n30102, A => n34005, ZN => n34004);
   U31826 : OAI222_X1 port map( A1 => n32026, A2 => n39774, B1 => n32317, B2 =>
                           n39768, C1 => n31966, C2 => n39762, ZN => n34005);
   U31827 : AOI221_X1 port map( B1 => n39534, B2 => n30038, C1 => n39528, C2 =>
                           n30102, A => n35279, ZN => n35278);
   U31828 : OAI222_X1 port map( A1 => n32026, A2 => n39522, B1 => n32317, B2 =>
                           n39516, C1 => n31966, C2 => n39510, ZN => n35279);
   U31829 : AOI221_X1 port map( B1 => n39786, B2 => n30037, C1 => n39780, C2 =>
                           n30101, A => n34024, ZN => n34023);
   U31830 : OAI222_X1 port map( A1 => n32025, A2 => n39774, B1 => n32316, B2 =>
                           n39768, C1 => n31965, C2 => n39762, ZN => n34024);
   U31831 : AOI221_X1 port map( B1 => n39534, B2 => n30037, C1 => n39528, C2 =>
                           n30101, A => n35298, ZN => n35297);
   U31832 : OAI222_X1 port map( A1 => n32025, A2 => n39522, B1 => n32316, B2 =>
                           n39516, C1 => n31965, C2 => n39510, ZN => n35298);
   U31833 : AOI221_X1 port map( B1 => n39786, B2 => n30036, C1 => n39780, C2 =>
                           n30100, A => n34043, ZN => n34042);
   U31834 : OAI222_X1 port map( A1 => n32024, A2 => n39774, B1 => n32315, B2 =>
                           n39768, C1 => n31964, C2 => n39762, ZN => n34043);
   U31835 : AOI221_X1 port map( B1 => n39534, B2 => n30036, C1 => n39528, C2 =>
                           n30100, A => n35317, ZN => n35316);
   U31836 : OAI222_X1 port map( A1 => n32024, A2 => n39522, B1 => n32315, B2 =>
                           n39516, C1 => n31964, C2 => n39510, ZN => n35317);
   U31837 : AOI221_X1 port map( B1 => n39786, B2 => n30035, C1 => n39780, C2 =>
                           n30099, A => n34062, ZN => n34061);
   U31838 : OAI222_X1 port map( A1 => n32023, A2 => n39774, B1 => n32314, B2 =>
                           n39768, C1 => n31963, C2 => n39762, ZN => n34062);
   U31839 : AOI221_X1 port map( B1 => n39534, B2 => n30035, C1 => n39528, C2 =>
                           n30099, A => n35336, ZN => n35335);
   U31840 : OAI222_X1 port map( A1 => n32023, A2 => n39522, B1 => n32314, B2 =>
                           n39516, C1 => n31963, C2 => n39510, ZN => n35336);
   U31841 : AOI221_X1 port map( B1 => n39786, B2 => n30034, C1 => n39780, C2 =>
                           n30098, A => n34081, ZN => n34080);
   U31842 : OAI222_X1 port map( A1 => n32022, A2 => n39774, B1 => n32313, B2 =>
                           n39768, C1 => n31962, C2 => n39762, ZN => n34081);
   U31843 : AOI221_X1 port map( B1 => n39534, B2 => n30034, C1 => n39528, C2 =>
                           n30098, A => n35355, ZN => n35354);
   U31844 : OAI222_X1 port map( A1 => n32022, A2 => n39522, B1 => n32313, B2 =>
                           n39516, C1 => n31962, C2 => n39510, ZN => n35355);
   U31845 : AOI221_X1 port map( B1 => n39786, B2 => n30033, C1 => n39780, C2 =>
                           n30097, A => n34100, ZN => n34099);
   U31846 : OAI222_X1 port map( A1 => n32021, A2 => n39774, B1 => n32312, B2 =>
                           n39768, C1 => n31961, C2 => n39762, ZN => n34100);
   U31847 : AOI221_X1 port map( B1 => n39534, B2 => n30033, C1 => n39528, C2 =>
                           n30097, A => n35374, ZN => n35373);
   U31848 : OAI222_X1 port map( A1 => n32021, A2 => n39522, B1 => n32312, B2 =>
                           n39516, C1 => n31961, C2 => n39510, ZN => n35374);
   U31849 : AOI221_X1 port map( B1 => n39786, B2 => n30032, C1 => n39780, C2 =>
                           n30096, A => n34119, ZN => n34118);
   U31850 : OAI222_X1 port map( A1 => n32020, A2 => n39774, B1 => n32311, B2 =>
                           n39768, C1 => n31960, C2 => n39762, ZN => n34119);
   U31851 : AOI221_X1 port map( B1 => n39534, B2 => n30032, C1 => n39528, C2 =>
                           n30096, A => n35393, ZN => n35392);
   U31852 : OAI222_X1 port map( A1 => n32020, A2 => n39522, B1 => n32311, B2 =>
                           n39516, C1 => n31960, C2 => n39510, ZN => n35393);
   U31853 : AOI221_X1 port map( B1 => n39786, B2 => n30031, C1 => n39780, C2 =>
                           n30095, A => n34138, ZN => n34137);
   U31854 : OAI222_X1 port map( A1 => n32019, A2 => n39774, B1 => n32310, B2 =>
                           n39768, C1 => n31959, C2 => n39762, ZN => n34138);
   U31855 : AOI221_X1 port map( B1 => n39534, B2 => n30031, C1 => n39528, C2 =>
                           n30095, A => n35412, ZN => n35411);
   U31856 : OAI222_X1 port map( A1 => n32019, A2 => n39522, B1 => n32310, B2 =>
                           n39516, C1 => n31959, C2 => n39510, ZN => n35412);
   U31857 : AOI221_X1 port map( B1 => n39786, B2 => n30030, C1 => n39780, C2 =>
                           n30094, A => n34157, ZN => n34156);
   U31858 : OAI222_X1 port map( A1 => n32018, A2 => n39774, B1 => n32309, B2 =>
                           n39768, C1 => n31958, C2 => n39762, ZN => n34157);
   U31859 : AOI221_X1 port map( B1 => n39534, B2 => n30030, C1 => n39528, C2 =>
                           n30094, A => n35431, ZN => n35430);
   U31860 : OAI222_X1 port map( A1 => n32018, A2 => n39522, B1 => n32309, B2 =>
                           n39516, C1 => n31958, C2 => n39510, ZN => n35431);
   U31861 : AOI221_X1 port map( B1 => n39786, B2 => n30029, C1 => n39780, C2 =>
                           n30093, A => n34176, ZN => n34175);
   U31862 : OAI222_X1 port map( A1 => n32017, A2 => n39774, B1 => n32308, B2 =>
                           n39768, C1 => n31957, C2 => n39762, ZN => n34176);
   U31863 : AOI221_X1 port map( B1 => n39534, B2 => n30029, C1 => n39528, C2 =>
                           n30093, A => n35450, ZN => n35449);
   U31864 : OAI222_X1 port map( A1 => n32017, A2 => n39522, B1 => n32308, B2 =>
                           n39516, C1 => n31957, C2 => n39510, ZN => n35450);
   U31865 : AOI221_X1 port map( B1 => n39786, B2 => n30028, C1 => n39780, C2 =>
                           n30092, A => n34195, ZN => n34194);
   U31866 : OAI222_X1 port map( A1 => n32016, A2 => n39774, B1 => n32307, B2 =>
                           n39768, C1 => n31956, C2 => n39762, ZN => n34195);
   U31867 : AOI221_X1 port map( B1 => n39534, B2 => n30028, C1 => n39528, C2 =>
                           n30092, A => n35469, ZN => n35468);
   U31868 : OAI222_X1 port map( A1 => n32016, A2 => n39522, B1 => n32307, B2 =>
                           n39516, C1 => n31956, C2 => n39510, ZN => n35469);
   U31869 : AOI221_X1 port map( B1 => n39786, B2 => n30027, C1 => n39780, C2 =>
                           n30091, A => n34214, ZN => n34213);
   U31870 : OAI222_X1 port map( A1 => n32015, A2 => n39774, B1 => n32306, B2 =>
                           n39768, C1 => n31955, C2 => n39762, ZN => n34214);
   U31871 : AOI221_X1 port map( B1 => n39534, B2 => n30027, C1 => n39528, C2 =>
                           n30091, A => n35488, ZN => n35487);
   U31872 : OAI222_X1 port map( A1 => n32015, A2 => n39522, B1 => n32306, B2 =>
                           n39516, C1 => n31955, C2 => n39510, ZN => n35488);
   U31873 : AOI221_X1 port map( B1 => n39785, B2 => n30026, C1 => n39779, C2 =>
                           n30090, A => n34233, ZN => n34232);
   U31874 : OAI222_X1 port map( A1 => n32014, A2 => n39773, B1 => n32305, B2 =>
                           n39767, C1 => n31954, C2 => n39761, ZN => n34233);
   U31875 : AOI221_X1 port map( B1 => n39533, B2 => n30026, C1 => n39527, C2 =>
                           n30090, A => n35507, ZN => n35506);
   U31876 : OAI222_X1 port map( A1 => n32014, A2 => n39521, B1 => n32305, B2 =>
                           n39515, C1 => n31954, C2 => n39509, ZN => n35507);
   U31877 : AOI221_X1 port map( B1 => n39785, B2 => n30025, C1 => n39779, C2 =>
                           n30089, A => n34252, ZN => n34251);
   U31878 : OAI222_X1 port map( A1 => n32013, A2 => n39773, B1 => n32304, B2 =>
                           n39767, C1 => n31953, C2 => n39761, ZN => n34252);
   U31879 : AOI221_X1 port map( B1 => n39533, B2 => n30025, C1 => n39527, C2 =>
                           n30089, A => n35526, ZN => n35525);
   U31880 : OAI222_X1 port map( A1 => n32013, A2 => n39521, B1 => n32304, B2 =>
                           n39515, C1 => n31953, C2 => n39509, ZN => n35526);
   U31881 : AOI221_X1 port map( B1 => n39785, B2 => n30024, C1 => n39779, C2 =>
                           n30088, A => n34271, ZN => n34270);
   U31882 : OAI222_X1 port map( A1 => n32012, A2 => n39773, B1 => n32303, B2 =>
                           n39767, C1 => n31952, C2 => n39761, ZN => n34271);
   U31883 : AOI221_X1 port map( B1 => n39533, B2 => n30024, C1 => n39527, C2 =>
                           n30088, A => n35545, ZN => n35544);
   U31884 : OAI222_X1 port map( A1 => n32012, A2 => n39521, B1 => n32303, B2 =>
                           n39515, C1 => n31952, C2 => n39509, ZN => n35545);
   U31885 : AOI221_X1 port map( B1 => n39785, B2 => n30023, C1 => n39779, C2 =>
                           n30087, A => n34290, ZN => n34289);
   U31886 : OAI222_X1 port map( A1 => n32011, A2 => n39773, B1 => n32302, B2 =>
                           n39767, C1 => n31951, C2 => n39761, ZN => n34290);
   U31887 : AOI221_X1 port map( B1 => n39533, B2 => n30023, C1 => n39527, C2 =>
                           n30087, A => n35564, ZN => n35563);
   U31888 : OAI222_X1 port map( A1 => n32011, A2 => n39521, B1 => n32302, B2 =>
                           n39515, C1 => n31951, C2 => n39509, ZN => n35564);
   U31889 : AOI221_X1 port map( B1 => n39785, B2 => n30022, C1 => n39779, C2 =>
                           n30086, A => n34309, ZN => n34308);
   U31890 : OAI222_X1 port map( A1 => n32010, A2 => n39773, B1 => n32301, B2 =>
                           n39767, C1 => n31950, C2 => n39761, ZN => n34309);
   U31891 : AOI221_X1 port map( B1 => n39533, B2 => n30022, C1 => n39527, C2 =>
                           n30086, A => n35583, ZN => n35582);
   U31892 : OAI222_X1 port map( A1 => n32010, A2 => n39521, B1 => n32301, B2 =>
                           n39515, C1 => n31950, C2 => n39509, ZN => n35583);
   U31893 : AOI221_X1 port map( B1 => n39785, B2 => n30021, C1 => n39779, C2 =>
                           n30085, A => n34328, ZN => n34327);
   U31894 : OAI222_X1 port map( A1 => n32009, A2 => n39773, B1 => n32300, B2 =>
                           n39767, C1 => n31949, C2 => n39761, ZN => n34328);
   U31895 : AOI221_X1 port map( B1 => n39533, B2 => n30021, C1 => n39527, C2 =>
                           n30085, A => n35602, ZN => n35601);
   U31896 : OAI222_X1 port map( A1 => n32009, A2 => n39521, B1 => n32300, B2 =>
                           n39515, C1 => n31949, C2 => n39509, ZN => n35602);
   U31897 : AOI221_X1 port map( B1 => n39785, B2 => n30020, C1 => n39779, C2 =>
                           n30084, A => n34347, ZN => n34346);
   U31898 : OAI222_X1 port map( A1 => n32008, A2 => n39773, B1 => n32299, B2 =>
                           n39767, C1 => n31948, C2 => n39761, ZN => n34347);
   U31899 : AOI221_X1 port map( B1 => n39533, B2 => n30020, C1 => n39527, C2 =>
                           n30084, A => n35621, ZN => n35620);
   U31900 : OAI222_X1 port map( A1 => n32008, A2 => n39521, B1 => n32299, B2 =>
                           n39515, C1 => n31948, C2 => n39509, ZN => n35621);
   U31901 : AOI221_X1 port map( B1 => n39785, B2 => n30019, C1 => n39779, C2 =>
                           n30083, A => n34366, ZN => n34365);
   U31902 : OAI222_X1 port map( A1 => n32007, A2 => n39773, B1 => n32298, B2 =>
                           n39767, C1 => n31947, C2 => n39761, ZN => n34366);
   U31903 : AOI221_X1 port map( B1 => n39533, B2 => n30019, C1 => n39527, C2 =>
                           n30083, A => n35640, ZN => n35639);
   U31904 : OAI222_X1 port map( A1 => n32007, A2 => n39521, B1 => n32298, B2 =>
                           n39515, C1 => n31947, C2 => n39509, ZN => n35640);
   U31905 : AOI221_X1 port map( B1 => n39785, B2 => n30018, C1 => n39779, C2 =>
                           n30082, A => n34385, ZN => n34384);
   U31906 : OAI222_X1 port map( A1 => n32006, A2 => n39773, B1 => n32297, B2 =>
                           n39767, C1 => n31946, C2 => n39761, ZN => n34385);
   U31907 : AOI221_X1 port map( B1 => n39533, B2 => n30018, C1 => n39527, C2 =>
                           n30082, A => n35659, ZN => n35658);
   U31908 : OAI222_X1 port map( A1 => n32006, A2 => n39521, B1 => n32297, B2 =>
                           n39515, C1 => n31946, C2 => n39509, ZN => n35659);
   U31909 : AOI221_X1 port map( B1 => n39785, B2 => n30017, C1 => n39779, C2 =>
                           n30081, A => n34404, ZN => n34403);
   U31910 : OAI222_X1 port map( A1 => n32005, A2 => n39773, B1 => n32296, B2 =>
                           n39767, C1 => n31945, C2 => n39761, ZN => n34404);
   U31911 : AOI221_X1 port map( B1 => n39533, B2 => n30017, C1 => n39527, C2 =>
                           n30081, A => n35678, ZN => n35677);
   U31912 : OAI222_X1 port map( A1 => n32005, A2 => n39521, B1 => n32296, B2 =>
                           n39515, C1 => n31945, C2 => n39509, ZN => n35678);
   U31913 : AOI221_X1 port map( B1 => n39785, B2 => n30016, C1 => n39779, C2 =>
                           n30080, A => n34423, ZN => n34422);
   U31914 : OAI222_X1 port map( A1 => n32004, A2 => n39773, B1 => n32295, B2 =>
                           n39767, C1 => n31944, C2 => n39761, ZN => n34423);
   U31915 : AOI221_X1 port map( B1 => n39533, B2 => n30016, C1 => n39527, C2 =>
                           n30080, A => n35697, ZN => n35696);
   U31916 : OAI222_X1 port map( A1 => n32004, A2 => n39521, B1 => n32295, B2 =>
                           n39515, C1 => n31944, C2 => n39509, ZN => n35697);
   U31917 : AOI221_X1 port map( B1 => n39785, B2 => n30015, C1 => n39779, C2 =>
                           n30079, A => n34442, ZN => n34441);
   U31918 : OAI222_X1 port map( A1 => n32003, A2 => n39773, B1 => n32294, B2 =>
                           n39767, C1 => n31943, C2 => n39761, ZN => n34442);
   U31919 : AOI221_X1 port map( B1 => n39533, B2 => n30015, C1 => n39527, C2 =>
                           n30079, A => n35716, ZN => n35715);
   U31920 : OAI222_X1 port map( A1 => n32003, A2 => n39521, B1 => n32294, B2 =>
                           n39515, C1 => n31943, C2 => n39509, ZN => n35716);
   U31921 : AOI221_X1 port map( B1 => n39784, B2 => n30014, C1 => n39778, C2 =>
                           n30078, A => n34461, ZN => n34460);
   U31922 : OAI222_X1 port map( A1 => n32002, A2 => n39772, B1 => n32293, B2 =>
                           n39766, C1 => n31942, C2 => n39760, ZN => n34461);
   U31923 : AOI221_X1 port map( B1 => n39532, B2 => n30014, C1 => n39526, C2 =>
                           n30078, A => n35735, ZN => n35734);
   U31924 : OAI222_X1 port map( A1 => n32002, A2 => n39520, B1 => n32293, B2 =>
                           n39514, C1 => n31942, C2 => n39508, ZN => n35735);
   U31925 : AOI221_X1 port map( B1 => n39784, B2 => n30013, C1 => n39778, C2 =>
                           n30077, A => n34480, ZN => n34479);
   U31926 : OAI222_X1 port map( A1 => n32001, A2 => n39772, B1 => n32292, B2 =>
                           n39766, C1 => n31941, C2 => n39760, ZN => n34480);
   U31927 : AOI221_X1 port map( B1 => n39532, B2 => n30013, C1 => n39526, C2 =>
                           n30077, A => n35754, ZN => n35753);
   U31928 : OAI222_X1 port map( A1 => n32001, A2 => n39520, B1 => n32292, B2 =>
                           n39514, C1 => n31941, C2 => n39508, ZN => n35754);
   U31929 : AOI221_X1 port map( B1 => n39784, B2 => n30012, C1 => n39778, C2 =>
                           n30076, A => n34499, ZN => n34498);
   U31930 : OAI222_X1 port map( A1 => n32000, A2 => n39772, B1 => n32291, B2 =>
                           n39766, C1 => n31940, C2 => n39760, ZN => n34499);
   U31931 : AOI221_X1 port map( B1 => n39532, B2 => n30012, C1 => n39526, C2 =>
                           n30076, A => n35773, ZN => n35772);
   U31932 : OAI222_X1 port map( A1 => n32000, A2 => n39520, B1 => n32291, B2 =>
                           n39514, C1 => n31940, C2 => n39508, ZN => n35773);
   U31933 : AOI221_X1 port map( B1 => n39784, B2 => n30011, C1 => n39778, C2 =>
                           n30075, A => n34518, ZN => n34517);
   U31934 : OAI222_X1 port map( A1 => n31999, A2 => n39772, B1 => n32290, B2 =>
                           n39766, C1 => n31939, C2 => n39760, ZN => n34518);
   U31935 : AOI221_X1 port map( B1 => n39532, B2 => n30011, C1 => n39526, C2 =>
                           n30075, A => n35792, ZN => n35791);
   U31936 : OAI222_X1 port map( A1 => n31999, A2 => n39520, B1 => n32290, B2 =>
                           n39514, C1 => n31939, C2 => n39508, ZN => n35792);
   U31937 : AOI221_X1 port map( B1 => n39784, B2 => n30010, C1 => n39778, C2 =>
                           n30074, A => n34537, ZN => n34536);
   U31938 : OAI222_X1 port map( A1 => n31998, A2 => n39772, B1 => n32289, B2 =>
                           n39766, C1 => n31938, C2 => n39760, ZN => n34537);
   U31939 : AOI221_X1 port map( B1 => n39532, B2 => n30010, C1 => n39526, C2 =>
                           n30074, A => n35811, ZN => n35810);
   U31940 : OAI222_X1 port map( A1 => n31998, A2 => n39520, B1 => n32289, B2 =>
                           n39514, C1 => n31938, C2 => n39508, ZN => n35811);
   U31941 : AOI221_X1 port map( B1 => n39784, B2 => n30009, C1 => n39778, C2 =>
                           n30073, A => n34556, ZN => n34555);
   U31942 : OAI222_X1 port map( A1 => n31997, A2 => n39772, B1 => n32288, B2 =>
                           n39766, C1 => n31937, C2 => n39760, ZN => n34556);
   U31943 : AOI221_X1 port map( B1 => n39532, B2 => n30009, C1 => n39526, C2 =>
                           n30073, A => n35830, ZN => n35829);
   U31944 : OAI222_X1 port map( A1 => n31997, A2 => n39520, B1 => n32288, B2 =>
                           n39514, C1 => n31937, C2 => n39508, ZN => n35830);
   U31945 : AOI221_X1 port map( B1 => n39784, B2 => n30008, C1 => n39778, C2 =>
                           n30072, A => n34575, ZN => n34574);
   U31946 : OAI222_X1 port map( A1 => n31996, A2 => n39772, B1 => n32287, B2 =>
                           n39766, C1 => n31936, C2 => n39760, ZN => n34575);
   U31947 : AOI221_X1 port map( B1 => n39532, B2 => n30008, C1 => n39526, C2 =>
                           n30072, A => n35849, ZN => n35848);
   U31948 : OAI222_X1 port map( A1 => n31996, A2 => n39520, B1 => n32287, B2 =>
                           n39514, C1 => n31936, C2 => n39508, ZN => n35849);
   U31949 : AOI221_X1 port map( B1 => n39784, B2 => n30007, C1 => n39778, C2 =>
                           n30071, A => n34594, ZN => n34593);
   U31950 : OAI222_X1 port map( A1 => n31995, A2 => n39772, B1 => n32054, B2 =>
                           n39766, C1 => n31935, C2 => n39760, ZN => n34594);
   U31951 : AOI221_X1 port map( B1 => n39532, B2 => n30007, C1 => n39526, C2 =>
                           n30071, A => n35868, ZN => n35867);
   U31952 : OAI222_X1 port map( A1 => n31995, A2 => n39520, B1 => n32054, B2 =>
                           n39514, C1 => n31935, C2 => n39508, ZN => n35868);
   U31953 : AOI221_X1 port map( B1 => n39784, B2 => n30006, C1 => n39778, C2 =>
                           n30070, A => n34613, ZN => n34612);
   U31954 : OAI222_X1 port map( A1 => n31994, A2 => n39772, B1 => n32286, B2 =>
                           n39766, C1 => n31934, C2 => n39760, ZN => n34613);
   U31955 : AOI221_X1 port map( B1 => n39532, B2 => n30006, C1 => n39526, C2 =>
                           n30070, A => n35887, ZN => n35886);
   U31956 : OAI222_X1 port map( A1 => n31994, A2 => n39520, B1 => n32286, B2 =>
                           n39514, C1 => n31934, C2 => n39508, ZN => n35887);
   U31957 : AOI221_X1 port map( B1 => n39784, B2 => n30005, C1 => n39778, C2 =>
                           n30069, A => n34632, ZN => n34631);
   U31958 : OAI222_X1 port map( A1 => n31993, A2 => n39772, B1 => n32053, B2 =>
                           n39766, C1 => n31933, C2 => n39760, ZN => n34632);
   U31959 : AOI221_X1 port map( B1 => n39532, B2 => n30005, C1 => n39526, C2 =>
                           n30069, A => n35906, ZN => n35905);
   U31960 : OAI222_X1 port map( A1 => n31993, A2 => n39520, B1 => n32053, B2 =>
                           n39514, C1 => n31933, C2 => n39508, ZN => n35906);
   U31961 : AOI221_X1 port map( B1 => n39784, B2 => n30004, C1 => n39778, C2 =>
                           n30068, A => n34651, ZN => n34650);
   U31962 : OAI222_X1 port map( A1 => n31992, A2 => n39772, B1 => n32052, B2 =>
                           n39766, C1 => n31932, C2 => n39760, ZN => n34651);
   U31963 : AOI221_X1 port map( B1 => n39532, B2 => n30004, C1 => n39526, C2 =>
                           n30068, A => n35925, ZN => n35924);
   U31964 : OAI222_X1 port map( A1 => n31992, A2 => n39520, B1 => n32052, B2 =>
                           n39514, C1 => n31932, C2 => n39508, ZN => n35925);
   U31965 : AOI221_X1 port map( B1 => n39784, B2 => n30003, C1 => n39778, C2 =>
                           n30067, A => n34670, ZN => n34669);
   U31966 : OAI222_X1 port map( A1 => n31991, A2 => n39772, B1 => n32051, B2 =>
                           n39766, C1 => n31931, C2 => n39760, ZN => n34670);
   U31967 : AOI221_X1 port map( B1 => n39532, B2 => n30003, C1 => n39526, C2 =>
                           n30067, A => n35944, ZN => n35943);
   U31968 : OAI222_X1 port map( A1 => n31991, A2 => n39520, B1 => n32051, B2 =>
                           n39514, C1 => n31931, C2 => n39508, ZN => n35944);
   U31969 : AOI221_X1 port map( B1 => n39252, B2 => n29735, C1 => n39246, C2 =>
                           n29799, A => n37017, ZN => n37014);
   U31970 : OAI222_X1 port map( A1 => n31863, A2 => n39240, B1 => n31923, B2 =>
                           n39234, C1 => n31803, C2 => n39228, ZN => n37017);
   U31971 : AOI221_X1 port map( B1 => n39253, B2 => n29734, C1 => n39247, C2 =>
                           n29798, A => n36998, ZN => n36995);
   U31972 : OAI222_X1 port map( A1 => n31862, A2 => n39241, B1 => n31922, B2 =>
                           n39235, C1 => n31802, C2 => n39229, ZN => n36998);
   U31973 : AOI221_X1 port map( B1 => n39253, B2 => n29733, C1 => n39247, C2 =>
                           n29797, A => n36979, ZN => n36976);
   U31974 : OAI222_X1 port map( A1 => n31861, A2 => n39241, B1 => n31921, B2 =>
                           n39235, C1 => n31801, C2 => n39229, ZN => n36979);
   U31975 : AOI221_X1 port map( B1 => n39253, B2 => n29732, C1 => n39247, C2 =>
                           n29796, A => n36960, ZN => n36957);
   U31976 : OAI222_X1 port map( A1 => n31860, A2 => n39241, B1 => n31920, B2 =>
                           n39235, C1 => n31800, C2 => n39229, ZN => n36960);
   U31977 : AOI221_X1 port map( B1 => n39253, B2 => n29731, C1 => n39247, C2 =>
                           n29795, A => n36941, ZN => n36938);
   U31978 : OAI222_X1 port map( A1 => n31859, A2 => n39241, B1 => n31919, B2 =>
                           n39235, C1 => n31799, C2 => n39229, ZN => n36941);
   U31979 : AOI221_X1 port map( B1 => n39253, B2 => n29730, C1 => n39247, C2 =>
                           n29794, A => n36922, ZN => n36919);
   U31980 : OAI222_X1 port map( A1 => n31858, A2 => n39241, B1 => n31918, B2 =>
                           n39235, C1 => n31798, C2 => n39229, ZN => n36922);
   U31981 : AOI221_X1 port map( B1 => n39253, B2 => n29729, C1 => n39247, C2 =>
                           n29793, A => n36903, ZN => n36900);
   U31982 : OAI222_X1 port map( A1 => n31857, A2 => n39241, B1 => n31917, B2 =>
                           n39235, C1 => n31797, C2 => n39229, ZN => n36903);
   U31983 : AOI221_X1 port map( B1 => n39253, B2 => n29728, C1 => n39247, C2 =>
                           n29792, A => n36884, ZN => n36881);
   U31984 : OAI222_X1 port map( A1 => n31856, A2 => n39241, B1 => n31916, B2 =>
                           n39235, C1 => n31796, C2 => n39229, ZN => n36884);
   U31985 : AOI221_X1 port map( B1 => n39253, B2 => n29727, C1 => n39247, C2 =>
                           n29791, A => n36865, ZN => n36862);
   U31986 : OAI222_X1 port map( A1 => n31855, A2 => n39241, B1 => n31915, B2 =>
                           n39235, C1 => n31795, C2 => n39229, ZN => n36865);
   U31987 : AOI221_X1 port map( B1 => n39253, B2 => n29726, C1 => n39247, C2 =>
                           n29790, A => n36846, ZN => n36843);
   U31988 : OAI222_X1 port map( A1 => n31854, A2 => n39241, B1 => n31914, B2 =>
                           n39235, C1 => n31794, C2 => n39229, ZN => n36846);
   U31989 : AOI221_X1 port map( B1 => n39253, B2 => n29725, C1 => n39247, C2 =>
                           n29789, A => n36827, ZN => n36824);
   U31990 : OAI222_X1 port map( A1 => n31853, A2 => n39241, B1 => n31913, B2 =>
                           n39235, C1 => n31793, C2 => n39229, ZN => n36827);
   U31991 : AOI221_X1 port map( B1 => n39253, B2 => n29724, C1 => n39247, C2 =>
                           n29788, A => n36808, ZN => n36805);
   U31992 : OAI222_X1 port map( A1 => n31852, A2 => n39241, B1 => n31912, B2 =>
                           n39235, C1 => n31792, C2 => n39229, ZN => n36808);
   U31993 : AOI221_X1 port map( B1 => n39253, B2 => n29723, C1 => n39247, C2 =>
                           n29787, A => n36789, ZN => n36786);
   U31994 : OAI222_X1 port map( A1 => n31851, A2 => n39241, B1 => n31911, B2 =>
                           n39235, C1 => n31791, C2 => n39229, ZN => n36789);
   U31995 : AOI221_X1 port map( B1 => n39254, B2 => n29722, C1 => n39248, C2 =>
                           n29786, A => n36770, ZN => n36767);
   U31996 : OAI222_X1 port map( A1 => n31850, A2 => n39242, B1 => n31910, B2 =>
                           n39236, C1 => n31790, C2 => n39230, ZN => n36770);
   U31997 : AOI221_X1 port map( B1 => n39254, B2 => n29721, C1 => n39248, C2 =>
                           n29785, A => n36751, ZN => n36748);
   U31998 : OAI222_X1 port map( A1 => n31849, A2 => n39242, B1 => n31909, B2 =>
                           n39236, C1 => n31789, C2 => n39230, ZN => n36751);
   U31999 : AOI221_X1 port map( B1 => n39254, B2 => n29720, C1 => n39248, C2 =>
                           n29784, A => n36732, ZN => n36729);
   U32000 : OAI222_X1 port map( A1 => n31848, A2 => n39242, B1 => n31908, B2 =>
                           n39236, C1 => n31788, C2 => n39230, ZN => n36732);
   U32001 : AOI221_X1 port map( B1 => n39254, B2 => n29719, C1 => n39248, C2 =>
                           n29783, A => n36713, ZN => n36710);
   U32002 : OAI222_X1 port map( A1 => n31847, A2 => n39242, B1 => n31907, B2 =>
                           n39236, C1 => n31787, C2 => n39230, ZN => n36713);
   U32003 : AOI221_X1 port map( B1 => n39254, B2 => n29718, C1 => n39248, C2 =>
                           n29782, A => n36694, ZN => n36691);
   U32004 : OAI222_X1 port map( A1 => n31846, A2 => n39242, B1 => n31906, B2 =>
                           n39236, C1 => n31786, C2 => n39230, ZN => n36694);
   U32005 : AOI221_X1 port map( B1 => n39254, B2 => n29717, C1 => n39248, C2 =>
                           n29781, A => n36675, ZN => n36672);
   U32006 : OAI222_X1 port map( A1 => n31845, A2 => n39242, B1 => n31905, B2 =>
                           n39236, C1 => n31785, C2 => n39230, ZN => n36675);
   U32007 : AOI221_X1 port map( B1 => n39254, B2 => n29716, C1 => n39248, C2 =>
                           n29780, A => n36656, ZN => n36653);
   U32008 : OAI222_X1 port map( A1 => n31844, A2 => n39242, B1 => n31904, B2 =>
                           n39236, C1 => n31784, C2 => n39230, ZN => n36656);
   U32009 : AOI221_X1 port map( B1 => n39254, B2 => n29715, C1 => n39248, C2 =>
                           n29779, A => n36637, ZN => n36634);
   U32010 : OAI222_X1 port map( A1 => n31843, A2 => n39242, B1 => n31903, B2 =>
                           n39236, C1 => n31783, C2 => n39230, ZN => n36637);
   U32011 : AOI221_X1 port map( B1 => n39254, B2 => n29714, C1 => n39248, C2 =>
                           n29778, A => n36618, ZN => n36615);
   U32012 : OAI222_X1 port map( A1 => n31842, A2 => n39242, B1 => n31902, B2 =>
                           n39236, C1 => n31782, C2 => n39230, ZN => n36618);
   U32013 : AOI221_X1 port map( B1 => n39254, B2 => n29713, C1 => n39248, C2 =>
                           n29777, A => n36599, ZN => n36596);
   U32014 : OAI222_X1 port map( A1 => n31841, A2 => n39242, B1 => n31901, B2 =>
                           n39236, C1 => n31781, C2 => n39230, ZN => n36599);
   U32015 : AOI221_X1 port map( B1 => n39254, B2 => n29712, C1 => n39248, C2 =>
                           n29776, A => n36580, ZN => n36577);
   U32016 : OAI222_X1 port map( A1 => n31840, A2 => n39242, B1 => n31900, B2 =>
                           n39236, C1 => n31780, C2 => n39230, ZN => n36580);
   U32017 : AOI221_X1 port map( B1 => n39254, B2 => n29711, C1 => n39248, C2 =>
                           n29775, A => n36561, ZN => n36558);
   U32018 : OAI222_X1 port map( A1 => n31839, A2 => n39242, B1 => n31899, B2 =>
                           n39236, C1 => n31779, C2 => n39230, ZN => n36561);
   U32019 : AOI221_X1 port map( B1 => n39255, B2 => n29710, C1 => n39249, C2 =>
                           n29774, A => n36542, ZN => n36539);
   U32020 : OAI222_X1 port map( A1 => n31838, A2 => n39243, B1 => n31898, B2 =>
                           n39237, C1 => n31778, C2 => n39231, ZN => n36542);
   U32021 : AOI221_X1 port map( B1 => n39255, B2 => n29709, C1 => n39249, C2 =>
                           n29773, A => n36523, ZN => n36520);
   U32022 : OAI222_X1 port map( A1 => n31837, A2 => n39243, B1 => n31897, B2 =>
                           n39237, C1 => n31777, C2 => n39231, ZN => n36523);
   U32023 : AOI221_X1 port map( B1 => n39255, B2 => n29708, C1 => n39249, C2 =>
                           n29772, A => n36504, ZN => n36501);
   U32024 : OAI222_X1 port map( A1 => n31836, A2 => n39243, B1 => n31896, B2 =>
                           n39237, C1 => n31776, C2 => n39231, ZN => n36504);
   U32025 : AOI221_X1 port map( B1 => n39255, B2 => n29707, C1 => n39249, C2 =>
                           n29771, A => n36485, ZN => n36482);
   U32026 : OAI222_X1 port map( A1 => n31835, A2 => n39243, B1 => n31895, B2 =>
                           n39237, C1 => n31775, C2 => n39231, ZN => n36485);
   U32027 : AOI221_X1 port map( B1 => n39255, B2 => n29706, C1 => n39249, C2 =>
                           n29770, A => n36466, ZN => n36463);
   U32028 : OAI222_X1 port map( A1 => n31834, A2 => n39243, B1 => n31894, B2 =>
                           n39237, C1 => n31774, C2 => n39231, ZN => n36466);
   U32029 : AOI221_X1 port map( B1 => n39255, B2 => n29705, C1 => n39249, C2 =>
                           n29769, A => n36447, ZN => n36444);
   U32030 : OAI222_X1 port map( A1 => n31833, A2 => n39243, B1 => n31893, B2 =>
                           n39237, C1 => n31773, C2 => n39231, ZN => n36447);
   U32031 : AOI221_X1 port map( B1 => n39255, B2 => n29704, C1 => n39249, C2 =>
                           n29768, A => n36428, ZN => n36425);
   U32032 : OAI222_X1 port map( A1 => n31832, A2 => n39243, B1 => n31892, B2 =>
                           n39237, C1 => n31772, C2 => n39231, ZN => n36428);
   U32033 : AOI221_X1 port map( B1 => n39255, B2 => n29703, C1 => n39249, C2 =>
                           n29767, A => n36409, ZN => n36406);
   U32034 : OAI222_X1 port map( A1 => n31831, A2 => n39243, B1 => n31891, B2 =>
                           n39237, C1 => n31771, C2 => n39231, ZN => n36409);
   U32035 : AOI221_X1 port map( B1 => n39255, B2 => n29702, C1 => n39249, C2 =>
                           n29766, A => n36390, ZN => n36387);
   U32036 : OAI222_X1 port map( A1 => n31830, A2 => n39243, B1 => n31890, B2 =>
                           n39237, C1 => n31770, C2 => n39231, ZN => n36390);
   U32037 : AOI221_X1 port map( B1 => n39255, B2 => n29701, C1 => n39249, C2 =>
                           n29765, A => n36371, ZN => n36368);
   U32038 : OAI222_X1 port map( A1 => n31829, A2 => n39243, B1 => n31889, B2 =>
                           n39237, C1 => n31769, C2 => n39231, ZN => n36371);
   U32039 : AOI221_X1 port map( B1 => n39255, B2 => n29700, C1 => n39249, C2 =>
                           n29764, A => n36352, ZN => n36349);
   U32040 : OAI222_X1 port map( A1 => n31828, A2 => n39243, B1 => n31888, B2 =>
                           n39237, C1 => n31768, C2 => n39231, ZN => n36352);
   U32041 : AOI221_X1 port map( B1 => n39255, B2 => n29699, C1 => n39249, C2 =>
                           n29763, A => n36333, ZN => n36330);
   U32042 : OAI222_X1 port map( A1 => n31827, A2 => n39243, B1 => n31887, B2 =>
                           n39237, C1 => n31767, C2 => n39231, ZN => n36333);
   U32043 : AOI221_X1 port map( B1 => n39256, B2 => n29698, C1 => n39250, C2 =>
                           n29762, A => n36314, ZN => n36311);
   U32044 : OAI222_X1 port map( A1 => n31826, A2 => n39244, B1 => n31886, B2 =>
                           n39238, C1 => n31766, C2 => n39232, ZN => n36314);
   U32045 : AOI221_X1 port map( B1 => n39256, B2 => n29697, C1 => n39250, C2 =>
                           n29761, A => n36295, ZN => n36292);
   U32046 : OAI222_X1 port map( A1 => n31825, A2 => n39244, B1 => n31885, B2 =>
                           n39238, C1 => n31765, C2 => n39232, ZN => n36295);
   U32047 : AOI221_X1 port map( B1 => n39256, B2 => n29696, C1 => n39250, C2 =>
                           n29760, A => n36276, ZN => n36273);
   U32048 : OAI222_X1 port map( A1 => n31824, A2 => n39244, B1 => n31884, B2 =>
                           n39238, C1 => n31764, C2 => n39232, ZN => n36276);
   U32049 : AOI221_X1 port map( B1 => n39256, B2 => n29695, C1 => n39250, C2 =>
                           n29759, A => n36257, ZN => n36254);
   U32050 : OAI222_X1 port map( A1 => n31823, A2 => n39244, B1 => n31883, B2 =>
                           n39238, C1 => n31763, C2 => n39232, ZN => n36257);
   U32051 : AOI221_X1 port map( B1 => n39256, B2 => n29694, C1 => n39250, C2 =>
                           n29758, A => n36238, ZN => n36235);
   U32052 : OAI222_X1 port map( A1 => n31822, A2 => n39244, B1 => n31882, B2 =>
                           n39238, C1 => n31762, C2 => n39232, ZN => n36238);
   U32053 : AOI221_X1 port map( B1 => n39256, B2 => n29693, C1 => n39250, C2 =>
                           n29757, A => n36219, ZN => n36216);
   U32054 : OAI222_X1 port map( A1 => n31821, A2 => n39244, B1 => n31881, B2 =>
                           n39238, C1 => n31761, C2 => n39232, ZN => n36219);
   U32055 : AOI221_X1 port map( B1 => n39252, B2 => n29745, C1 => n39246, C2 =>
                           n29809, A => n37207, ZN => n37204);
   U32056 : OAI222_X1 port map( A1 => n32268, A2 => n39240, B1 => n32272, B2 =>
                           n39234, C1 => n32276, C2 => n39228, ZN => n37207);
   U32057 : AOI221_X1 port map( B1 => n39252, B2 => n29744, C1 => n39246, C2 =>
                           n29808, A => n37188, ZN => n37185);
   U32058 : OAI222_X1 port map( A1 => n32267, A2 => n39240, B1 => n32271, B2 =>
                           n39234, C1 => n32275, C2 => n39228, ZN => n37188);
   U32059 : AOI221_X1 port map( B1 => n39252, B2 => n29743, C1 => n39246, C2 =>
                           n29807, A => n37169, ZN => n37166);
   U32060 : OAI222_X1 port map( A1 => n32266, A2 => n39240, B1 => n32270, B2 =>
                           n39234, C1 => n32274, C2 => n39228, ZN => n37169);
   U32061 : AOI221_X1 port map( B1 => n39252, B2 => n29742, C1 => n39246, C2 =>
                           n29806, A => n37150, ZN => n37147);
   U32062 : OAI222_X1 port map( A1 => n31870, A2 => n39240, B1 => n31930, B2 =>
                           n39234, C1 => n31810, C2 => n39228, ZN => n37150);
   U32063 : AOI221_X1 port map( B1 => n39252, B2 => n29741, C1 => n39246, C2 =>
                           n29805, A => n37131, ZN => n37128);
   U32064 : OAI222_X1 port map( A1 => n31869, A2 => n39240, B1 => n31929, B2 =>
                           n39234, C1 => n31809, C2 => n39228, ZN => n37131);
   U32065 : AOI221_X1 port map( B1 => n39257, B2 => n29686, C1 => n39251, C2 =>
                           n29750, A => n36086, ZN => n36083);
   U32066 : OAI222_X1 port map( A1 => n31814, A2 => n39245, B1 => n31874, B2 =>
                           n39239, C1 => n31754, C2 => n39233, ZN => n36086);
   U32067 : AOI221_X1 port map( B1 => n39257, B2 => n29685, C1 => n39251, C2 =>
                           n29749, A => n36067, ZN => n36064);
   U32068 : OAI222_X1 port map( A1 => n31813, A2 => n39245, B1 => n31873, B2 =>
                           n39239, C1 => n31753, C2 => n39233, ZN => n36067);
   U32069 : AOI221_X1 port map( B1 => n39257, B2 => n29684, C1 => n39251, C2 =>
                           n29748, A => n36048, ZN => n36045);
   U32070 : OAI222_X1 port map( A1 => n31812, A2 => n39245, B1 => n31872, B2 =>
                           n39239, C1 => n31752, C2 => n39233, ZN => n36048);
   U32071 : AOI221_X1 port map( B1 => n39257, B2 => n29683, C1 => n39251, C2 =>
                           n29747, A => n35996, ZN => n35986);
   U32072 : OAI222_X1 port map( A1 => n31811, A2 => n39245, B1 => n31871, B2 =>
                           n39239, C1 => n31751, C2 => n39233, ZN => n35996);
   U32073 : AOI221_X1 port map( B1 => n39252, B2 => n29746, C1 => n39246, C2 =>
                           n29810, A => n37232, ZN => n37223);
   U32074 : OAI222_X1 port map( A1 => n32269, A2 => n39240, B1 => n32273, B2 =>
                           n39234, C1 => n32277, C2 => n39228, ZN => n37232);
   U32075 : AOI221_X1 port map( B1 => n39252, B2 => n29740, C1 => n39246, C2 =>
                           n29804, A => n37112, ZN => n37109);
   U32076 : OAI222_X1 port map( A1 => n31868, A2 => n39240, B1 => n31928, B2 =>
                           n39234, C1 => n31808, C2 => n39228, ZN => n37112);
   U32077 : AOI221_X1 port map( B1 => n39252, B2 => n29739, C1 => n39246, C2 =>
                           n29803, A => n37093, ZN => n37090);
   U32078 : OAI222_X1 port map( A1 => n31867, A2 => n39240, B1 => n31927, B2 =>
                           n39234, C1 => n31807, C2 => n39228, ZN => n37093);
   U32079 : AOI221_X1 port map( B1 => n39252, B2 => n29738, C1 => n39246, C2 =>
                           n29802, A => n37074, ZN => n37071);
   U32080 : OAI222_X1 port map( A1 => n31866, A2 => n39240, B1 => n31926, B2 =>
                           n39234, C1 => n31806, C2 => n39228, ZN => n37074);
   U32081 : AOI221_X1 port map( B1 => n39252, B2 => n29737, C1 => n39246, C2 =>
                           n29801, A => n37055, ZN => n37052);
   U32082 : OAI222_X1 port map( A1 => n31865, A2 => n39240, B1 => n31925, B2 =>
                           n39234, C1 => n31805, C2 => n39228, ZN => n37055);
   U32083 : AOI221_X1 port map( B1 => n39252, B2 => n29736, C1 => n39246, C2 =>
                           n29800, A => n37036, ZN => n37033);
   U32084 : OAI222_X1 port map( A1 => n31864, A2 => n39240, B1 => n31924, B2 =>
                           n39234, C1 => n31804, C2 => n39228, ZN => n37036);
   U32085 : AOI221_X1 port map( B1 => n39256, B2 => n29692, C1 => n39250, C2 =>
                           n29756, A => n36200, ZN => n36197);
   U32086 : OAI222_X1 port map( A1 => n31820, A2 => n39244, B1 => n31880, B2 =>
                           n39238, C1 => n31760, C2 => n39232, ZN => n36200);
   U32087 : AOI221_X1 port map( B1 => n39256, B2 => n29691, C1 => n39250, C2 =>
                           n29755, A => n36181, ZN => n36178);
   U32088 : OAI222_X1 port map( A1 => n31819, A2 => n39244, B1 => n31879, B2 =>
                           n39238, C1 => n31759, C2 => n39232, ZN => n36181);
   U32089 : AOI221_X1 port map( B1 => n39256, B2 => n29690, C1 => n39250, C2 =>
                           n29754, A => n36162, ZN => n36159);
   U32090 : OAI222_X1 port map( A1 => n31818, A2 => n39244, B1 => n31878, B2 =>
                           n39238, C1 => n31758, C2 => n39232, ZN => n36162);
   U32091 : AOI221_X1 port map( B1 => n39256, B2 => n29689, C1 => n39250, C2 =>
                           n29753, A => n36143, ZN => n36140);
   U32092 : OAI222_X1 port map( A1 => n31817, A2 => n39244, B1 => n31877, B2 =>
                           n39238, C1 => n31757, C2 => n39232, ZN => n36143);
   U32093 : AOI221_X1 port map( B1 => n39256, B2 => n29688, C1 => n39250, C2 =>
                           n29752, A => n36124, ZN => n36121);
   U32094 : OAI222_X1 port map( A1 => n31816, A2 => n39244, B1 => n31876, B2 =>
                           n39238, C1 => n31756, C2 => n39232, ZN => n36124);
   U32095 : AOI221_X1 port map( B1 => n39256, B2 => n29687, C1 => n39250, C2 =>
                           n29751, A => n36105, ZN => n36102);
   U32096 : OAI222_X1 port map( A1 => n31815, A2 => n39244, B1 => n31875, B2 =>
                           n39238, C1 => n31755, C2 => n39232, ZN => n36105);
   U32097 : AOI221_X1 port map( B1 => n39759, B2 => n29746, C1 => n39753, C2 =>
                           n29810, A => n33441, ZN => n33431);
   U32098 : OAI222_X1 port map( A1 => n32269, A2 => n39747, B1 => n32273, B2 =>
                           n39741, C1 => n32277, C2 => n39735, ZN => n33441);
   U32099 : AOI221_X1 port map( B1 => n39507, B2 => n29746, C1 => n39501, C2 =>
                           n29810, A => n34715, ZN => n34705);
   U32100 : OAI222_X1 port map( A1 => n32269, A2 => n39495, B1 => n32273, B2 =>
                           n39489, C1 => n32277, C2 => n39483, ZN => n34715);
   U32101 : AOI221_X1 port map( B1 => n39759, B2 => n29745, C1 => n39753, C2 =>
                           n29809, A => n33493, ZN => n33490);
   U32102 : OAI222_X1 port map( A1 => n32268, A2 => n39747, B1 => n32272, B2 =>
                           n39741, C1 => n32276, C2 => n39735, ZN => n33493);
   U32103 : AOI221_X1 port map( B1 => n39507, B2 => n29745, C1 => n39501, C2 =>
                           n29809, A => n34767, ZN => n34764);
   U32104 : OAI222_X1 port map( A1 => n32268, A2 => n39495, B1 => n32272, B2 =>
                           n39489, C1 => n32276, C2 => n39483, ZN => n34767);
   U32105 : AOI221_X1 port map( B1 => n39759, B2 => n29744, C1 => n39753, C2 =>
                           n29808, A => n33512, ZN => n33509);
   U32106 : OAI222_X1 port map( A1 => n32267, A2 => n39747, B1 => n32271, B2 =>
                           n39741, C1 => n32275, C2 => n39735, ZN => n33512);
   U32107 : AOI221_X1 port map( B1 => n39507, B2 => n29744, C1 => n39501, C2 =>
                           n29808, A => n34786, ZN => n34783);
   U32108 : OAI222_X1 port map( A1 => n32267, A2 => n39495, B1 => n32271, B2 =>
                           n39489, C1 => n32275, C2 => n39483, ZN => n34786);
   U32109 : AOI221_X1 port map( B1 => n39759, B2 => n29743, C1 => n39753, C2 =>
                           n29807, A => n33531, ZN => n33528);
   U32110 : OAI222_X1 port map( A1 => n32266, A2 => n39747, B1 => n32270, B2 =>
                           n39741, C1 => n32274, C2 => n39735, ZN => n33531);
   U32111 : AOI221_X1 port map( B1 => n39507, B2 => n29743, C1 => n39501, C2 =>
                           n29807, A => n34805, ZN => n34802);
   U32112 : OAI222_X1 port map( A1 => n32266, A2 => n39495, B1 => n32270, B2 =>
                           n39489, C1 => n32274, C2 => n39483, ZN => n34805);
   U32113 : AOI221_X1 port map( B1 => n39758, B2 => n29742, C1 => n39752, C2 =>
                           n29806, A => n33550, ZN => n33547);
   U32114 : OAI222_X1 port map( A1 => n31870, A2 => n39746, B1 => n31930, B2 =>
                           n39740, C1 => n31810, C2 => n39734, ZN => n33550);
   U32115 : AOI221_X1 port map( B1 => n39506, B2 => n29742, C1 => n39500, C2 =>
                           n29806, A => n34824, ZN => n34821);
   U32116 : OAI222_X1 port map( A1 => n31870, A2 => n39494, B1 => n31930, B2 =>
                           n39488, C1 => n31810, C2 => n39482, ZN => n34824);
   U32117 : AOI221_X1 port map( B1 => n39758, B2 => n29741, C1 => n39752, C2 =>
                           n29805, A => n33569, ZN => n33566);
   U32118 : OAI222_X1 port map( A1 => n31869, A2 => n39746, B1 => n31929, B2 =>
                           n39740, C1 => n31809, C2 => n39734, ZN => n33569);
   U32119 : AOI221_X1 port map( B1 => n39506, B2 => n29741, C1 => n39500, C2 =>
                           n29805, A => n34843, ZN => n34840);
   U32120 : OAI222_X1 port map( A1 => n31869, A2 => n39494, B1 => n31929, B2 =>
                           n39488, C1 => n31809, C2 => n39482, ZN => n34843);
   U32121 : AOI221_X1 port map( B1 => n39758, B2 => n29740, C1 => n39752, C2 =>
                           n29804, A => n33588, ZN => n33585);
   U32122 : OAI222_X1 port map( A1 => n31868, A2 => n39746, B1 => n31928, B2 =>
                           n39740, C1 => n31808, C2 => n39734, ZN => n33588);
   U32123 : AOI221_X1 port map( B1 => n39506, B2 => n29740, C1 => n39500, C2 =>
                           n29804, A => n34862, ZN => n34859);
   U32124 : OAI222_X1 port map( A1 => n31868, A2 => n39494, B1 => n31928, B2 =>
                           n39488, C1 => n31808, C2 => n39482, ZN => n34862);
   U32125 : AOI221_X1 port map( B1 => n39758, B2 => n29739, C1 => n39752, C2 =>
                           n29803, A => n33607, ZN => n33604);
   U32126 : OAI222_X1 port map( A1 => n31867, A2 => n39746, B1 => n31927, B2 =>
                           n39740, C1 => n31807, C2 => n39734, ZN => n33607);
   U32127 : AOI221_X1 port map( B1 => n39506, B2 => n29739, C1 => n39500, C2 =>
                           n29803, A => n34881, ZN => n34878);
   U32128 : OAI222_X1 port map( A1 => n31867, A2 => n39494, B1 => n31927, B2 =>
                           n39488, C1 => n31807, C2 => n39482, ZN => n34881);
   U32129 : AOI221_X1 port map( B1 => n39758, B2 => n29738, C1 => n39752, C2 =>
                           n29802, A => n33626, ZN => n33623);
   U32130 : OAI222_X1 port map( A1 => n31866, A2 => n39746, B1 => n31926, B2 =>
                           n39740, C1 => n31806, C2 => n39734, ZN => n33626);
   U32131 : AOI221_X1 port map( B1 => n39506, B2 => n29738, C1 => n39500, C2 =>
                           n29802, A => n34900, ZN => n34897);
   U32132 : OAI222_X1 port map( A1 => n31866, A2 => n39494, B1 => n31926, B2 =>
                           n39488, C1 => n31806, C2 => n39482, ZN => n34900);
   U32133 : AOI221_X1 port map( B1 => n39758, B2 => n29737, C1 => n39752, C2 =>
                           n29801, A => n33645, ZN => n33642);
   U32134 : OAI222_X1 port map( A1 => n31865, A2 => n39746, B1 => n31925, B2 =>
                           n39740, C1 => n31805, C2 => n39734, ZN => n33645);
   U32135 : AOI221_X1 port map( B1 => n39506, B2 => n29737, C1 => n39500, C2 =>
                           n29801, A => n34919, ZN => n34916);
   U32136 : OAI222_X1 port map( A1 => n31865, A2 => n39494, B1 => n31925, B2 =>
                           n39488, C1 => n31805, C2 => n39482, ZN => n34919);
   U32137 : AOI221_X1 port map( B1 => n39758, B2 => n29736, C1 => n39752, C2 =>
                           n29800, A => n33664, ZN => n33661);
   U32138 : OAI222_X1 port map( A1 => n31864, A2 => n39746, B1 => n31924, B2 =>
                           n39740, C1 => n31804, C2 => n39734, ZN => n33664);
   U32139 : AOI221_X1 port map( B1 => n39506, B2 => n29736, C1 => n39500, C2 =>
                           n29800, A => n34938, ZN => n34935);
   U32140 : OAI222_X1 port map( A1 => n31864, A2 => n39494, B1 => n31924, B2 =>
                           n39488, C1 => n31804, C2 => n39482, ZN => n34938);
   U32141 : AOI221_X1 port map( B1 => n39758, B2 => n29735, C1 => n39752, C2 =>
                           n29799, A => n33683, ZN => n33680);
   U32142 : OAI222_X1 port map( A1 => n31863, A2 => n39746, B1 => n31923, B2 =>
                           n39740, C1 => n31803, C2 => n39734, ZN => n33683);
   U32143 : AOI221_X1 port map( B1 => n39506, B2 => n29735, C1 => n39500, C2 =>
                           n29799, A => n34957, ZN => n34954);
   U32144 : OAI222_X1 port map( A1 => n31863, A2 => n39494, B1 => n31923, B2 =>
                           n39488, C1 => n31803, C2 => n39482, ZN => n34957);
   U32145 : AOI221_X1 port map( B1 => n39758, B2 => n29734, C1 => n39752, C2 =>
                           n29798, A => n33702, ZN => n33699);
   U32146 : OAI222_X1 port map( A1 => n31862, A2 => n39746, B1 => n31922, B2 =>
                           n39740, C1 => n31802, C2 => n39734, ZN => n33702);
   U32147 : AOI221_X1 port map( B1 => n39506, B2 => n29734, C1 => n39500, C2 =>
                           n29798, A => n34976, ZN => n34973);
   U32148 : OAI222_X1 port map( A1 => n31862, A2 => n39494, B1 => n31922, B2 =>
                           n39488, C1 => n31802, C2 => n39482, ZN => n34976);
   U32149 : AOI221_X1 port map( B1 => n39758, B2 => n29733, C1 => n39752, C2 =>
                           n29797, A => n33721, ZN => n33718);
   U32150 : OAI222_X1 port map( A1 => n31861, A2 => n39746, B1 => n31921, B2 =>
                           n39740, C1 => n31801, C2 => n39734, ZN => n33721);
   U32151 : AOI221_X1 port map( B1 => n39506, B2 => n29733, C1 => n39500, C2 =>
                           n29797, A => n34995, ZN => n34992);
   U32152 : OAI222_X1 port map( A1 => n31861, A2 => n39494, B1 => n31921, B2 =>
                           n39488, C1 => n31801, C2 => n39482, ZN => n34995);
   U32153 : AOI221_X1 port map( B1 => n39758, B2 => n29732, C1 => n39752, C2 =>
                           n29796, A => n33740, ZN => n33737);
   U32154 : OAI222_X1 port map( A1 => n31860, A2 => n39746, B1 => n31920, B2 =>
                           n39740, C1 => n31800, C2 => n39734, ZN => n33740);
   U32155 : AOI221_X1 port map( B1 => n39506, B2 => n29732, C1 => n39500, C2 =>
                           n29796, A => n35014, ZN => n35011);
   U32156 : OAI222_X1 port map( A1 => n31860, A2 => n39494, B1 => n31920, B2 =>
                           n39488, C1 => n31800, C2 => n39482, ZN => n35014);
   U32157 : AOI221_X1 port map( B1 => n39758, B2 => n29731, C1 => n39752, C2 =>
                           n29795, A => n33759, ZN => n33756);
   U32158 : OAI222_X1 port map( A1 => n31859, A2 => n39746, B1 => n31919, B2 =>
                           n39740, C1 => n31799, C2 => n39734, ZN => n33759);
   U32159 : AOI221_X1 port map( B1 => n39506, B2 => n29731, C1 => n39500, C2 =>
                           n29795, A => n35033, ZN => n35030);
   U32160 : OAI222_X1 port map( A1 => n31859, A2 => n39494, B1 => n31919, B2 =>
                           n39488, C1 => n31799, C2 => n39482, ZN => n35033);
   U32161 : AOI221_X1 port map( B1 => n39757, B2 => n29730, C1 => n39751, C2 =>
                           n29794, A => n33778, ZN => n33775);
   U32162 : OAI222_X1 port map( A1 => n31858, A2 => n39745, B1 => n31918, B2 =>
                           n39739, C1 => n31798, C2 => n39733, ZN => n33778);
   U32163 : AOI221_X1 port map( B1 => n39505, B2 => n29730, C1 => n39499, C2 =>
                           n29794, A => n35052, ZN => n35049);
   U32164 : OAI222_X1 port map( A1 => n31858, A2 => n39493, B1 => n31918, B2 =>
                           n39487, C1 => n31798, C2 => n39481, ZN => n35052);
   U32165 : AOI221_X1 port map( B1 => n39757, B2 => n29729, C1 => n39751, C2 =>
                           n29793, A => n33797, ZN => n33794);
   U32166 : OAI222_X1 port map( A1 => n31857, A2 => n39745, B1 => n31917, B2 =>
                           n39739, C1 => n31797, C2 => n39733, ZN => n33797);
   U32167 : AOI221_X1 port map( B1 => n39505, B2 => n29729, C1 => n39499, C2 =>
                           n29793, A => n35071, ZN => n35068);
   U32168 : OAI222_X1 port map( A1 => n31857, A2 => n39493, B1 => n31917, B2 =>
                           n39487, C1 => n31797, C2 => n39481, ZN => n35071);
   U32169 : AOI221_X1 port map( B1 => n39757, B2 => n29728, C1 => n39751, C2 =>
                           n29792, A => n33816, ZN => n33813);
   U32170 : OAI222_X1 port map( A1 => n31856, A2 => n39745, B1 => n31916, B2 =>
                           n39739, C1 => n31796, C2 => n39733, ZN => n33816);
   U32171 : AOI221_X1 port map( B1 => n39505, B2 => n29728, C1 => n39499, C2 =>
                           n29792, A => n35090, ZN => n35087);
   U32172 : OAI222_X1 port map( A1 => n31856, A2 => n39493, B1 => n31916, B2 =>
                           n39487, C1 => n31796, C2 => n39481, ZN => n35090);
   U32173 : AOI221_X1 port map( B1 => n39757, B2 => n29727, C1 => n39751, C2 =>
                           n29791, A => n33835, ZN => n33832);
   U32174 : OAI222_X1 port map( A1 => n31855, A2 => n39745, B1 => n31915, B2 =>
                           n39739, C1 => n31795, C2 => n39733, ZN => n33835);
   U32175 : AOI221_X1 port map( B1 => n39505, B2 => n29727, C1 => n39499, C2 =>
                           n29791, A => n35109, ZN => n35106);
   U32176 : OAI222_X1 port map( A1 => n31855, A2 => n39493, B1 => n31915, B2 =>
                           n39487, C1 => n31795, C2 => n39481, ZN => n35109);
   U32177 : AOI221_X1 port map( B1 => n39757, B2 => n29726, C1 => n39751, C2 =>
                           n29790, A => n33854, ZN => n33851);
   U32178 : OAI222_X1 port map( A1 => n31854, A2 => n39745, B1 => n31914, B2 =>
                           n39739, C1 => n31794, C2 => n39733, ZN => n33854);
   U32179 : AOI221_X1 port map( B1 => n39505, B2 => n29726, C1 => n39499, C2 =>
                           n29790, A => n35128, ZN => n35125);
   U32180 : OAI222_X1 port map( A1 => n31854, A2 => n39493, B1 => n31914, B2 =>
                           n39487, C1 => n31794, C2 => n39481, ZN => n35128);
   U32181 : AOI221_X1 port map( B1 => n39757, B2 => n29725, C1 => n39751, C2 =>
                           n29789, A => n33873, ZN => n33870);
   U32182 : OAI222_X1 port map( A1 => n31853, A2 => n39745, B1 => n31913, B2 =>
                           n39739, C1 => n31793, C2 => n39733, ZN => n33873);
   U32183 : AOI221_X1 port map( B1 => n39505, B2 => n29725, C1 => n39499, C2 =>
                           n29789, A => n35147, ZN => n35144);
   U32184 : OAI222_X1 port map( A1 => n31853, A2 => n39493, B1 => n31913, B2 =>
                           n39487, C1 => n31793, C2 => n39481, ZN => n35147);
   U32185 : AOI221_X1 port map( B1 => n39757, B2 => n29724, C1 => n39751, C2 =>
                           n29788, A => n33892, ZN => n33889);
   U32186 : OAI222_X1 port map( A1 => n31852, A2 => n39745, B1 => n31912, B2 =>
                           n39739, C1 => n31792, C2 => n39733, ZN => n33892);
   U32187 : AOI221_X1 port map( B1 => n39505, B2 => n29724, C1 => n39499, C2 =>
                           n29788, A => n35166, ZN => n35163);
   U32188 : OAI222_X1 port map( A1 => n31852, A2 => n39493, B1 => n31912, B2 =>
                           n39487, C1 => n31792, C2 => n39481, ZN => n35166);
   U32189 : AOI221_X1 port map( B1 => n39757, B2 => n29723, C1 => n39751, C2 =>
                           n29787, A => n33911, ZN => n33908);
   U32190 : OAI222_X1 port map( A1 => n31851, A2 => n39745, B1 => n31911, B2 =>
                           n39739, C1 => n31791, C2 => n39733, ZN => n33911);
   U32191 : AOI221_X1 port map( B1 => n39505, B2 => n29723, C1 => n39499, C2 =>
                           n29787, A => n35185, ZN => n35182);
   U32192 : OAI222_X1 port map( A1 => n31851, A2 => n39493, B1 => n31911, B2 =>
                           n39487, C1 => n31791, C2 => n39481, ZN => n35185);
   U32193 : AOI221_X1 port map( B1 => n39757, B2 => n29722, C1 => n39751, C2 =>
                           n29786, A => n33930, ZN => n33927);
   U32194 : OAI222_X1 port map( A1 => n31850, A2 => n39745, B1 => n31910, B2 =>
                           n39739, C1 => n31790, C2 => n39733, ZN => n33930);
   U32195 : AOI221_X1 port map( B1 => n39505, B2 => n29722, C1 => n39499, C2 =>
                           n29786, A => n35204, ZN => n35201);
   U32196 : OAI222_X1 port map( A1 => n31850, A2 => n39493, B1 => n31910, B2 =>
                           n39487, C1 => n31790, C2 => n39481, ZN => n35204);
   U32197 : AOI221_X1 port map( B1 => n39757, B2 => n29721, C1 => n39751, C2 =>
                           n29785, A => n33949, ZN => n33946);
   U32198 : OAI222_X1 port map( A1 => n31849, A2 => n39745, B1 => n31909, B2 =>
                           n39739, C1 => n31789, C2 => n39733, ZN => n33949);
   U32199 : AOI221_X1 port map( B1 => n39505, B2 => n29721, C1 => n39499, C2 =>
                           n29785, A => n35223, ZN => n35220);
   U32200 : OAI222_X1 port map( A1 => n31849, A2 => n39493, B1 => n31909, B2 =>
                           n39487, C1 => n31789, C2 => n39481, ZN => n35223);
   U32201 : AOI221_X1 port map( B1 => n39757, B2 => n29720, C1 => n39751, C2 =>
                           n29784, A => n33968, ZN => n33965);
   U32202 : OAI222_X1 port map( A1 => n31848, A2 => n39745, B1 => n31908, B2 =>
                           n39739, C1 => n31788, C2 => n39733, ZN => n33968);
   U32203 : AOI221_X1 port map( B1 => n39505, B2 => n29720, C1 => n39499, C2 =>
                           n29784, A => n35242, ZN => n35239);
   U32204 : OAI222_X1 port map( A1 => n31848, A2 => n39493, B1 => n31908, B2 =>
                           n39487, C1 => n31788, C2 => n39481, ZN => n35242);
   U32205 : AOI221_X1 port map( B1 => n39757, B2 => n29719, C1 => n39751, C2 =>
                           n29783, A => n33987, ZN => n33984);
   U32206 : OAI222_X1 port map( A1 => n31847, A2 => n39745, B1 => n31907, B2 =>
                           n39739, C1 => n31787, C2 => n39733, ZN => n33987);
   U32207 : AOI221_X1 port map( B1 => n39505, B2 => n29719, C1 => n39499, C2 =>
                           n29783, A => n35261, ZN => n35258);
   U32208 : OAI222_X1 port map( A1 => n31847, A2 => n39493, B1 => n31907, B2 =>
                           n39487, C1 => n31787, C2 => n39481, ZN => n35261);
   U32209 : AOI221_X1 port map( B1 => n39756, B2 => n29718, C1 => n39750, C2 =>
                           n29782, A => n34006, ZN => n34003);
   U32210 : OAI222_X1 port map( A1 => n31846, A2 => n39744, B1 => n31906, B2 =>
                           n39738, C1 => n31786, C2 => n39732, ZN => n34006);
   U32211 : AOI221_X1 port map( B1 => n39504, B2 => n29718, C1 => n39498, C2 =>
                           n29782, A => n35280, ZN => n35277);
   U32212 : OAI222_X1 port map( A1 => n31846, A2 => n39492, B1 => n31906, B2 =>
                           n39486, C1 => n31786, C2 => n39480, ZN => n35280);
   U32213 : AOI221_X1 port map( B1 => n39756, B2 => n29717, C1 => n39750, C2 =>
                           n29781, A => n34025, ZN => n34022);
   U32214 : OAI222_X1 port map( A1 => n31845, A2 => n39744, B1 => n31905, B2 =>
                           n39738, C1 => n31785, C2 => n39732, ZN => n34025);
   U32215 : AOI221_X1 port map( B1 => n39504, B2 => n29717, C1 => n39498, C2 =>
                           n29781, A => n35299, ZN => n35296);
   U32216 : OAI222_X1 port map( A1 => n31845, A2 => n39492, B1 => n31905, B2 =>
                           n39486, C1 => n31785, C2 => n39480, ZN => n35299);
   U32217 : AOI221_X1 port map( B1 => n39756, B2 => n29716, C1 => n39750, C2 =>
                           n29780, A => n34044, ZN => n34041);
   U32218 : OAI222_X1 port map( A1 => n31844, A2 => n39744, B1 => n31904, B2 =>
                           n39738, C1 => n31784, C2 => n39732, ZN => n34044);
   U32219 : AOI221_X1 port map( B1 => n39504, B2 => n29716, C1 => n39498, C2 =>
                           n29780, A => n35318, ZN => n35315);
   U32220 : OAI222_X1 port map( A1 => n31844, A2 => n39492, B1 => n31904, B2 =>
                           n39486, C1 => n31784, C2 => n39480, ZN => n35318);
   U32221 : AOI221_X1 port map( B1 => n39756, B2 => n29715, C1 => n39750, C2 =>
                           n29779, A => n34063, ZN => n34060);
   U32222 : OAI222_X1 port map( A1 => n31843, A2 => n39744, B1 => n31903, B2 =>
                           n39738, C1 => n31783, C2 => n39732, ZN => n34063);
   U32223 : AOI221_X1 port map( B1 => n39504, B2 => n29715, C1 => n39498, C2 =>
                           n29779, A => n35337, ZN => n35334);
   U32224 : OAI222_X1 port map( A1 => n31843, A2 => n39492, B1 => n31903, B2 =>
                           n39486, C1 => n31783, C2 => n39480, ZN => n35337);
   U32225 : AOI221_X1 port map( B1 => n39756, B2 => n29714, C1 => n39750, C2 =>
                           n29778, A => n34082, ZN => n34079);
   U32226 : OAI222_X1 port map( A1 => n31842, A2 => n39744, B1 => n31902, B2 =>
                           n39738, C1 => n31782, C2 => n39732, ZN => n34082);
   U32227 : AOI221_X1 port map( B1 => n39504, B2 => n29714, C1 => n39498, C2 =>
                           n29778, A => n35356, ZN => n35353);
   U32228 : OAI222_X1 port map( A1 => n31842, A2 => n39492, B1 => n31902, B2 =>
                           n39486, C1 => n31782, C2 => n39480, ZN => n35356);
   U32229 : AOI221_X1 port map( B1 => n39756, B2 => n29713, C1 => n39750, C2 =>
                           n29777, A => n34101, ZN => n34098);
   U32230 : OAI222_X1 port map( A1 => n31841, A2 => n39744, B1 => n31901, B2 =>
                           n39738, C1 => n31781, C2 => n39732, ZN => n34101);
   U32231 : AOI221_X1 port map( B1 => n39504, B2 => n29713, C1 => n39498, C2 =>
                           n29777, A => n35375, ZN => n35372);
   U32232 : OAI222_X1 port map( A1 => n31841, A2 => n39492, B1 => n31901, B2 =>
                           n39486, C1 => n31781, C2 => n39480, ZN => n35375);
   U32233 : AOI221_X1 port map( B1 => n39756, B2 => n29712, C1 => n39750, C2 =>
                           n29776, A => n34120, ZN => n34117);
   U32234 : OAI222_X1 port map( A1 => n31840, A2 => n39744, B1 => n31900, B2 =>
                           n39738, C1 => n31780, C2 => n39732, ZN => n34120);
   U32235 : AOI221_X1 port map( B1 => n39504, B2 => n29712, C1 => n39498, C2 =>
                           n29776, A => n35394, ZN => n35391);
   U32236 : OAI222_X1 port map( A1 => n31840, A2 => n39492, B1 => n31900, B2 =>
                           n39486, C1 => n31780, C2 => n39480, ZN => n35394);
   U32237 : AOI221_X1 port map( B1 => n39756, B2 => n29711, C1 => n39750, C2 =>
                           n29775, A => n34139, ZN => n34136);
   U32238 : OAI222_X1 port map( A1 => n31839, A2 => n39744, B1 => n31899, B2 =>
                           n39738, C1 => n31779, C2 => n39732, ZN => n34139);
   U32239 : AOI221_X1 port map( B1 => n39504, B2 => n29711, C1 => n39498, C2 =>
                           n29775, A => n35413, ZN => n35410);
   U32240 : OAI222_X1 port map( A1 => n31839, A2 => n39492, B1 => n31899, B2 =>
                           n39486, C1 => n31779, C2 => n39480, ZN => n35413);
   U32241 : AOI221_X1 port map( B1 => n39756, B2 => n29710, C1 => n39750, C2 =>
                           n29774, A => n34158, ZN => n34155);
   U32242 : OAI222_X1 port map( A1 => n31838, A2 => n39744, B1 => n31898, B2 =>
                           n39738, C1 => n31778, C2 => n39732, ZN => n34158);
   U32243 : AOI221_X1 port map( B1 => n39504, B2 => n29710, C1 => n39498, C2 =>
                           n29774, A => n35432, ZN => n35429);
   U32244 : OAI222_X1 port map( A1 => n31838, A2 => n39492, B1 => n31898, B2 =>
                           n39486, C1 => n31778, C2 => n39480, ZN => n35432);
   U32245 : AOI221_X1 port map( B1 => n39756, B2 => n29709, C1 => n39750, C2 =>
                           n29773, A => n34177, ZN => n34174);
   U32246 : OAI222_X1 port map( A1 => n31837, A2 => n39744, B1 => n31897, B2 =>
                           n39738, C1 => n31777, C2 => n39732, ZN => n34177);
   U32247 : AOI221_X1 port map( B1 => n39504, B2 => n29709, C1 => n39498, C2 =>
                           n29773, A => n35451, ZN => n35448);
   U32248 : OAI222_X1 port map( A1 => n31837, A2 => n39492, B1 => n31897, B2 =>
                           n39486, C1 => n31777, C2 => n39480, ZN => n35451);
   U32249 : AOI221_X1 port map( B1 => n39756, B2 => n29708, C1 => n39750, C2 =>
                           n29772, A => n34196, ZN => n34193);
   U32250 : OAI222_X1 port map( A1 => n31836, A2 => n39744, B1 => n31896, B2 =>
                           n39738, C1 => n31776, C2 => n39732, ZN => n34196);
   U32251 : AOI221_X1 port map( B1 => n39504, B2 => n29708, C1 => n39498, C2 =>
                           n29772, A => n35470, ZN => n35467);
   U32252 : OAI222_X1 port map( A1 => n31836, A2 => n39492, B1 => n31896, B2 =>
                           n39486, C1 => n31776, C2 => n39480, ZN => n35470);
   U32253 : AOI221_X1 port map( B1 => n39756, B2 => n29707, C1 => n39750, C2 =>
                           n29771, A => n34215, ZN => n34212);
   U32254 : OAI222_X1 port map( A1 => n31835, A2 => n39744, B1 => n31895, B2 =>
                           n39738, C1 => n31775, C2 => n39732, ZN => n34215);
   U32255 : AOI221_X1 port map( B1 => n39504, B2 => n29707, C1 => n39498, C2 =>
                           n29771, A => n35489, ZN => n35486);
   U32256 : OAI222_X1 port map( A1 => n31835, A2 => n39492, B1 => n31895, B2 =>
                           n39486, C1 => n31775, C2 => n39480, ZN => n35489);
   U32257 : AOI221_X1 port map( B1 => n39755, B2 => n29706, C1 => n39749, C2 =>
                           n29770, A => n34234, ZN => n34231);
   U32258 : OAI222_X1 port map( A1 => n31834, A2 => n39743, B1 => n31894, B2 =>
                           n39737, C1 => n31774, C2 => n39731, ZN => n34234);
   U32259 : AOI221_X1 port map( B1 => n39503, B2 => n29706, C1 => n39497, C2 =>
                           n29770, A => n35508, ZN => n35505);
   U32260 : OAI222_X1 port map( A1 => n31834, A2 => n39491, B1 => n31894, B2 =>
                           n39485, C1 => n31774, C2 => n39479, ZN => n35508);
   U32261 : AOI221_X1 port map( B1 => n39755, B2 => n29705, C1 => n39749, C2 =>
                           n29769, A => n34253, ZN => n34250);
   U32262 : OAI222_X1 port map( A1 => n31833, A2 => n39743, B1 => n31893, B2 =>
                           n39737, C1 => n31773, C2 => n39731, ZN => n34253);
   U32263 : AOI221_X1 port map( B1 => n39503, B2 => n29705, C1 => n39497, C2 =>
                           n29769, A => n35527, ZN => n35524);
   U32264 : OAI222_X1 port map( A1 => n31833, A2 => n39491, B1 => n31893, B2 =>
                           n39485, C1 => n31773, C2 => n39479, ZN => n35527);
   U32265 : AOI221_X1 port map( B1 => n39755, B2 => n29704, C1 => n39749, C2 =>
                           n29768, A => n34272, ZN => n34269);
   U32266 : OAI222_X1 port map( A1 => n31832, A2 => n39743, B1 => n31892, B2 =>
                           n39737, C1 => n31772, C2 => n39731, ZN => n34272);
   U32267 : AOI221_X1 port map( B1 => n39503, B2 => n29704, C1 => n39497, C2 =>
                           n29768, A => n35546, ZN => n35543);
   U32268 : OAI222_X1 port map( A1 => n31832, A2 => n39491, B1 => n31892, B2 =>
                           n39485, C1 => n31772, C2 => n39479, ZN => n35546);
   U32269 : AOI221_X1 port map( B1 => n39755, B2 => n29703, C1 => n39749, C2 =>
                           n29767, A => n34291, ZN => n34288);
   U32270 : OAI222_X1 port map( A1 => n31831, A2 => n39743, B1 => n31891, B2 =>
                           n39737, C1 => n31771, C2 => n39731, ZN => n34291);
   U32271 : AOI221_X1 port map( B1 => n39503, B2 => n29703, C1 => n39497, C2 =>
                           n29767, A => n35565, ZN => n35562);
   U32272 : OAI222_X1 port map( A1 => n31831, A2 => n39491, B1 => n31891, B2 =>
                           n39485, C1 => n31771, C2 => n39479, ZN => n35565);
   U32273 : AOI221_X1 port map( B1 => n39755, B2 => n29702, C1 => n39749, C2 =>
                           n29766, A => n34310, ZN => n34307);
   U32274 : OAI222_X1 port map( A1 => n31830, A2 => n39743, B1 => n31890, B2 =>
                           n39737, C1 => n31770, C2 => n39731, ZN => n34310);
   U32275 : AOI221_X1 port map( B1 => n39503, B2 => n29702, C1 => n39497, C2 =>
                           n29766, A => n35584, ZN => n35581);
   U32276 : OAI222_X1 port map( A1 => n31830, A2 => n39491, B1 => n31890, B2 =>
                           n39485, C1 => n31770, C2 => n39479, ZN => n35584);
   U32277 : AOI221_X1 port map( B1 => n39755, B2 => n29701, C1 => n39749, C2 =>
                           n29765, A => n34329, ZN => n34326);
   U32278 : OAI222_X1 port map( A1 => n31829, A2 => n39743, B1 => n31889, B2 =>
                           n39737, C1 => n31769, C2 => n39731, ZN => n34329);
   U32279 : AOI221_X1 port map( B1 => n39503, B2 => n29701, C1 => n39497, C2 =>
                           n29765, A => n35603, ZN => n35600);
   U32280 : OAI222_X1 port map( A1 => n31829, A2 => n39491, B1 => n31889, B2 =>
                           n39485, C1 => n31769, C2 => n39479, ZN => n35603);
   U32281 : AOI221_X1 port map( B1 => n39755, B2 => n29700, C1 => n39749, C2 =>
                           n29764, A => n34348, ZN => n34345);
   U32282 : OAI222_X1 port map( A1 => n31828, A2 => n39743, B1 => n31888, B2 =>
                           n39737, C1 => n31768, C2 => n39731, ZN => n34348);
   U32283 : AOI221_X1 port map( B1 => n39503, B2 => n29700, C1 => n39497, C2 =>
                           n29764, A => n35622, ZN => n35619);
   U32284 : OAI222_X1 port map( A1 => n31828, A2 => n39491, B1 => n31888, B2 =>
                           n39485, C1 => n31768, C2 => n39479, ZN => n35622);
   U32285 : AOI221_X1 port map( B1 => n39755, B2 => n29699, C1 => n39749, C2 =>
                           n29763, A => n34367, ZN => n34364);
   U32286 : OAI222_X1 port map( A1 => n31827, A2 => n39743, B1 => n31887, B2 =>
                           n39737, C1 => n31767, C2 => n39731, ZN => n34367);
   U32287 : AOI221_X1 port map( B1 => n39503, B2 => n29699, C1 => n39497, C2 =>
                           n29763, A => n35641, ZN => n35638);
   U32288 : OAI222_X1 port map( A1 => n31827, A2 => n39491, B1 => n31887, B2 =>
                           n39485, C1 => n31767, C2 => n39479, ZN => n35641);
   U32289 : AOI221_X1 port map( B1 => n39755, B2 => n29698, C1 => n39749, C2 =>
                           n29762, A => n34386, ZN => n34383);
   U32290 : OAI222_X1 port map( A1 => n31826, A2 => n39743, B1 => n31886, B2 =>
                           n39737, C1 => n31766, C2 => n39731, ZN => n34386);
   U32291 : AOI221_X1 port map( B1 => n39503, B2 => n29698, C1 => n39497, C2 =>
                           n29762, A => n35660, ZN => n35657);
   U32292 : OAI222_X1 port map( A1 => n31826, A2 => n39491, B1 => n31886, B2 =>
                           n39485, C1 => n31766, C2 => n39479, ZN => n35660);
   U32293 : AOI221_X1 port map( B1 => n39755, B2 => n29697, C1 => n39749, C2 =>
                           n29761, A => n34405, ZN => n34402);
   U32294 : OAI222_X1 port map( A1 => n31825, A2 => n39743, B1 => n31885, B2 =>
                           n39737, C1 => n31765, C2 => n39731, ZN => n34405);
   U32295 : AOI221_X1 port map( B1 => n39503, B2 => n29697, C1 => n39497, C2 =>
                           n29761, A => n35679, ZN => n35676);
   U32296 : OAI222_X1 port map( A1 => n31825, A2 => n39491, B1 => n31885, B2 =>
                           n39485, C1 => n31765, C2 => n39479, ZN => n35679);
   U32297 : AOI221_X1 port map( B1 => n39755, B2 => n29696, C1 => n39749, C2 =>
                           n29760, A => n34424, ZN => n34421);
   U32298 : OAI222_X1 port map( A1 => n31824, A2 => n39743, B1 => n31884, B2 =>
                           n39737, C1 => n31764, C2 => n39731, ZN => n34424);
   U32299 : AOI221_X1 port map( B1 => n39503, B2 => n29696, C1 => n39497, C2 =>
                           n29760, A => n35698, ZN => n35695);
   U32300 : OAI222_X1 port map( A1 => n31824, A2 => n39491, B1 => n31884, B2 =>
                           n39485, C1 => n31764, C2 => n39479, ZN => n35698);
   U32301 : AOI221_X1 port map( B1 => n39755, B2 => n29695, C1 => n39749, C2 =>
                           n29759, A => n34443, ZN => n34440);
   U32302 : OAI222_X1 port map( A1 => n31823, A2 => n39743, B1 => n31883, B2 =>
                           n39737, C1 => n31763, C2 => n39731, ZN => n34443);
   U32303 : AOI221_X1 port map( B1 => n39503, B2 => n29695, C1 => n39497, C2 =>
                           n29759, A => n35717, ZN => n35714);
   U32304 : OAI222_X1 port map( A1 => n31823, A2 => n39491, B1 => n31883, B2 =>
                           n39485, C1 => n31763, C2 => n39479, ZN => n35717);
   U32305 : AOI221_X1 port map( B1 => n39754, B2 => n29694, C1 => n39748, C2 =>
                           n29758, A => n34462, ZN => n34459);
   U32306 : OAI222_X1 port map( A1 => n31822, A2 => n39742, B1 => n31882, B2 =>
                           n39736, C1 => n31762, C2 => n39730, ZN => n34462);
   U32307 : AOI221_X1 port map( B1 => n39502, B2 => n29694, C1 => n39496, C2 =>
                           n29758, A => n35736, ZN => n35733);
   U32308 : OAI222_X1 port map( A1 => n31822, A2 => n39490, B1 => n31882, B2 =>
                           n39484, C1 => n31762, C2 => n39478, ZN => n35736);
   U32309 : AOI221_X1 port map( B1 => n39754, B2 => n29693, C1 => n39748, C2 =>
                           n29757, A => n34481, ZN => n34478);
   U32310 : OAI222_X1 port map( A1 => n31821, A2 => n39742, B1 => n31881, B2 =>
                           n39736, C1 => n31761, C2 => n39730, ZN => n34481);
   U32311 : AOI221_X1 port map( B1 => n39502, B2 => n29693, C1 => n39496, C2 =>
                           n29757, A => n35755, ZN => n35752);
   U32312 : OAI222_X1 port map( A1 => n31821, A2 => n39490, B1 => n31881, B2 =>
                           n39484, C1 => n31761, C2 => n39478, ZN => n35755);
   U32313 : AOI221_X1 port map( B1 => n39754, B2 => n29692, C1 => n39748, C2 =>
                           n29756, A => n34500, ZN => n34497);
   U32314 : OAI222_X1 port map( A1 => n31820, A2 => n39742, B1 => n31880, B2 =>
                           n39736, C1 => n31760, C2 => n39730, ZN => n34500);
   U32315 : AOI221_X1 port map( B1 => n39502, B2 => n29692, C1 => n39496, C2 =>
                           n29756, A => n35774, ZN => n35771);
   U32316 : OAI222_X1 port map( A1 => n31820, A2 => n39490, B1 => n31880, B2 =>
                           n39484, C1 => n31760, C2 => n39478, ZN => n35774);
   U32317 : AOI221_X1 port map( B1 => n39754, B2 => n29691, C1 => n39748, C2 =>
                           n29755, A => n34519, ZN => n34516);
   U32318 : OAI222_X1 port map( A1 => n31819, A2 => n39742, B1 => n31879, B2 =>
                           n39736, C1 => n31759, C2 => n39730, ZN => n34519);
   U32319 : AOI221_X1 port map( B1 => n39502, B2 => n29691, C1 => n39496, C2 =>
                           n29755, A => n35793, ZN => n35790);
   U32320 : OAI222_X1 port map( A1 => n31819, A2 => n39490, B1 => n31879, B2 =>
                           n39484, C1 => n31759, C2 => n39478, ZN => n35793);
   U32321 : AOI221_X1 port map( B1 => n39754, B2 => n29690, C1 => n39748, C2 =>
                           n29754, A => n34538, ZN => n34535);
   U32322 : OAI222_X1 port map( A1 => n31818, A2 => n39742, B1 => n31878, B2 =>
                           n39736, C1 => n31758, C2 => n39730, ZN => n34538);
   U32323 : AOI221_X1 port map( B1 => n39502, B2 => n29690, C1 => n39496, C2 =>
                           n29754, A => n35812, ZN => n35809);
   U32324 : OAI222_X1 port map( A1 => n31818, A2 => n39490, B1 => n31878, B2 =>
                           n39484, C1 => n31758, C2 => n39478, ZN => n35812);
   U32325 : AOI221_X1 port map( B1 => n39754, B2 => n29689, C1 => n39748, C2 =>
                           n29753, A => n34557, ZN => n34554);
   U32326 : OAI222_X1 port map( A1 => n31817, A2 => n39742, B1 => n31877, B2 =>
                           n39736, C1 => n31757, C2 => n39730, ZN => n34557);
   U32327 : AOI221_X1 port map( B1 => n39502, B2 => n29689, C1 => n39496, C2 =>
                           n29753, A => n35831, ZN => n35828);
   U32328 : OAI222_X1 port map( A1 => n31817, A2 => n39490, B1 => n31877, B2 =>
                           n39484, C1 => n31757, C2 => n39478, ZN => n35831);
   U32329 : AOI221_X1 port map( B1 => n39754, B2 => n29688, C1 => n39748, C2 =>
                           n29752, A => n34576, ZN => n34573);
   U32330 : OAI222_X1 port map( A1 => n31816, A2 => n39742, B1 => n31876, B2 =>
                           n39736, C1 => n31756, C2 => n39730, ZN => n34576);
   U32331 : AOI221_X1 port map( B1 => n39502, B2 => n29688, C1 => n39496, C2 =>
                           n29752, A => n35850, ZN => n35847);
   U32332 : OAI222_X1 port map( A1 => n31816, A2 => n39490, B1 => n31876, B2 =>
                           n39484, C1 => n31756, C2 => n39478, ZN => n35850);
   U32333 : AOI221_X1 port map( B1 => n39754, B2 => n29687, C1 => n39748, C2 =>
                           n29751, A => n34595, ZN => n34592);
   U32334 : OAI222_X1 port map( A1 => n31815, A2 => n39742, B1 => n31875, B2 =>
                           n39736, C1 => n31755, C2 => n39730, ZN => n34595);
   U32335 : AOI221_X1 port map( B1 => n39502, B2 => n29687, C1 => n39496, C2 =>
                           n29751, A => n35869, ZN => n35866);
   U32336 : OAI222_X1 port map( A1 => n31815, A2 => n39490, B1 => n31875, B2 =>
                           n39484, C1 => n31755, C2 => n39478, ZN => n35869);
   U32337 : AOI221_X1 port map( B1 => n39754, B2 => n29686, C1 => n39748, C2 =>
                           n29750, A => n34614, ZN => n34611);
   U32338 : OAI222_X1 port map( A1 => n31814, A2 => n39742, B1 => n31874, B2 =>
                           n39736, C1 => n31754, C2 => n39730, ZN => n34614);
   U32339 : AOI221_X1 port map( B1 => n39502, B2 => n29686, C1 => n39496, C2 =>
                           n29750, A => n35888, ZN => n35885);
   U32340 : OAI222_X1 port map( A1 => n31814, A2 => n39490, B1 => n31874, B2 =>
                           n39484, C1 => n31754, C2 => n39478, ZN => n35888);
   U32341 : AOI221_X1 port map( B1 => n39754, B2 => n29685, C1 => n39748, C2 =>
                           n29749, A => n34633, ZN => n34630);
   U32342 : OAI222_X1 port map( A1 => n31813, A2 => n39742, B1 => n31873, B2 =>
                           n39736, C1 => n31753, C2 => n39730, ZN => n34633);
   U32343 : AOI221_X1 port map( B1 => n39502, B2 => n29685, C1 => n39496, C2 =>
                           n29749, A => n35907, ZN => n35904);
   U32344 : OAI222_X1 port map( A1 => n31813, A2 => n39490, B1 => n31873, B2 =>
                           n39484, C1 => n31753, C2 => n39478, ZN => n35907);
   U32345 : AOI221_X1 port map( B1 => n39754, B2 => n29684, C1 => n39748, C2 =>
                           n29748, A => n34652, ZN => n34649);
   U32346 : OAI222_X1 port map( A1 => n31812, A2 => n39742, B1 => n31872, B2 =>
                           n39736, C1 => n31752, C2 => n39730, ZN => n34652);
   U32347 : AOI221_X1 port map( B1 => n39502, B2 => n29684, C1 => n39496, C2 =>
                           n29748, A => n35926, ZN => n35923);
   U32348 : OAI222_X1 port map( A1 => n31812, A2 => n39490, B1 => n31872, B2 =>
                           n39484, C1 => n31752, C2 => n39478, ZN => n35926);
   U32349 : AOI221_X1 port map( B1 => n39754, B2 => n29683, C1 => n39748, C2 =>
                           n29747, A => n34677, ZN => n34668);
   U32350 : OAI222_X1 port map( A1 => n31811, A2 => n39742, B1 => n31871, B2 =>
                           n39736, C1 => n31751, C2 => n39730, ZN => n34677);
   U32351 : AOI221_X1 port map( B1 => n39502, B2 => n29683, C1 => n39496, C2 =>
                           n29747, A => n35951, ZN => n35942);
   U32352 : OAI222_X1 port map( A1 => n31811, A2 => n39490, B1 => n31871, B2 =>
                           n39484, C1 => n31751, C2 => n39478, ZN => n35951);
   U32353 : OAI222_X1 port map( A1 => n40910, A2 => n39914, B1 => n41294, B2 =>
                           n39907, C1 => n390, C2 => n39901, ZN => n7662);
   U32354 : OAI222_X1 port map( A1 => n40916, A2 => n39914, B1 => n41300, B2 =>
                           n39907, C1 => n389, C2 => n39901, ZN => n7661);
   U32355 : OAI222_X1 port map( A1 => n40922, A2 => n39914, B1 => n41306, B2 =>
                           n39907, C1 => n388, C2 => n39901, ZN => n7660);
   U32356 : OAI222_X1 port map( A1 => n40928, A2 => n39914, B1 => n41312, B2 =>
                           n39907, C1 => n387, C2 => n39901, ZN => n7659);
   U32357 : OAI222_X1 port map( A1 => n40934, A2 => n39914, B1 => n41318, B2 =>
                           n39907, C1 => n386, C2 => n39901, ZN => n7658);
   U32358 : OAI222_X1 port map( A1 => n40940, A2 => n39914, B1 => n41324, B2 =>
                           n39907, C1 => n385, C2 => n39901, ZN => n7657);
   U32359 : OAI222_X1 port map( A1 => n40946, A2 => n39914, B1 => n41330, B2 =>
                           n39907, C1 => n384, C2 => n39901, ZN => n7656);
   U32360 : OAI222_X1 port map( A1 => n40952, A2 => n39914, B1 => n41336, B2 =>
                           n39907, C1 => n383, C2 => n39901, ZN => n7655);
   U32361 : OAI222_X1 port map( A1 => n40958, A2 => n39914, B1 => n41342, B2 =>
                           n39907, C1 => n382, C2 => n39901, ZN => n7654);
   U32362 : OAI222_X1 port map( A1 => n40964, A2 => n39914, B1 => n41348, B2 =>
                           n39907, C1 => n381, C2 => n39901, ZN => n7653);
   U32363 : OAI222_X1 port map( A1 => n40970, A2 => n39914, B1 => n41354, B2 =>
                           n39907, C1 => n380, C2 => n39901, ZN => n7652);
   U32364 : OAI222_X1 port map( A1 => n40976, A2 => n39914, B1 => n41360, B2 =>
                           n39907, C1 => n379, C2 => n39901, ZN => n7651);
   U32365 : OAI222_X1 port map( A1 => n40910, A2 => n39933, B1 => n41294, B2 =>
                           n39926, C1 => n454, C2 => n39920, ZN => n7726);
   U32366 : OAI222_X1 port map( A1 => n40916, A2 => n39933, B1 => n41300, B2 =>
                           n39926, C1 => n453, C2 => n39920, ZN => n7725);
   U32367 : OAI222_X1 port map( A1 => n40922, A2 => n39933, B1 => n41306, B2 =>
                           n39926, C1 => n452, C2 => n39920, ZN => n7724);
   U32368 : OAI222_X1 port map( A1 => n40928, A2 => n39933, B1 => n41312, B2 =>
                           n39926, C1 => n451, C2 => n39920, ZN => n7723);
   U32369 : OAI222_X1 port map( A1 => n40934, A2 => n39933, B1 => n41318, B2 =>
                           n39926, C1 => n450, C2 => n39920, ZN => n7722);
   U32370 : OAI222_X1 port map( A1 => n40940, A2 => n39933, B1 => n41324, B2 =>
                           n39926, C1 => n449, C2 => n39920, ZN => n7721);
   U32371 : OAI222_X1 port map( A1 => n40946, A2 => n39933, B1 => n41330, B2 =>
                           n39926, C1 => n448, C2 => n39920, ZN => n7720);
   U32372 : OAI222_X1 port map( A1 => n40952, A2 => n39933, B1 => n41336, B2 =>
                           n39926, C1 => n447, C2 => n39920, ZN => n7719);
   U32373 : OAI222_X1 port map( A1 => n40958, A2 => n39933, B1 => n41342, B2 =>
                           n39926, C1 => n446, C2 => n39920, ZN => n7718);
   U32374 : OAI222_X1 port map( A1 => n40964, A2 => n39933, B1 => n41348, B2 =>
                           n39926, C1 => n445, C2 => n39920, ZN => n7717);
   U32375 : OAI222_X1 port map( A1 => n40970, A2 => n39933, B1 => n41354, B2 =>
                           n39926, C1 => n444, C2 => n39920, ZN => n7716);
   U32376 : OAI222_X1 port map( A1 => n40976, A2 => n39933, B1 => n41360, B2 =>
                           n39926, C1 => n443, C2 => n39920, ZN => n7715);
   U32377 : OAI222_X1 port map( A1 => n40622, A2 => n39918, B1 => n41006, B2 =>
                           n39911, C1 => n438, C2 => n39905, ZN => n7710);
   U32378 : OAI222_X1 port map( A1 => n40628, A2 => n39918, B1 => n41012, B2 =>
                           n39911, C1 => n437, C2 => n39905, ZN => n7709);
   U32379 : OAI222_X1 port map( A1 => n40634, A2 => n39918, B1 => n41018, B2 =>
                           n39911, C1 => n436, C2 => n39905, ZN => n7708);
   U32380 : OAI222_X1 port map( A1 => n40640, A2 => n39918, B1 => n41024, B2 =>
                           n39911, C1 => n435, C2 => n39905, ZN => n7707);
   U32381 : OAI222_X1 port map( A1 => n40646, A2 => n39918, B1 => n41030, B2 =>
                           n39911, C1 => n434, C2 => n39905, ZN => n7706);
   U32382 : OAI222_X1 port map( A1 => n40652, A2 => n39918, B1 => n41036, B2 =>
                           n39911, C1 => n433, C2 => n39905, ZN => n7705);
   U32383 : OAI222_X1 port map( A1 => n40658, A2 => n39918, B1 => n41042, B2 =>
                           n39911, C1 => n432, C2 => n39905, ZN => n7704);
   U32384 : OAI222_X1 port map( A1 => n40664, A2 => n39918, B1 => n41048, B2 =>
                           n39911, C1 => n431, C2 => n39905, ZN => n7703);
   U32385 : OAI222_X1 port map( A1 => n40670, A2 => n39918, B1 => n41054, B2 =>
                           n39911, C1 => n430, C2 => n39905, ZN => n7702);
   U32386 : OAI222_X1 port map( A1 => n40676, A2 => n39918, B1 => n41060, B2 =>
                           n39911, C1 => n429, C2 => n39904, ZN => n7701);
   U32387 : OAI222_X1 port map( A1 => n40682, A2 => n39918, B1 => n41066, B2 =>
                           n39911, C1 => n428, C2 => n39904, ZN => n7700);
   U32388 : OAI222_X1 port map( A1 => n40688, A2 => n39918, B1 => n41072, B2 =>
                           n39911, C1 => n427, C2 => n39904, ZN => n7699);
   U32389 : OAI222_X1 port map( A1 => n40694, A2 => n39917, B1 => n41078, B2 =>
                           n39910, C1 => n426, C2 => n39904, ZN => n7698);
   U32390 : OAI222_X1 port map( A1 => n40700, A2 => n39917, B1 => n41084, B2 =>
                           n39910, C1 => n425, C2 => n39904, ZN => n7697);
   U32391 : OAI222_X1 port map( A1 => n40706, A2 => n39917, B1 => n41090, B2 =>
                           n39910, C1 => n424, C2 => n39904, ZN => n7696);
   U32392 : OAI222_X1 port map( A1 => n40712, A2 => n39917, B1 => n41096, B2 =>
                           n39910, C1 => n423, C2 => n39904, ZN => n7695);
   U32393 : OAI222_X1 port map( A1 => n40718, A2 => n39917, B1 => n41102, B2 =>
                           n39910, C1 => n422, C2 => n39904, ZN => n7694);
   U32394 : OAI222_X1 port map( A1 => n40724, A2 => n39917, B1 => n41108, B2 =>
                           n39910, C1 => n421, C2 => n39904, ZN => n7693);
   U32395 : OAI222_X1 port map( A1 => n40730, A2 => n39917, B1 => n41114, B2 =>
                           n39910, C1 => n420, C2 => n39904, ZN => n7692);
   U32396 : OAI222_X1 port map( A1 => n40736, A2 => n39917, B1 => n41120, B2 =>
                           n39910, C1 => n419, C2 => n39904, ZN => n7691);
   U32397 : OAI222_X1 port map( A1 => n40742, A2 => n39917, B1 => n41126, B2 =>
                           n39910, C1 => n418, C2 => n39904, ZN => n7690);
   U32398 : OAI222_X1 port map( A1 => n40748, A2 => n39917, B1 => n41132, B2 =>
                           n39910, C1 => n417, C2 => n39904, ZN => n7689);
   U32399 : OAI222_X1 port map( A1 => n40754, A2 => n39917, B1 => n41138, B2 =>
                           n39910, C1 => n416, C2 => n39903, ZN => n7688);
   U32400 : OAI222_X1 port map( A1 => n40760, A2 => n39917, B1 => n41144, B2 =>
                           n39910, C1 => n415, C2 => n39903, ZN => n7687);
   U32401 : OAI222_X1 port map( A1 => n40766, A2 => n39916, B1 => n41150, B2 =>
                           n39909, C1 => n414, C2 => n39903, ZN => n7686);
   U32402 : OAI222_X1 port map( A1 => n40772, A2 => n39916, B1 => n41156, B2 =>
                           n39909, C1 => n413, C2 => n39903, ZN => n7685);
   U32403 : OAI222_X1 port map( A1 => n40778, A2 => n39916, B1 => n41162, B2 =>
                           n39909, C1 => n412, C2 => n39903, ZN => n7684);
   U32404 : OAI222_X1 port map( A1 => n40784, A2 => n39916, B1 => n41168, B2 =>
                           n39909, C1 => n411, C2 => n39903, ZN => n7683);
   U32405 : OAI222_X1 port map( A1 => n40790, A2 => n39916, B1 => n41174, B2 =>
                           n39909, C1 => n410, C2 => n39903, ZN => n7682);
   U32406 : OAI222_X1 port map( A1 => n40796, A2 => n39916, B1 => n41180, B2 =>
                           n39909, C1 => n409, C2 => n39903, ZN => n7681);
   U32407 : OAI222_X1 port map( A1 => n40802, A2 => n39916, B1 => n41186, B2 =>
                           n39909, C1 => n408, C2 => n39903, ZN => n7680);
   U32408 : OAI222_X1 port map( A1 => n40808, A2 => n39916, B1 => n41192, B2 =>
                           n39909, C1 => n407, C2 => n39903, ZN => n7679);
   U32409 : OAI222_X1 port map( A1 => n40814, A2 => n39916, B1 => n41198, B2 =>
                           n39909, C1 => n406, C2 => n39903, ZN => n7678);
   U32410 : OAI222_X1 port map( A1 => n40820, A2 => n39916, B1 => n41204, B2 =>
                           n39909, C1 => n405, C2 => n39903, ZN => n7677);
   U32411 : OAI222_X1 port map( A1 => n40826, A2 => n39916, B1 => n41210, B2 =>
                           n39909, C1 => n404, C2 => n39903, ZN => n7676);
   U32412 : OAI222_X1 port map( A1 => n40832, A2 => n39916, B1 => n41216, B2 =>
                           n39909, C1 => n403, C2 => n39902, ZN => n7675);
   U32413 : OAI222_X1 port map( A1 => n40838, A2 => n39915, B1 => n41222, B2 =>
                           n39908, C1 => n402, C2 => n39902, ZN => n7674);
   U32414 : OAI222_X1 port map( A1 => n40844, A2 => n39915, B1 => n41228, B2 =>
                           n39908, C1 => n401, C2 => n39902, ZN => n7673);
   U32415 : OAI222_X1 port map( A1 => n40850, A2 => n39915, B1 => n41234, B2 =>
                           n39908, C1 => n400, C2 => n39902, ZN => n7672);
   U32416 : OAI222_X1 port map( A1 => n40856, A2 => n39915, B1 => n41240, B2 =>
                           n39908, C1 => n399, C2 => n39902, ZN => n7671);
   U32417 : OAI222_X1 port map( A1 => n40862, A2 => n39915, B1 => n41246, B2 =>
                           n39908, C1 => n398, C2 => n39902, ZN => n7670);
   U32418 : OAI222_X1 port map( A1 => n40868, A2 => n39915, B1 => n41252, B2 =>
                           n39908, C1 => n397, C2 => n39902, ZN => n7669);
   U32419 : OAI222_X1 port map( A1 => n40874, A2 => n39915, B1 => n41258, B2 =>
                           n39908, C1 => n396, C2 => n39902, ZN => n7668);
   U32420 : OAI222_X1 port map( A1 => n40880, A2 => n39915, B1 => n41264, B2 =>
                           n39908, C1 => n395, C2 => n39902, ZN => n7667);
   U32421 : OAI222_X1 port map( A1 => n40886, A2 => n39915, B1 => n41270, B2 =>
                           n39908, C1 => n394, C2 => n39902, ZN => n7666);
   U32422 : OAI222_X1 port map( A1 => n40892, A2 => n39915, B1 => n41276, B2 =>
                           n39908, C1 => n393, C2 => n39902, ZN => n7665);
   U32423 : OAI222_X1 port map( A1 => n40898, A2 => n39915, B1 => n41282, B2 =>
                           n39908, C1 => n392, C2 => n39902, ZN => n7664);
   U32424 : OAI222_X1 port map( A1 => n40904, A2 => n39915, B1 => n41288, B2 =>
                           n39908, C1 => n391, C2 => n39902, ZN => n7663);
   U32425 : OAI222_X1 port map( A1 => n40622, A2 => n39937, B1 => n41006, B2 =>
                           n39930, C1 => n502, C2 => n39924, ZN => n7774);
   U32426 : OAI222_X1 port map( A1 => n40628, A2 => n39937, B1 => n41012, B2 =>
                           n39930, C1 => n501, C2 => n39924, ZN => n7773);
   U32427 : OAI222_X1 port map( A1 => n40634, A2 => n39937, B1 => n41018, B2 =>
                           n39930, C1 => n500, C2 => n39924, ZN => n7772);
   U32428 : OAI222_X1 port map( A1 => n40640, A2 => n39937, B1 => n41024, B2 =>
                           n39930, C1 => n499, C2 => n39924, ZN => n7771);
   U32429 : OAI222_X1 port map( A1 => n40646, A2 => n39937, B1 => n41030, B2 =>
                           n39930, C1 => n498, C2 => n39924, ZN => n7770);
   U32430 : OAI222_X1 port map( A1 => n40652, A2 => n39937, B1 => n41036, B2 =>
                           n39930, C1 => n497, C2 => n39924, ZN => n7769);
   U32431 : OAI222_X1 port map( A1 => n40658, A2 => n39937, B1 => n41042, B2 =>
                           n39930, C1 => n496, C2 => n39924, ZN => n7768);
   U32432 : OAI222_X1 port map( A1 => n40664, A2 => n39937, B1 => n41048, B2 =>
                           n39930, C1 => n495, C2 => n39924, ZN => n7767);
   U32433 : OAI222_X1 port map( A1 => n40670, A2 => n39937, B1 => n41054, B2 =>
                           n39930, C1 => n494, C2 => n39924, ZN => n7766);
   U32434 : OAI222_X1 port map( A1 => n40676, A2 => n39937, B1 => n41060, B2 =>
                           n39930, C1 => n493, C2 => n39923, ZN => n7765);
   U32435 : OAI222_X1 port map( A1 => n40682, A2 => n39937, B1 => n41066, B2 =>
                           n39930, C1 => n492, C2 => n39923, ZN => n7764);
   U32436 : OAI222_X1 port map( A1 => n40688, A2 => n39937, B1 => n41072, B2 =>
                           n39930, C1 => n491, C2 => n39923, ZN => n7763);
   U32437 : OAI222_X1 port map( A1 => n40694, A2 => n39936, B1 => n41078, B2 =>
                           n39929, C1 => n490, C2 => n39923, ZN => n7762);
   U32438 : OAI222_X1 port map( A1 => n40700, A2 => n39936, B1 => n41084, B2 =>
                           n39929, C1 => n489, C2 => n39923, ZN => n7761);
   U32439 : OAI222_X1 port map( A1 => n40706, A2 => n39936, B1 => n41090, B2 =>
                           n39929, C1 => n488, C2 => n39923, ZN => n7760);
   U32440 : OAI222_X1 port map( A1 => n40712, A2 => n39936, B1 => n41096, B2 =>
                           n39929, C1 => n487, C2 => n39923, ZN => n7759);
   U32441 : OAI222_X1 port map( A1 => n40718, A2 => n39936, B1 => n41102, B2 =>
                           n39929, C1 => n486, C2 => n39923, ZN => n7758);
   U32442 : OAI222_X1 port map( A1 => n40724, A2 => n39936, B1 => n41108, B2 =>
                           n39929, C1 => n485, C2 => n39923, ZN => n7757);
   U32443 : OAI222_X1 port map( A1 => n40730, A2 => n39936, B1 => n41114, B2 =>
                           n39929, C1 => n484, C2 => n39923, ZN => n7756);
   U32444 : OAI222_X1 port map( A1 => n40736, A2 => n39936, B1 => n41120, B2 =>
                           n39929, C1 => n483, C2 => n39923, ZN => n7755);
   U32445 : OAI222_X1 port map( A1 => n40742, A2 => n39936, B1 => n41126, B2 =>
                           n39929, C1 => n482, C2 => n39923, ZN => n7754);
   U32446 : OAI222_X1 port map( A1 => n40748, A2 => n39936, B1 => n41132, B2 =>
                           n39929, C1 => n481, C2 => n39923, ZN => n7753);
   U32447 : OAI222_X1 port map( A1 => n40754, A2 => n39936, B1 => n41138, B2 =>
                           n39929, C1 => n480, C2 => n39922, ZN => n7752);
   U32448 : OAI222_X1 port map( A1 => n40760, A2 => n39936, B1 => n41144, B2 =>
                           n39929, C1 => n479, C2 => n39922, ZN => n7751);
   U32449 : OAI222_X1 port map( A1 => n40766, A2 => n39935, B1 => n41150, B2 =>
                           n39928, C1 => n478, C2 => n39922, ZN => n7750);
   U32450 : OAI222_X1 port map( A1 => n40772, A2 => n39935, B1 => n41156, B2 =>
                           n39928, C1 => n477, C2 => n39922, ZN => n7749);
   U32451 : OAI222_X1 port map( A1 => n40778, A2 => n39935, B1 => n41162, B2 =>
                           n39928, C1 => n476, C2 => n39922, ZN => n7748);
   U32452 : OAI222_X1 port map( A1 => n40784, A2 => n39935, B1 => n41168, B2 =>
                           n39928, C1 => n475, C2 => n39922, ZN => n7747);
   U32453 : OAI222_X1 port map( A1 => n40790, A2 => n39935, B1 => n41174, B2 =>
                           n39928, C1 => n474, C2 => n39922, ZN => n7746);
   U32454 : OAI222_X1 port map( A1 => n40796, A2 => n39935, B1 => n41180, B2 =>
                           n39928, C1 => n473, C2 => n39922, ZN => n7745);
   U32455 : OAI222_X1 port map( A1 => n40802, A2 => n39935, B1 => n41186, B2 =>
                           n39928, C1 => n472, C2 => n39922, ZN => n7744);
   U32456 : OAI222_X1 port map( A1 => n40808, A2 => n39935, B1 => n41192, B2 =>
                           n39928, C1 => n471, C2 => n39922, ZN => n7743);
   U32457 : OAI222_X1 port map( A1 => n40814, A2 => n39935, B1 => n41198, B2 =>
                           n39928, C1 => n470, C2 => n39922, ZN => n7742);
   U32458 : OAI222_X1 port map( A1 => n40820, A2 => n39935, B1 => n41204, B2 =>
                           n39928, C1 => n469, C2 => n39922, ZN => n7741);
   U32459 : OAI222_X1 port map( A1 => n40826, A2 => n39935, B1 => n41210, B2 =>
                           n39928, C1 => n468, C2 => n39922, ZN => n7740);
   U32460 : OAI222_X1 port map( A1 => n40832, A2 => n39935, B1 => n41216, B2 =>
                           n39928, C1 => n467, C2 => n39921, ZN => n7739);
   U32461 : OAI222_X1 port map( A1 => n40838, A2 => n39934, B1 => n41222, B2 =>
                           n39927, C1 => n466, C2 => n39921, ZN => n7738);
   U32462 : OAI222_X1 port map( A1 => n40844, A2 => n39934, B1 => n41228, B2 =>
                           n39927, C1 => n465, C2 => n39921, ZN => n7737);
   U32463 : OAI222_X1 port map( A1 => n40850, A2 => n39934, B1 => n41234, B2 =>
                           n39927, C1 => n464, C2 => n39921, ZN => n7736);
   U32464 : OAI222_X1 port map( A1 => n40856, A2 => n39934, B1 => n41240, B2 =>
                           n39927, C1 => n463, C2 => n39921, ZN => n7735);
   U32465 : OAI222_X1 port map( A1 => n40862, A2 => n39934, B1 => n41246, B2 =>
                           n39927, C1 => n462, C2 => n39921, ZN => n7734);
   U32466 : OAI222_X1 port map( A1 => n40868, A2 => n39934, B1 => n41252, B2 =>
                           n39927, C1 => n461, C2 => n39921, ZN => n7733);
   U32467 : OAI222_X1 port map( A1 => n40874, A2 => n39934, B1 => n41258, B2 =>
                           n39927, C1 => n460, C2 => n39921, ZN => n7732);
   U32468 : OAI222_X1 port map( A1 => n40880, A2 => n39934, B1 => n41264, B2 =>
                           n39927, C1 => n459, C2 => n39921, ZN => n7731);
   U32469 : OAI222_X1 port map( A1 => n40886, A2 => n39934, B1 => n41270, B2 =>
                           n39927, C1 => n458, C2 => n39921, ZN => n7730);
   U32470 : OAI222_X1 port map( A1 => n40892, A2 => n39934, B1 => n41276, B2 =>
                           n39927, C1 => n457, C2 => n39921, ZN => n7729);
   U32471 : OAI222_X1 port map( A1 => n40898, A2 => n39934, B1 => n41282, B2 =>
                           n39927, C1 => n456, C2 => n39921, ZN => n7728);
   U32472 : OAI222_X1 port map( A1 => n40904, A2 => n39934, B1 => n41288, B2 =>
                           n39927, C1 => n455, C2 => n39921, ZN => n7727);
   U32473 : OAI222_X1 port map( A1 => n40910, A2 => n40012, B1 => n41294, B2 =>
                           n40005, C1 => n710, C2 => n39999, ZN => n7982);
   U32474 : OAI222_X1 port map( A1 => n40916, A2 => n40012, B1 => n41300, B2 =>
                           n40005, C1 => n709, C2 => n39999, ZN => n7981);
   U32475 : OAI222_X1 port map( A1 => n40922, A2 => n40012, B1 => n41306, B2 =>
                           n40005, C1 => n708, C2 => n39999, ZN => n7980);
   U32476 : OAI222_X1 port map( A1 => n40928, A2 => n40012, B1 => n41312, B2 =>
                           n40005, C1 => n707, C2 => n39999, ZN => n7979);
   U32477 : OAI222_X1 port map( A1 => n40934, A2 => n40012, B1 => n41318, B2 =>
                           n40005, C1 => n706, C2 => n39999, ZN => n7978);
   U32478 : OAI222_X1 port map( A1 => n40940, A2 => n40012, B1 => n41324, B2 =>
                           n40005, C1 => n705, C2 => n39999, ZN => n7977);
   U32479 : OAI222_X1 port map( A1 => n40946, A2 => n40012, B1 => n41330, B2 =>
                           n40005, C1 => n704, C2 => n39999, ZN => n7976);
   U32480 : OAI222_X1 port map( A1 => n40952, A2 => n40012, B1 => n41336, B2 =>
                           n40005, C1 => n703, C2 => n39999, ZN => n7975);
   U32481 : OAI222_X1 port map( A1 => n40958, A2 => n40012, B1 => n41342, B2 =>
                           n40005, C1 => n702, C2 => n39999, ZN => n7974);
   U32482 : OAI222_X1 port map( A1 => n40964, A2 => n40012, B1 => n41348, B2 =>
                           n40005, C1 => n701, C2 => n39999, ZN => n7973);
   U32483 : OAI222_X1 port map( A1 => n40970, A2 => n40012, B1 => n41354, B2 =>
                           n40005, C1 => n700, C2 => n39999, ZN => n7972);
   U32484 : OAI222_X1 port map( A1 => n40976, A2 => n40012, B1 => n41360, B2 =>
                           n40005, C1 => n699, C2 => n39999, ZN => n7971);
   U32485 : OAI222_X1 port map( A1 => n40910, A2 => n40031, B1 => n41294, B2 =>
                           n40024, C1 => n774, C2 => n40018, ZN => n8046);
   U32486 : OAI222_X1 port map( A1 => n40916, A2 => n40031, B1 => n41300, B2 =>
                           n40024, C1 => n773, C2 => n40018, ZN => n8045);
   U32487 : OAI222_X1 port map( A1 => n40922, A2 => n40031, B1 => n41306, B2 =>
                           n40024, C1 => n772, C2 => n40018, ZN => n8044);
   U32488 : OAI222_X1 port map( A1 => n40928, A2 => n40031, B1 => n41312, B2 =>
                           n40024, C1 => n771, C2 => n40018, ZN => n8043);
   U32489 : OAI222_X1 port map( A1 => n40934, A2 => n40031, B1 => n41318, B2 =>
                           n40024, C1 => n770, C2 => n40018, ZN => n8042);
   U32490 : OAI222_X1 port map( A1 => n40940, A2 => n40031, B1 => n41324, B2 =>
                           n40024, C1 => n769, C2 => n40018, ZN => n8041);
   U32491 : OAI222_X1 port map( A1 => n40946, A2 => n40031, B1 => n41330, B2 =>
                           n40024, C1 => n768, C2 => n40018, ZN => n8040);
   U32492 : OAI222_X1 port map( A1 => n40952, A2 => n40031, B1 => n41336, B2 =>
                           n40024, C1 => n767, C2 => n40018, ZN => n8039);
   U32493 : OAI222_X1 port map( A1 => n40958, A2 => n40031, B1 => n41342, B2 =>
                           n40024, C1 => n766, C2 => n40018, ZN => n8038);
   U32494 : OAI222_X1 port map( A1 => n40964, A2 => n40031, B1 => n41348, B2 =>
                           n40024, C1 => n765, C2 => n40018, ZN => n8037);
   U32495 : OAI222_X1 port map( A1 => n40970, A2 => n40031, B1 => n41354, B2 =>
                           n40024, C1 => n764, C2 => n40018, ZN => n8036);
   U32496 : OAI222_X1 port map( A1 => n40976, A2 => n40031, B1 => n41360, B2 =>
                           n40024, C1 => n763, C2 => n40018, ZN => n8035);
   U32497 : OAI222_X1 port map( A1 => n40622, A2 => n40016, B1 => n41006, B2 =>
                           n40009, C1 => n758, C2 => n40003, ZN => n8030);
   U32498 : OAI222_X1 port map( A1 => n40628, A2 => n40016, B1 => n41012, B2 =>
                           n40009, C1 => n757, C2 => n40003, ZN => n8029);
   U32499 : OAI222_X1 port map( A1 => n40634, A2 => n40016, B1 => n41018, B2 =>
                           n40009, C1 => n756, C2 => n40003, ZN => n8028);
   U32500 : OAI222_X1 port map( A1 => n40640, A2 => n40016, B1 => n41024, B2 =>
                           n40009, C1 => n755, C2 => n40003, ZN => n8027);
   U32501 : OAI222_X1 port map( A1 => n40646, A2 => n40016, B1 => n41030, B2 =>
                           n40009, C1 => n754, C2 => n40003, ZN => n8026);
   U32502 : OAI222_X1 port map( A1 => n40652, A2 => n40016, B1 => n41036, B2 =>
                           n40009, C1 => n753, C2 => n40003, ZN => n8025);
   U32503 : OAI222_X1 port map( A1 => n40658, A2 => n40016, B1 => n41042, B2 =>
                           n40009, C1 => n752, C2 => n40003, ZN => n8024);
   U32504 : OAI222_X1 port map( A1 => n40664, A2 => n40016, B1 => n41048, B2 =>
                           n40009, C1 => n751, C2 => n40003, ZN => n8023);
   U32505 : OAI222_X1 port map( A1 => n40670, A2 => n40016, B1 => n41054, B2 =>
                           n40009, C1 => n750, C2 => n40003, ZN => n8022);
   U32506 : OAI222_X1 port map( A1 => n40676, A2 => n40016, B1 => n41060, B2 =>
                           n40009, C1 => n749, C2 => n40002, ZN => n8021);
   U32507 : OAI222_X1 port map( A1 => n40682, A2 => n40016, B1 => n41066, B2 =>
                           n40009, C1 => n748, C2 => n40002, ZN => n8020);
   U32508 : OAI222_X1 port map( A1 => n40688, A2 => n40016, B1 => n41072, B2 =>
                           n40009, C1 => n747, C2 => n40002, ZN => n8019);
   U32509 : OAI222_X1 port map( A1 => n40694, A2 => n40015, B1 => n41078, B2 =>
                           n40008, C1 => n746, C2 => n40002, ZN => n8018);
   U32510 : OAI222_X1 port map( A1 => n40700, A2 => n40015, B1 => n41084, B2 =>
                           n40008, C1 => n745, C2 => n40002, ZN => n8017);
   U32511 : OAI222_X1 port map( A1 => n40706, A2 => n40015, B1 => n41090, B2 =>
                           n40008, C1 => n744, C2 => n40002, ZN => n8016);
   U32512 : OAI222_X1 port map( A1 => n40712, A2 => n40015, B1 => n41096, B2 =>
                           n40008, C1 => n743, C2 => n40002, ZN => n8015);
   U32513 : OAI222_X1 port map( A1 => n40718, A2 => n40015, B1 => n41102, B2 =>
                           n40008, C1 => n742, C2 => n40002, ZN => n8014);
   U32514 : OAI222_X1 port map( A1 => n40724, A2 => n40015, B1 => n41108, B2 =>
                           n40008, C1 => n741, C2 => n40002, ZN => n8013);
   U32515 : OAI222_X1 port map( A1 => n40730, A2 => n40015, B1 => n41114, B2 =>
                           n40008, C1 => n740, C2 => n40002, ZN => n8012);
   U32516 : OAI222_X1 port map( A1 => n40736, A2 => n40015, B1 => n41120, B2 =>
                           n40008, C1 => n739, C2 => n40002, ZN => n8011);
   U32517 : OAI222_X1 port map( A1 => n40742, A2 => n40015, B1 => n41126, B2 =>
                           n40008, C1 => n738, C2 => n40002, ZN => n8010);
   U32518 : OAI222_X1 port map( A1 => n40748, A2 => n40015, B1 => n41132, B2 =>
                           n40008, C1 => n737, C2 => n40002, ZN => n8009);
   U32519 : OAI222_X1 port map( A1 => n40754, A2 => n40015, B1 => n41138, B2 =>
                           n40008, C1 => n736, C2 => n40001, ZN => n8008);
   U32520 : OAI222_X1 port map( A1 => n40760, A2 => n40015, B1 => n41144, B2 =>
                           n40008, C1 => n735, C2 => n40001, ZN => n8007);
   U32521 : OAI222_X1 port map( A1 => n40766, A2 => n40014, B1 => n41150, B2 =>
                           n40007, C1 => n734, C2 => n40001, ZN => n8006);
   U32522 : OAI222_X1 port map( A1 => n40772, A2 => n40014, B1 => n41156, B2 =>
                           n40007, C1 => n733, C2 => n40001, ZN => n8005);
   U32523 : OAI222_X1 port map( A1 => n40778, A2 => n40014, B1 => n41162, B2 =>
                           n40007, C1 => n732, C2 => n40001, ZN => n8004);
   U32524 : OAI222_X1 port map( A1 => n40784, A2 => n40014, B1 => n41168, B2 =>
                           n40007, C1 => n731, C2 => n40001, ZN => n8003);
   U32525 : OAI222_X1 port map( A1 => n40790, A2 => n40014, B1 => n41174, B2 =>
                           n40007, C1 => n730, C2 => n40001, ZN => n8002);
   U32526 : OAI222_X1 port map( A1 => n40796, A2 => n40014, B1 => n41180, B2 =>
                           n40007, C1 => n729, C2 => n40001, ZN => n8001);
   U32527 : OAI222_X1 port map( A1 => n40802, A2 => n40014, B1 => n41186, B2 =>
                           n40007, C1 => n728, C2 => n40001, ZN => n8000);
   U32528 : OAI222_X1 port map( A1 => n40808, A2 => n40014, B1 => n41192, B2 =>
                           n40007, C1 => n727, C2 => n40001, ZN => n7999);
   U32529 : OAI222_X1 port map( A1 => n40814, A2 => n40014, B1 => n41198, B2 =>
                           n40007, C1 => n726, C2 => n40001, ZN => n7998);
   U32530 : OAI222_X1 port map( A1 => n40820, A2 => n40014, B1 => n41204, B2 =>
                           n40007, C1 => n725, C2 => n40001, ZN => n7997);
   U32531 : OAI222_X1 port map( A1 => n40826, A2 => n40014, B1 => n41210, B2 =>
                           n40007, C1 => n724, C2 => n40001, ZN => n7996);
   U32532 : OAI222_X1 port map( A1 => n40832, A2 => n40014, B1 => n41216, B2 =>
                           n40007, C1 => n723, C2 => n40000, ZN => n7995);
   U32533 : OAI222_X1 port map( A1 => n40838, A2 => n40013, B1 => n41222, B2 =>
                           n40006, C1 => n722, C2 => n40000, ZN => n7994);
   U32534 : OAI222_X1 port map( A1 => n40844, A2 => n40013, B1 => n41228, B2 =>
                           n40006, C1 => n721, C2 => n40000, ZN => n7993);
   U32535 : OAI222_X1 port map( A1 => n40850, A2 => n40013, B1 => n41234, B2 =>
                           n40006, C1 => n720, C2 => n40000, ZN => n7992);
   U32536 : OAI222_X1 port map( A1 => n40856, A2 => n40013, B1 => n41240, B2 =>
                           n40006, C1 => n719, C2 => n40000, ZN => n7991);
   U32537 : OAI222_X1 port map( A1 => n40862, A2 => n40013, B1 => n41246, B2 =>
                           n40006, C1 => n718, C2 => n40000, ZN => n7990);
   U32538 : OAI222_X1 port map( A1 => n40868, A2 => n40013, B1 => n41252, B2 =>
                           n40006, C1 => n717, C2 => n40000, ZN => n7989);
   U32539 : OAI222_X1 port map( A1 => n40874, A2 => n40013, B1 => n41258, B2 =>
                           n40006, C1 => n716, C2 => n40000, ZN => n7988);
   U32540 : OAI222_X1 port map( A1 => n40880, A2 => n40013, B1 => n41264, B2 =>
                           n40006, C1 => n715, C2 => n40000, ZN => n7987);
   U32541 : OAI222_X1 port map( A1 => n40886, A2 => n40013, B1 => n41270, B2 =>
                           n40006, C1 => n714, C2 => n40000, ZN => n7986);
   U32542 : OAI222_X1 port map( A1 => n40892, A2 => n40013, B1 => n41276, B2 =>
                           n40006, C1 => n713, C2 => n40000, ZN => n7985);
   U32543 : OAI222_X1 port map( A1 => n40898, A2 => n40013, B1 => n41282, B2 =>
                           n40006, C1 => n712, C2 => n40000, ZN => n7984);
   U32544 : OAI222_X1 port map( A1 => n40904, A2 => n40013, B1 => n41288, B2 =>
                           n40006, C1 => n711, C2 => n40000, ZN => n7983);
   U32545 : OAI222_X1 port map( A1 => n40622, A2 => n40035, B1 => n41006, B2 =>
                           n40028, C1 => n822, C2 => n40022, ZN => n8094);
   U32546 : OAI222_X1 port map( A1 => n40628, A2 => n40035, B1 => n41012, B2 =>
                           n40028, C1 => n821, C2 => n40022, ZN => n8093);
   U32547 : OAI222_X1 port map( A1 => n40634, A2 => n40035, B1 => n41018, B2 =>
                           n40028, C1 => n820, C2 => n40022, ZN => n8092);
   U32548 : OAI222_X1 port map( A1 => n40640, A2 => n40035, B1 => n41024, B2 =>
                           n40028, C1 => n819, C2 => n40022, ZN => n8091);
   U32549 : OAI222_X1 port map( A1 => n40646, A2 => n40035, B1 => n41030, B2 =>
                           n40028, C1 => n818, C2 => n40022, ZN => n8090);
   U32550 : OAI222_X1 port map( A1 => n40652, A2 => n40035, B1 => n41036, B2 =>
                           n40028, C1 => n817, C2 => n40022, ZN => n8089);
   U32551 : OAI222_X1 port map( A1 => n40658, A2 => n40035, B1 => n41042, B2 =>
                           n40028, C1 => n816, C2 => n40022, ZN => n8088);
   U32552 : OAI222_X1 port map( A1 => n40664, A2 => n40035, B1 => n41048, B2 =>
                           n40028, C1 => n815, C2 => n40022, ZN => n8087);
   U32553 : OAI222_X1 port map( A1 => n40670, A2 => n40035, B1 => n41054, B2 =>
                           n40028, C1 => n814, C2 => n40022, ZN => n8086);
   U32554 : OAI222_X1 port map( A1 => n40676, A2 => n40035, B1 => n41060, B2 =>
                           n40028, C1 => n813_port, C2 => n40021, ZN => n8085);
   U32555 : OAI222_X1 port map( A1 => n40682, A2 => n40035, B1 => n41066, B2 =>
                           n40028, C1 => n812_port, C2 => n40021, ZN => n8084);
   U32556 : OAI222_X1 port map( A1 => n40688, A2 => n40035, B1 => n41072, B2 =>
                           n40028, C1 => n811_port, C2 => n40021, ZN => n8083);
   U32557 : OAI222_X1 port map( A1 => n40694, A2 => n40034, B1 => n41078, B2 =>
                           n40027, C1 => n810, C2 => n40021, ZN => n8082);
   U32558 : OAI222_X1 port map( A1 => n40700, A2 => n40034, B1 => n41084, B2 =>
                           n40027, C1 => n809, C2 => n40021, ZN => n8081);
   U32559 : OAI222_X1 port map( A1 => n40706, A2 => n40034, B1 => n41090, B2 =>
                           n40027, C1 => n808, C2 => n40021, ZN => n8080);
   U32560 : OAI222_X1 port map( A1 => n40712, A2 => n40034, B1 => n41096, B2 =>
                           n40027, C1 => n807, C2 => n40021, ZN => n8079);
   U32561 : OAI222_X1 port map( A1 => n40718, A2 => n40034, B1 => n41102, B2 =>
                           n40027, C1 => n806, C2 => n40021, ZN => n8078);
   U32562 : OAI222_X1 port map( A1 => n40724, A2 => n40034, B1 => n41108, B2 =>
                           n40027, C1 => n805, C2 => n40021, ZN => n8077);
   U32563 : OAI222_X1 port map( A1 => n40730, A2 => n40034, B1 => n41114, B2 =>
                           n40027, C1 => n804, C2 => n40021, ZN => n8076);
   U32564 : OAI222_X1 port map( A1 => n40736, A2 => n40034, B1 => n41120, B2 =>
                           n40027, C1 => n803, C2 => n40021, ZN => n8075);
   U32565 : OAI222_X1 port map( A1 => n40742, A2 => n40034, B1 => n41126, B2 =>
                           n40027, C1 => n802, C2 => n40021, ZN => n8074);
   U32566 : OAI222_X1 port map( A1 => n40748, A2 => n40034, B1 => n41132, B2 =>
                           n40027, C1 => n801, C2 => n40021, ZN => n8073);
   U32567 : OAI222_X1 port map( A1 => n40754, A2 => n40034, B1 => n41138, B2 =>
                           n40027, C1 => n800, C2 => n40020, ZN => n8072);
   U32568 : OAI222_X1 port map( A1 => n40760, A2 => n40034, B1 => n41144, B2 =>
                           n40027, C1 => n799, C2 => n40020, ZN => n8071);
   U32569 : OAI222_X1 port map( A1 => n40766, A2 => n40033, B1 => n41150, B2 =>
                           n40026, C1 => n798, C2 => n40020, ZN => n8070);
   U32570 : OAI222_X1 port map( A1 => n40772, A2 => n40033, B1 => n41156, B2 =>
                           n40026, C1 => n797, C2 => n40020, ZN => n8069);
   U32571 : OAI222_X1 port map( A1 => n40778, A2 => n40033, B1 => n41162, B2 =>
                           n40026, C1 => n796, C2 => n40020, ZN => n8068);
   U32572 : OAI222_X1 port map( A1 => n40784, A2 => n40033, B1 => n41168, B2 =>
                           n40026, C1 => n795, C2 => n40020, ZN => n8067);
   U32573 : OAI222_X1 port map( A1 => n40790, A2 => n40033, B1 => n41174, B2 =>
                           n40026, C1 => n794, C2 => n40020, ZN => n8066);
   U32574 : OAI222_X1 port map( A1 => n40796, A2 => n40033, B1 => n41180, B2 =>
                           n40026, C1 => n793, C2 => n40020, ZN => n8065);
   U32575 : OAI222_X1 port map( A1 => n40802, A2 => n40033, B1 => n41186, B2 =>
                           n40026, C1 => n792, C2 => n40020, ZN => n8064);
   U32576 : OAI222_X1 port map( A1 => n40808, A2 => n40033, B1 => n41192, B2 =>
                           n40026, C1 => n791, C2 => n40020, ZN => n8063);
   U32577 : OAI222_X1 port map( A1 => n40814, A2 => n40033, B1 => n41198, B2 =>
                           n40026, C1 => n790, C2 => n40020, ZN => n8062);
   U32578 : OAI222_X1 port map( A1 => n40820, A2 => n40033, B1 => n41204, B2 =>
                           n40026, C1 => n789, C2 => n40020, ZN => n8061);
   U32579 : OAI222_X1 port map( A1 => n40826, A2 => n40033, B1 => n41210, B2 =>
                           n40026, C1 => n788, C2 => n40020, ZN => n8060);
   U32580 : OAI222_X1 port map( A1 => n40832, A2 => n40033, B1 => n41216, B2 =>
                           n40026, C1 => n787, C2 => n40019, ZN => n8059);
   U32581 : OAI222_X1 port map( A1 => n40838, A2 => n40032, B1 => n41222, B2 =>
                           n40025, C1 => n786, C2 => n40019, ZN => n8058);
   U32582 : OAI222_X1 port map( A1 => n40844, A2 => n40032, B1 => n41228, B2 =>
                           n40025, C1 => n785, C2 => n40019, ZN => n8057);
   U32583 : OAI222_X1 port map( A1 => n40850, A2 => n40032, B1 => n41234, B2 =>
                           n40025, C1 => n784, C2 => n40019, ZN => n8056);
   U32584 : OAI222_X1 port map( A1 => n40856, A2 => n40032, B1 => n41240, B2 =>
                           n40025, C1 => n783, C2 => n40019, ZN => n8055);
   U32585 : OAI222_X1 port map( A1 => n40862, A2 => n40032, B1 => n41246, B2 =>
                           n40025, C1 => n782, C2 => n40019, ZN => n8054);
   U32586 : OAI222_X1 port map( A1 => n40868, A2 => n40032, B1 => n41252, B2 =>
                           n40025, C1 => n781, C2 => n40019, ZN => n8053);
   U32587 : OAI222_X1 port map( A1 => n40874, A2 => n40032, B1 => n41258, B2 =>
                           n40025, C1 => n780, C2 => n40019, ZN => n8052);
   U32588 : OAI222_X1 port map( A1 => n40880, A2 => n40032, B1 => n41264, B2 =>
                           n40025, C1 => n779, C2 => n40019, ZN => n8051);
   U32589 : OAI222_X1 port map( A1 => n40886, A2 => n40032, B1 => n41270, B2 =>
                           n40025, C1 => n778, C2 => n40019, ZN => n8050);
   U32590 : OAI222_X1 port map( A1 => n40892, A2 => n40032, B1 => n41276, B2 =>
                           n40025, C1 => n777, C2 => n40019, ZN => n8049);
   U32591 : OAI222_X1 port map( A1 => n40898, A2 => n40032, B1 => n41282, B2 =>
                           n40025, C1 => n776, C2 => n40019, ZN => n8048);
   U32592 : OAI222_X1 port map( A1 => n40904, A2 => n40032, B1 => n41288, B2 =>
                           n40025, C1 => n775, C2 => n40019, ZN => n8047);
   U32593 : OAI222_X1 port map( A1 => n40736, A2 => n39818, B1 => n41120, B2 =>
                           n39811, C1 => n99, C2 => n39805, ZN => n7371);
   U32594 : OAI222_X1 port map( A1 => n40742, A2 => n39818, B1 => n41126, B2 =>
                           n39811, C1 => n98, C2 => n39805, ZN => n7370);
   U32595 : OAI222_X1 port map( A1 => n40748, A2 => n39818, B1 => n41132, B2 =>
                           n39811, C1 => n97, C2 => n39805, ZN => n7369);
   U32596 : OAI222_X1 port map( A1 => n40754, A2 => n39818, B1 => n41138, B2 =>
                           n39811, C1 => n96, C2 => n39804, ZN => n7368);
   U32597 : OAI222_X1 port map( A1 => n40760, A2 => n39818, B1 => n41144, B2 =>
                           n39811, C1 => n95, C2 => n39804, ZN => n7367);
   U32598 : OAI222_X1 port map( A1 => n40766, A2 => n39817, B1 => n41150, B2 =>
                           n39810, C1 => n94, C2 => n39804, ZN => n7366);
   U32599 : OAI222_X1 port map( A1 => n40772, A2 => n39817, B1 => n41156, B2 =>
                           n39810, C1 => n93, C2 => n39804, ZN => n7365);
   U32600 : OAI222_X1 port map( A1 => n40778, A2 => n39817, B1 => n41162, B2 =>
                           n39810, C1 => n92, C2 => n39804, ZN => n7364);
   U32601 : OAI222_X1 port map( A1 => n40784, A2 => n39817, B1 => n41168, B2 =>
                           n39810, C1 => n91, C2 => n39804, ZN => n7363);
   U32602 : OAI222_X1 port map( A1 => n40790, A2 => n39817, B1 => n41174, B2 =>
                           n39810, C1 => n90, C2 => n39804, ZN => n7362);
   U32603 : OAI222_X1 port map( A1 => n40796, A2 => n39817, B1 => n41180, B2 =>
                           n39810, C1 => n89, C2 => n39804, ZN => n7361);
   U32604 : OAI222_X1 port map( A1 => n40802, A2 => n39817, B1 => n41186, B2 =>
                           n39810, C1 => n88, C2 => n39804, ZN => n7360);
   U32605 : OAI222_X1 port map( A1 => n40808, A2 => n39817, B1 => n41192, B2 =>
                           n39810, C1 => n87, C2 => n39804, ZN => n7359);
   U32606 : OAI222_X1 port map( A1 => n40814, A2 => n39817, B1 => n41198, B2 =>
                           n39810, C1 => n86, C2 => n39804, ZN => n7358);
   U32607 : OAI222_X1 port map( A1 => n40820, A2 => n39817, B1 => n41204, B2 =>
                           n39810, C1 => n85, C2 => n39804, ZN => n7357);
   U32608 : OAI222_X1 port map( A1 => n40826, A2 => n39817, B1 => n41210, B2 =>
                           n39810, C1 => n84, C2 => n39804, ZN => n7356);
   U32609 : OAI222_X1 port map( A1 => n40832, A2 => n39817, B1 => n41216, B2 =>
                           n39810, C1 => n83, C2 => n39803, ZN => n7355);
   U32610 : OAI222_X1 port map( A1 => n40838, A2 => n39816, B1 => n41222, B2 =>
                           n39809, C1 => n82, C2 => n39803, ZN => n7354);
   U32611 : OAI222_X1 port map( A1 => n40844, A2 => n39816, B1 => n41228, B2 =>
                           n39809, C1 => n81, C2 => n39803, ZN => n7353);
   U32612 : OAI222_X1 port map( A1 => n40850, A2 => n39816, B1 => n41234, B2 =>
                           n39809, C1 => n80, C2 => n39803, ZN => n7352);
   U32613 : OAI222_X1 port map( A1 => n40856, A2 => n39816, B1 => n41240, B2 =>
                           n39809, C1 => n79, C2 => n39803, ZN => n7351);
   U32614 : OAI222_X1 port map( A1 => n40862, A2 => n39816, B1 => n41246, B2 =>
                           n39809, C1 => n78, C2 => n39803, ZN => n7350);
   U32615 : OAI222_X1 port map( A1 => n40868, A2 => n39816, B1 => n41252, B2 =>
                           n39809, C1 => n77, C2 => n39803, ZN => n7349);
   U32616 : OAI222_X1 port map( A1 => n40874, A2 => n39816, B1 => n41258, B2 =>
                           n39809, C1 => n76, C2 => n39803, ZN => n7348);
   U32617 : OAI222_X1 port map( A1 => n40880, A2 => n39816, B1 => n41264, B2 =>
                           n39809, C1 => n75, C2 => n39803, ZN => n7347);
   U32618 : OAI222_X1 port map( A1 => n40886, A2 => n39816, B1 => n41270, B2 =>
                           n39809, C1 => n74, C2 => n39803, ZN => n7346);
   U32619 : OAI222_X1 port map( A1 => n40892, A2 => n39816, B1 => n41276, B2 =>
                           n39809, C1 => n73, C2 => n39803, ZN => n7345);
   U32620 : OAI222_X1 port map( A1 => n40898, A2 => n39816, B1 => n41282, B2 =>
                           n39809, C1 => n72, C2 => n39803, ZN => n7344);
   U32621 : OAI222_X1 port map( A1 => n40904, A2 => n39816, B1 => n41288, B2 =>
                           n39809, C1 => n71, C2 => n39803, ZN => n7343);
   U32622 : OAI222_X1 port map( A1 => n40910, A2 => n39815, B1 => n41294, B2 =>
                           n39808, C1 => n70, C2 => n39802, ZN => n7342);
   U32623 : OAI222_X1 port map( A1 => n40916, A2 => n39815, B1 => n41300, B2 =>
                           n39808, C1 => n69, C2 => n39802, ZN => n7341);
   U32624 : OAI222_X1 port map( A1 => n40922, A2 => n39815, B1 => n41306, B2 =>
                           n39808, C1 => n68, C2 => n39802, ZN => n7340);
   U32625 : OAI222_X1 port map( A1 => n40928, A2 => n39815, B1 => n41312, B2 =>
                           n39808, C1 => n67, C2 => n39802, ZN => n7339);
   U32626 : OAI222_X1 port map( A1 => n40934, A2 => n39815, B1 => n41318, B2 =>
                           n39808, C1 => n66, C2 => n39802, ZN => n7338);
   U32627 : OAI222_X1 port map( A1 => n40940, A2 => n39815, B1 => n41324, B2 =>
                           n39808, C1 => n65, C2 => n39802, ZN => n7337);
   U32628 : OAI222_X1 port map( A1 => n40946, A2 => n39815, B1 => n41330, B2 =>
                           n39808, C1 => n64, C2 => n39802, ZN => n7336);
   U32629 : OAI222_X1 port map( A1 => n40952, A2 => n39815, B1 => n41336, B2 =>
                           n39808, C1 => n63, C2 => n39802, ZN => n7335);
   U32630 : OAI222_X1 port map( A1 => n40970, A2 => n39815, B1 => n41354, B2 =>
                           n39808, C1 => n60, C2 => n39802, ZN => n7332);
   U32631 : OAI222_X1 port map( A1 => n40976, A2 => n39815, B1 => n41360, B2 =>
                           n39808, C1 => n59, C2 => n39802, ZN => n7331);
   U32632 : OAI222_X1 port map( A1 => n40958, A2 => n39815, B1 => n41342, B2 =>
                           n39808, C1 => n62, C2 => n39802, ZN => n7334);
   U32633 : OAI222_X1 port map( A1 => n40964, A2 => n39815, B1 => n41348, B2 =>
                           n39808, C1 => n61, C2 => n39802, ZN => n7333);
   U32634 : OAI222_X1 port map( A1 => n40598, A2 => n39919, B1 => n40982, B2 =>
                           n39912, C1 => n442, C2 => n39905, ZN => n7714);
   U32635 : OAI222_X1 port map( A1 => n40604, A2 => n39919, B1 => n40988, B2 =>
                           n39912, C1 => n441, C2 => n39905, ZN => n7713);
   U32636 : OAI222_X1 port map( A1 => n40610, A2 => n39919, B1 => n40994, B2 =>
                           n39912, C1 => n440, C2 => n39905, ZN => n7712);
   U32637 : OAI222_X1 port map( A1 => n40616, A2 => n39919, B1 => n41000, B2 =>
                           n39912, C1 => n439, C2 => n39905, ZN => n7711);
   U32638 : OAI222_X1 port map( A1 => n40598, A2 => n39938, B1 => n40982, B2 =>
                           n39931, C1 => n506, C2 => n39924, ZN => n7778);
   U32639 : OAI222_X1 port map( A1 => n40604, A2 => n39938, B1 => n40988, B2 =>
                           n39931, C1 => n505, C2 => n39924, ZN => n7777);
   U32640 : OAI222_X1 port map( A1 => n40610, A2 => n39938, B1 => n40994, B2 =>
                           n39931, C1 => n504, C2 => n39924, ZN => n7776);
   U32641 : OAI222_X1 port map( A1 => n40616, A2 => n39938, B1 => n41000, B2 =>
                           n39931, C1 => n503, C2 => n39924, ZN => n7775);
   U32642 : OAI222_X1 port map( A1 => n40598, A2 => n40017, B1 => n40982, B2 =>
                           n40010, C1 => n762, C2 => n40003, ZN => n8034);
   U32643 : OAI222_X1 port map( A1 => n40604, A2 => n40017, B1 => n40988, B2 =>
                           n40010, C1 => n761, C2 => n40003, ZN => n8033);
   U32644 : OAI222_X1 port map( A1 => n40610, A2 => n40017, B1 => n40994, B2 =>
                           n40010, C1 => n760, C2 => n40003, ZN => n8032);
   U32645 : OAI222_X1 port map( A1 => n40616, A2 => n40017, B1 => n41000, B2 =>
                           n40010, C1 => n759, C2 => n40003, ZN => n8031);
   U32646 : OAI222_X1 port map( A1 => n40598, A2 => n40036, B1 => n40982, B2 =>
                           n40029, C1 => n826, C2 => n40022, ZN => n8098);
   U32647 : OAI222_X1 port map( A1 => n40604, A2 => n40036, B1 => n40988, B2 =>
                           n40029, C1 => n825, C2 => n40022, ZN => n8097);
   U32648 : OAI222_X1 port map( A1 => n40610, A2 => n40036, B1 => n40994, B2 =>
                           n40029, C1 => n824, C2 => n40022, ZN => n8096);
   U32649 : OAI222_X1 port map( A1 => n40616, A2 => n40036, B1 => n41000, B2 =>
                           n40029, C1 => n823, C2 => n40022, ZN => n8095);
   U32650 : OAI222_X1 port map( A1 => n40659, A2 => n40134, B1 => n41043, B2 =>
                           n40127, C1 => n25458, C2 => n40117, ZN => n8408);
   U32651 : OAI222_X1 port map( A1 => n40665, A2 => n40134, B1 => n41049, B2 =>
                           n40127, C1 => n25459, C2 => n40117, ZN => n8407);
   U32652 : OAI222_X1 port map( A1 => n40671, A2 => n40134, B1 => n41055, B2 =>
                           n40127, C1 => n25460, C2 => n40117, ZN => n8406);
   U32653 : OAI222_X1 port map( A1 => n40677, A2 => n40134, B1 => n41061, B2 =>
                           n40127, C1 => n25461, C2 => n40117, ZN => n8405);
   U32654 : OAI222_X1 port map( A1 => n40683, A2 => n40134, B1 => n41067, B2 =>
                           n40127, C1 => n25462, C2 => n40117, ZN => n8404);
   U32655 : OAI222_X1 port map( A1 => n40689, A2 => n40134, B1 => n41073, B2 =>
                           n40127, C1 => n25463, C2 => n40118, ZN => n8403);
   U32656 : OAI222_X1 port map( A1 => n40695, A2 => n40133, B1 => n41079, B2 =>
                           n40126, C1 => n25464, C2 => n40117, ZN => n8402);
   U32657 : OAI222_X1 port map( A1 => n40701, A2 => n40133, B1 => n41085, B2 =>
                           n40126, C1 => n25465, C2 => n40117, ZN => n8401);
   U32658 : OAI222_X1 port map( A1 => n40707, A2 => n40133, B1 => n41091, B2 =>
                           n40126, C1 => n25466, C2 => n40117, ZN => n8400);
   U32659 : OAI222_X1 port map( A1 => n40713, A2 => n40133, B1 => n41097, B2 =>
                           n40126, C1 => n25467, C2 => n40117, ZN => n8399);
   U32660 : OAI222_X1 port map( A1 => n40719, A2 => n40133, B1 => n41103, B2 =>
                           n40126, C1 => n25468, C2 => n40117, ZN => n8398);
   U32661 : OAI222_X1 port map( A1 => n40725, A2 => n40133, B1 => n41109, B2 =>
                           n40126, C1 => n25469, C2 => n40117, ZN => n8397);
   U32662 : OAI222_X1 port map( A1 => n40731, A2 => n40133, B1 => n41115, B2 =>
                           n40126, C1 => n25470, C2 => n40117, ZN => n8396);
   U32663 : OAI222_X1 port map( A1 => n40737, A2 => n40133, B1 => n41121, B2 =>
                           n40126, C1 => n25471, C2 => n40117, ZN => n8395);
   U32664 : OAI222_X1 port map( A1 => n40743, A2 => n40133, B1 => n41127, B2 =>
                           n40126, C1 => n25472, C2 => n40118, ZN => n8394);
   U32665 : OAI222_X1 port map( A1 => n40749, A2 => n40133, B1 => n41133, B2 =>
                           n40126, C1 => n25473, C2 => n40118, ZN => n8393);
   U32666 : OAI222_X1 port map( A1 => n40755, A2 => n40133, B1 => n41139, B2 =>
                           n40126, C1 => n25474, C2 => n40118, ZN => n8392);
   U32667 : OAI222_X1 port map( A1 => n40761, A2 => n40133, B1 => n41145, B2 =>
                           n40126, C1 => n25475, C2 => n40118, ZN => n8391);
   U32668 : OAI222_X1 port map( A1 => n40767, A2 => n40132, B1 => n41151, B2 =>
                           n40125, C1 => n25476, C2 => n40118, ZN => n8390);
   U32669 : OAI222_X1 port map( A1 => n40773, A2 => n40132, B1 => n41157, B2 =>
                           n40125, C1 => n25477, C2 => n40118, ZN => n8389);
   U32670 : OAI222_X1 port map( A1 => n40779, A2 => n40132, B1 => n41163, B2 =>
                           n40125, C1 => n25478, C2 => n40118, ZN => n8388);
   U32671 : OAI222_X1 port map( A1 => n40785, A2 => n40132, B1 => n41169, B2 =>
                           n40125, C1 => n25479, C2 => n40118, ZN => n8387);
   U32672 : OAI222_X1 port map( A1 => n40791, A2 => n40132, B1 => n41175, B2 =>
                           n40125, C1 => n25480, C2 => n40118, ZN => n8386);
   U32673 : OAI222_X1 port map( A1 => n40797, A2 => n40132, B1 => n41181, B2 =>
                           n40125, C1 => n25481, C2 => n40118, ZN => n8385);
   U32674 : OAI222_X1 port map( A1 => n40803, A2 => n40132, B1 => n41187, B2 =>
                           n40125, C1 => n25482, C2 => n40118, ZN => n8384);
   U32675 : OAI222_X1 port map( A1 => n40809, A2 => n40132, B1 => n41193, B2 =>
                           n40125, C1 => n25483, C2 => n40118, ZN => n8383);
   U32676 : OAI222_X1 port map( A1 => n40815, A2 => n40132, B1 => n41199, B2 =>
                           n40125, C1 => n25484, C2 => n40119, ZN => n8382);
   U32677 : OAI222_X1 port map( A1 => n40821, A2 => n40132, B1 => n41205, B2 =>
                           n40125, C1 => n25485, C2 => n40119, ZN => n8381);
   U32678 : OAI222_X1 port map( A1 => n40827, A2 => n40132, B1 => n41211, B2 =>
                           n40125, C1 => n25486, C2 => n40119, ZN => n8380);
   U32679 : OAI222_X1 port map( A1 => n40833, A2 => n40132, B1 => n41217, B2 =>
                           n40125, C1 => n25487, C2 => n40119, ZN => n8379);
   U32680 : OAI222_X1 port map( A1 => n40839, A2 => n40131, B1 => n41223, B2 =>
                           n40124, C1 => n25488, C2 => n40119, ZN => n8378);
   U32681 : OAI222_X1 port map( A1 => n40845, A2 => n40131, B1 => n41229, B2 =>
                           n40124, C1 => n25489, C2 => n40119, ZN => n8377);
   U32682 : OAI222_X1 port map( A1 => n40851, A2 => n40131, B1 => n41235, B2 =>
                           n40124, C1 => n25490, C2 => n40119, ZN => n8376);
   U32683 : OAI222_X1 port map( A1 => n40857, A2 => n40131, B1 => n41241, B2 =>
                           n40124, C1 => n25491, C2 => n40119, ZN => n8375);
   U32684 : OAI222_X1 port map( A1 => n40863, A2 => n40131, B1 => n41247, B2 =>
                           n40124, C1 => n25492, C2 => n40119, ZN => n8374);
   U32685 : OAI222_X1 port map( A1 => n40869, A2 => n40131, B1 => n41253, B2 =>
                           n40124, C1 => n25493, C2 => n40119, ZN => n8373);
   U32686 : OAI222_X1 port map( A1 => n40875, A2 => n40131, B1 => n41259, B2 =>
                           n40124, C1 => n25494, C2 => n40119, ZN => n8372);
   U32687 : OAI222_X1 port map( A1 => n40881, A2 => n40131, B1 => n41265, B2 =>
                           n40124, C1 => n25495, C2 => n40119, ZN => n8371);
   U32688 : OAI222_X1 port map( A1 => n40887, A2 => n40131, B1 => n41271, B2 =>
                           n40124, C1 => n25496, C2 => n40119, ZN => n8370);
   U32689 : OAI222_X1 port map( A1 => n40893, A2 => n40131, B1 => n41277, B2 =>
                           n40124, C1 => n25497, C2 => n40120, ZN => n8369);
   U32690 : OAI222_X1 port map( A1 => n40899, A2 => n40131, B1 => n41283, B2 =>
                           n40124, C1 => n25498, C2 => n40120, ZN => n8368);
   U32691 : OAI222_X1 port map( A1 => n40905, A2 => n40131, B1 => n41289, B2 =>
                           n40124, C1 => n25499, C2 => n40120, ZN => n8367);
   U32692 : OAI222_X1 port map( A1 => n40911, A2 => n40130, B1 => n41295, B2 =>
                           n40123, C1 => n25500, C2 => n40120, ZN => n8366);
   U32693 : OAI222_X1 port map( A1 => n40917, A2 => n40130, B1 => n41301, B2 =>
                           n40123, C1 => n25501, C2 => n40120, ZN => n8365);
   U32694 : OAI222_X1 port map( A1 => n40923, A2 => n40130, B1 => n41307, B2 =>
                           n40123, C1 => n25502, C2 => n40120, ZN => n8364);
   U32695 : OAI222_X1 port map( A1 => n40929, A2 => n40130, B1 => n41313, B2 =>
                           n40123, C1 => n25503, C2 => n40120, ZN => n8363);
   U32696 : OAI222_X1 port map( A1 => n40935, A2 => n40130, B1 => n41319, B2 =>
                           n40123, C1 => n25504, C2 => n40120, ZN => n8362);
   U32697 : OAI222_X1 port map( A1 => n40941, A2 => n40130, B1 => n41325, B2 =>
                           n40123, C1 => n25505, C2 => n40120, ZN => n8361);
   U32698 : OAI222_X1 port map( A1 => n40947, A2 => n40130, B1 => n41331, B2 =>
                           n40123, C1 => n25506, C2 => n40120, ZN => n8360);
   U32699 : OAI222_X1 port map( A1 => n40953, A2 => n40130, B1 => n41337, B2 =>
                           n40123, C1 => n25507, C2 => n40120, ZN => n8359);
   U32700 : OAI222_X1 port map( A1 => n40959, A2 => n40130, B1 => n41343, B2 =>
                           n40123, C1 => n25508, C2 => n40120, ZN => n8358);
   U32701 : OAI222_X1 port map( A1 => n40965, A2 => n40130, B1 => n41349, B2 =>
                           n40123, C1 => n25509, C2 => n40121, ZN => n8357);
   U32702 : OAI222_X1 port map( A1 => n40971, A2 => n40130, B1 => n41355, B2 =>
                           n40123, C1 => n25510, C2 => n40120, ZN => n8356);
   U32703 : OAI222_X1 port map( A1 => n40977, A2 => n40130, B1 => n41361, B2 =>
                           n40123, C1 => n25511, C2 => n40116, ZN => n8355);
   U32704 : OAI222_X1 port map( A1 => n40599, A2 => n40115, B1 => n40983, B2 =>
                           n40108, C1 => n25398, C2 => n40101, ZN => n8354);
   U32705 : OAI222_X1 port map( A1 => n40605, A2 => n40115, B1 => n40989, B2 =>
                           n40108, C1 => n25399, C2 => n40101, ZN => n8353);
   U32706 : OAI222_X1 port map( A1 => n40611, A2 => n40115, B1 => n40995, B2 =>
                           n40108, C1 => n25400, C2 => n40101, ZN => n8352);
   U32707 : OAI222_X1 port map( A1 => n40617, A2 => n40115, B1 => n41001, B2 =>
                           n40108, C1 => n25401, C2 => n40101, ZN => n8351);
   U32708 : OAI222_X1 port map( A1 => n40623, A2 => n40114, B1 => n41007, B2 =>
                           n40107, C1 => n25402, C2 => n40101, ZN => n8350);
   U32709 : OAI222_X1 port map( A1 => n40629, A2 => n40114, B1 => n41013, B2 =>
                           n40107, C1 => n25403, C2 => n40101, ZN => n8349);
   U32710 : OAI222_X1 port map( A1 => n40635, A2 => n40114, B1 => n41019, B2 =>
                           n40107, C1 => n25404, C2 => n40101, ZN => n8348);
   U32711 : OAI222_X1 port map( A1 => n40641, A2 => n40114, B1 => n41025, B2 =>
                           n40107, C1 => n25405, C2 => n40101, ZN => n8347);
   U32712 : OAI222_X1 port map( A1 => n40647, A2 => n40114, B1 => n41031, B2 =>
                           n40107, C1 => n25406, C2 => n40101, ZN => n8346);
   U32713 : OAI222_X1 port map( A1 => n40653, A2 => n40114, B1 => n41037, B2 =>
                           n40107, C1 => n25407, C2 => n40101, ZN => n8345);
   U32714 : OAI222_X1 port map( A1 => n40659, A2 => n40114, B1 => n41043, B2 =>
                           n40107, C1 => n25408, C2 => n40101, ZN => n8344);
   U32715 : OAI222_X1 port map( A1 => n40665, A2 => n40114, B1 => n41049, B2 =>
                           n40107, C1 => n25409, C2 => n40101, ZN => n8343);
   U32716 : OAI222_X1 port map( A1 => n40671, A2 => n40114, B1 => n41055, B2 =>
                           n40107, C1 => n25410, C2 => n40101, ZN => n8342);
   U32717 : OAI222_X1 port map( A1 => n40677, A2 => n40114, B1 => n41061, B2 =>
                           n40107, C1 => n25411, C2 => n40100, ZN => n8341);
   U32718 : OAI222_X1 port map( A1 => n40683, A2 => n40114, B1 => n41067, B2 =>
                           n40107, C1 => n25412, C2 => n40100, ZN => n8340);
   U32719 : OAI222_X1 port map( A1 => n40689, A2 => n40114, B1 => n41073, B2 =>
                           n40107, C1 => n25413, C2 => n40100, ZN => n8339);
   U32720 : OAI222_X1 port map( A1 => n40695, A2 => n40113, B1 => n41079, B2 =>
                           n40106, C1 => n25414, C2 => n40100, ZN => n8338);
   U32721 : OAI222_X1 port map( A1 => n40701, A2 => n40113, B1 => n41085, B2 =>
                           n40106, C1 => n25415, C2 => n40100, ZN => n8337);
   U32722 : OAI222_X1 port map( A1 => n40707, A2 => n40113, B1 => n41091, B2 =>
                           n40106, C1 => n25416, C2 => n40100, ZN => n8336);
   U32723 : OAI222_X1 port map( A1 => n40713, A2 => n40113, B1 => n41097, B2 =>
                           n40106, C1 => n25417, C2 => n40100, ZN => n8335);
   U32724 : OAI222_X1 port map( A1 => n40719, A2 => n40113, B1 => n41103, B2 =>
                           n40106, C1 => n25418, C2 => n40100, ZN => n8334);
   U32725 : OAI222_X1 port map( A1 => n40725, A2 => n40113, B1 => n41109, B2 =>
                           n40106, C1 => n25419, C2 => n40100, ZN => n8333);
   U32726 : OAI222_X1 port map( A1 => n40731, A2 => n40113, B1 => n41115, B2 =>
                           n40106, C1 => n25420, C2 => n40100, ZN => n8332);
   U32727 : OAI222_X1 port map( A1 => n40737, A2 => n40113, B1 => n41121, B2 =>
                           n40106, C1 => n25421, C2 => n40100, ZN => n8331);
   U32728 : OAI222_X1 port map( A1 => n40743, A2 => n40113, B1 => n41127, B2 =>
                           n40106, C1 => n25422, C2 => n40100, ZN => n8330);
   U32729 : OAI222_X1 port map( A1 => n40749, A2 => n40113, B1 => n41133, B2 =>
                           n40106, C1 => n25423, C2 => n40100, ZN => n8329);
   U32730 : OAI222_X1 port map( A1 => n40755, A2 => n40113, B1 => n41139, B2 =>
                           n40106, C1 => n25424, C2 => n40099, ZN => n8328);
   U32731 : OAI222_X1 port map( A1 => n40761, A2 => n40113, B1 => n41145, B2 =>
                           n40106, C1 => n25425, C2 => n40099, ZN => n8327);
   U32732 : OAI222_X1 port map( A1 => n40767, A2 => n40112, B1 => n41151, B2 =>
                           n40105, C1 => n25426, C2 => n40099, ZN => n8326);
   U32733 : OAI222_X1 port map( A1 => n40773, A2 => n40112, B1 => n41157, B2 =>
                           n40105, C1 => n25427, C2 => n40099, ZN => n8325);
   U32734 : OAI222_X1 port map( A1 => n40779, A2 => n40112, B1 => n41163, B2 =>
                           n40105, C1 => n25428, C2 => n40099, ZN => n8324);
   U32735 : OAI222_X1 port map( A1 => n40785, A2 => n40112, B1 => n41169, B2 =>
                           n40105, C1 => n25429, C2 => n40099, ZN => n8323);
   U32736 : OAI222_X1 port map( A1 => n40791, A2 => n40112, B1 => n41175, B2 =>
                           n40105, C1 => n25430, C2 => n40099, ZN => n8322);
   U32737 : OAI222_X1 port map( A1 => n40797, A2 => n40112, B1 => n41181, B2 =>
                           n40105, C1 => n25431, C2 => n40099, ZN => n8321);
   U32738 : OAI222_X1 port map( A1 => n40803, A2 => n40112, B1 => n41187, B2 =>
                           n40105, C1 => n25432, C2 => n40099, ZN => n8320);
   U32739 : OAI222_X1 port map( A1 => n40809, A2 => n40112, B1 => n41193, B2 =>
                           n40105, C1 => n25433, C2 => n40099, ZN => n8319);
   U32740 : OAI222_X1 port map( A1 => n40815, A2 => n40112, B1 => n41199, B2 =>
                           n40105, C1 => n25434, C2 => n40099, ZN => n8318);
   U32741 : OAI222_X1 port map( A1 => n40821, A2 => n40112, B1 => n41205, B2 =>
                           n40105, C1 => n25435, C2 => n40099, ZN => n8317);
   U32742 : OAI222_X1 port map( A1 => n40827, A2 => n40112, B1 => n41211, B2 =>
                           n40105, C1 => n25436, C2 => n40099, ZN => n8316);
   U32743 : OAI222_X1 port map( A1 => n40833, A2 => n40112, B1 => n41217, B2 =>
                           n40105, C1 => n25437, C2 => n40098, ZN => n8315);
   U32744 : OAI222_X1 port map( A1 => n40839, A2 => n40111, B1 => n41223, B2 =>
                           n40104, C1 => n25438, C2 => n40098, ZN => n8314);
   U32745 : OAI222_X1 port map( A1 => n40845, A2 => n40111, B1 => n41229, B2 =>
                           n40104, C1 => n25439, C2 => n40098, ZN => n8313);
   U32746 : OAI222_X1 port map( A1 => n40851, A2 => n40111, B1 => n41235, B2 =>
                           n40104, C1 => n25440, C2 => n40098, ZN => n8312);
   U32747 : OAI222_X1 port map( A1 => n40857, A2 => n40111, B1 => n41241, B2 =>
                           n40104, C1 => n25441, C2 => n40098, ZN => n8311);
   U32748 : OAI222_X1 port map( A1 => n40863, A2 => n40111, B1 => n41247, B2 =>
                           n40104, C1 => n25442, C2 => n40098, ZN => n8310);
   U32749 : OAI222_X1 port map( A1 => n40869, A2 => n40111, B1 => n41253, B2 =>
                           n40104, C1 => n25443, C2 => n40098, ZN => n8309);
   U32750 : OAI222_X1 port map( A1 => n40875, A2 => n40111, B1 => n41259, B2 =>
                           n40104, C1 => n25444, C2 => n40098, ZN => n8308);
   U32751 : OAI222_X1 port map( A1 => n40881, A2 => n40111, B1 => n41265, B2 =>
                           n40104, C1 => n25445, C2 => n40098, ZN => n8307);
   U32752 : OAI222_X1 port map( A1 => n40887, A2 => n40111, B1 => n41271, B2 =>
                           n40104, C1 => n25446, C2 => n40098, ZN => n8306);
   U32753 : OAI222_X1 port map( A1 => n40893, A2 => n40111, B1 => n41277, B2 =>
                           n40104, C1 => n25447, C2 => n40098, ZN => n8305);
   U32754 : OAI222_X1 port map( A1 => n40899, A2 => n40111, B1 => n41283, B2 =>
                           n40104, C1 => n25448, C2 => n40098, ZN => n8304);
   U32755 : OAI222_X1 port map( A1 => n40905, A2 => n40111, B1 => n41289, B2 =>
                           n40104, C1 => n25449, C2 => n40098, ZN => n8303);
   U32756 : OAI222_X1 port map( A1 => n40911, A2 => n40110, B1 => n41295, B2 =>
                           n40103, C1 => n25450, C2 => n40097, ZN => n8302);
   U32757 : OAI222_X1 port map( A1 => n40917, A2 => n40110, B1 => n41301, B2 =>
                           n40103, C1 => n25451, C2 => n40097, ZN => n8301);
   U32758 : OAI222_X1 port map( A1 => n40923, A2 => n40110, B1 => n41307, B2 =>
                           n40103, C1 => n25452, C2 => n40097, ZN => n8300);
   U32759 : OAI222_X1 port map( A1 => n40929, A2 => n40110, B1 => n41313, B2 =>
                           n40103, C1 => n25453, C2 => n40097, ZN => n8299);
   U32760 : OAI222_X1 port map( A1 => n40935, A2 => n40110, B1 => n41319, B2 =>
                           n40103, C1 => n25454, C2 => n40097, ZN => n8298);
   U32761 : OAI222_X1 port map( A1 => n40941, A2 => n40110, B1 => n41325, B2 =>
                           n40103, C1 => n25455, C2 => n40097, ZN => n8297);
   U32762 : OAI222_X1 port map( A1 => n40947, A2 => n40110, B1 => n41331, B2 =>
                           n40103, C1 => n25456, C2 => n40097, ZN => n8296);
   U32763 : OAI222_X1 port map( A1 => n40953, A2 => n40110, B1 => n41337, B2 =>
                           n40103, C1 => n28840, C2 => n40097, ZN => n8295);
   U32764 : OAI222_X1 port map( A1 => n40959, A2 => n40110, B1 => n41343, B2 =>
                           n40103, C1 => n25457, C2 => n40097, ZN => n8294);
   U32765 : OAI222_X1 port map( A1 => n40965, A2 => n40110, B1 => n41349, B2 =>
                           n40103, C1 => n25395, C2 => n40097, ZN => n8293);
   U32766 : OAI222_X1 port map( A1 => n40971, A2 => n40110, B1 => n41355, B2 =>
                           n40103, C1 => n25396, C2 => n40097, ZN => n8292);
   U32767 : OAI222_X1 port map( A1 => n40977, A2 => n40110, B1 => n41361, B2 =>
                           n40103, C1 => n25397, C2 => n40097, ZN => n8291);
   U32768 : OAI222_X1 port map( A1 => n40598, A2 => n39820, B1 => n40982, B2 =>
                           n39813, C1 => n27943, C2 => n39806, ZN => n7394);
   U32769 : OAI222_X1 port map( A1 => n40604, A2 => n39820, B1 => n40988, B2 =>
                           n39813, C1 => n27942, C2 => n39806, ZN => n7393);
   U32770 : OAI222_X1 port map( A1 => n40610, A2 => n39820, B1 => n40994, B2 =>
                           n39813, C1 => n27941, C2 => n39806, ZN => n7392);
   U32771 : OAI222_X1 port map( A1 => n40616, A2 => n39820, B1 => n41000, B2 =>
                           n39813, C1 => n27940, C2 => n39806, ZN => n7391);
   U32772 : OAI222_X1 port map( A1 => n40622, A2 => n39819, B1 => n41006, B2 =>
                           n39812, C1 => n27939, C2 => n39806, ZN => n7390);
   U32773 : OAI222_X1 port map( A1 => n40628, A2 => n39819, B1 => n41012, B2 =>
                           n39812, C1 => n27938, C2 => n39806, ZN => n7389);
   U32774 : OAI222_X1 port map( A1 => n40634, A2 => n39819, B1 => n41018, B2 =>
                           n39812, C1 => n27937, C2 => n39806, ZN => n7388);
   U32775 : OAI222_X1 port map( A1 => n40640, A2 => n39819, B1 => n41024, B2 =>
                           n39812, C1 => n27936, C2 => n39806, ZN => n7387);
   U32776 : OAI222_X1 port map( A1 => n40646, A2 => n39819, B1 => n41030, B2 =>
                           n39812, C1 => n27935, C2 => n39806, ZN => n7386);
   U32777 : OAI222_X1 port map( A1 => n40652, A2 => n39819, B1 => n41036, B2 =>
                           n39812, C1 => n27934, C2 => n39806, ZN => n7385);
   U32778 : OAI222_X1 port map( A1 => n40658, A2 => n39819, B1 => n41042, B2 =>
                           n39812, C1 => n27933, C2 => n39806, ZN => n7384);
   U32779 : OAI222_X1 port map( A1 => n40664, A2 => n39819, B1 => n41048, B2 =>
                           n39812, C1 => n27932, C2 => n39806, ZN => n7383);
   U32780 : OAI222_X1 port map( A1 => n40670, A2 => n39819, B1 => n41054, B2 =>
                           n39812, C1 => n27931, C2 => n39806, ZN => n7382);
   U32781 : OAI222_X1 port map( A1 => n40676, A2 => n39819, B1 => n41060, B2 =>
                           n39812, C1 => n27930, C2 => n39805, ZN => n7381);
   U32782 : OAI222_X1 port map( A1 => n40682, A2 => n39819, B1 => n41066, B2 =>
                           n39812, C1 => n27929, C2 => n39805, ZN => n7380);
   U32783 : OAI222_X1 port map( A1 => n40688, A2 => n39819, B1 => n41072, B2 =>
                           n39812, C1 => n27928, C2 => n39805, ZN => n7379);
   U32784 : OAI222_X1 port map( A1 => n40694, A2 => n39818, B1 => n41078, B2 =>
                           n39811, C1 => n27927, C2 => n39805, ZN => n7378);
   U32785 : OAI222_X1 port map( A1 => n40700, A2 => n39818, B1 => n41084, B2 =>
                           n39811, C1 => n27926, C2 => n39805, ZN => n7377);
   U32786 : OAI222_X1 port map( A1 => n40706, A2 => n39818, B1 => n41090, B2 =>
                           n39811, C1 => n27925, C2 => n39805, ZN => n7376);
   U32787 : OAI222_X1 port map( A1 => n40712, A2 => n39818, B1 => n41096, B2 =>
                           n39811, C1 => n27924, C2 => n39805, ZN => n7375);
   U32788 : OAI222_X1 port map( A1 => n40718, A2 => n39818, B1 => n41102, B2 =>
                           n39811, C1 => n27923, C2 => n39805, ZN => n7374);
   U32789 : OAI222_X1 port map( A1 => n40724, A2 => n39818, B1 => n41108, B2 =>
                           n39811, C1 => n27922, C2 => n39805, ZN => n7373);
   U32790 : OAI222_X1 port map( A1 => n40730, A2 => n39818, B1 => n41114, B2 =>
                           n39811, C1 => n27921, C2 => n39805, ZN => n7372);
   U32791 : OAI222_X1 port map( A1 => n40912, A2 => n40430, B1 => n41296, B2 =>
                           n40423, C1 => n40420, C2 => n38794, ZN => n9326);
   U32792 : OAI222_X1 port map( A1 => n40918, A2 => n40430, B1 => n41302, B2 =>
                           n40423, C1 => n40420, C2 => n38795, ZN => n9325);
   U32793 : OAI222_X1 port map( A1 => n40924, A2 => n40430, B1 => n41308, B2 =>
                           n40423, C1 => n40420, C2 => n38796, ZN => n9324);
   U32794 : OAI222_X1 port map( A1 => n40930, A2 => n40430, B1 => n41314, B2 =>
                           n40423, C1 => n40420, C2 => n38797, ZN => n9323);
   U32795 : OAI222_X1 port map( A1 => n40936, A2 => n40430, B1 => n41320, B2 =>
                           n40423, C1 => n40420, C2 => n38798, ZN => n9322);
   U32796 : OAI222_X1 port map( A1 => n40942, A2 => n40430, B1 => n41326, B2 =>
                           n40423, C1 => n40420, C2 => n38799, ZN => n9321);
   U32797 : OAI222_X1 port map( A1 => n40948, A2 => n40430, B1 => n41332, B2 =>
                           n40423, C1 => n40420, C2 => n38800, ZN => n9320);
   U32798 : OAI222_X1 port map( A1 => n40960, A2 => n40430, B1 => n41344, B2 =>
                           n40423, C1 => n40420, C2 => n38801, ZN => n9318);
   U32799 : OAI222_X1 port map( A1 => n40624, A2 => n40434, B1 => n41008, B2 =>
                           n40427, C1 => n40416, C2 => n38802, ZN => n9374);
   U32800 : OAI222_X1 port map( A1 => n40630, A2 => n40434, B1 => n41014, B2 =>
                           n40427, C1 => n40416, C2 => n38803, ZN => n9373);
   U32801 : OAI222_X1 port map( A1 => n40636, A2 => n40434, B1 => n41020, B2 =>
                           n40427, C1 => n40416, C2 => n38804, ZN => n9372);
   U32802 : OAI222_X1 port map( A1 => n40642, A2 => n40434, B1 => n41026, B2 =>
                           n40427, C1 => n40416, C2 => n38805, ZN => n9371);
   U32803 : OAI222_X1 port map( A1 => n40648, A2 => n40434, B1 => n41032, B2 =>
                           n40427, C1 => n40416, C2 => n38806, ZN => n9370);
   U32804 : OAI222_X1 port map( A1 => n40654, A2 => n40434, B1 => n41038, B2 =>
                           n40427, C1 => n40416, C2 => n38807, ZN => n9369);
   U32805 : OAI222_X1 port map( A1 => n40660, A2 => n40434, B1 => n41044, B2 =>
                           n40427, C1 => n40416, C2 => n38808, ZN => n9368);
   U32806 : OAI222_X1 port map( A1 => n40666, A2 => n40434, B1 => n41050, B2 =>
                           n40427, C1 => n40416, C2 => n38809, ZN => n9367);
   U32807 : OAI222_X1 port map( A1 => n40672, A2 => n40434, B1 => n41056, B2 =>
                           n40427, C1 => n40417, C2 => n38810, ZN => n9366);
   U32808 : OAI222_X1 port map( A1 => n40678, A2 => n40434, B1 => n41062, B2 =>
                           n40427, C1 => n40417, C2 => n38811, ZN => n9365);
   U32809 : OAI222_X1 port map( A1 => n40684, A2 => n40434, B1 => n41068, B2 =>
                           n40427, C1 => n40417, C2 => n38812, ZN => n9364);
   U32810 : OAI222_X1 port map( A1 => n40690, A2 => n40434, B1 => n41074, B2 =>
                           n40427, C1 => n40418, C2 => n38813, ZN => n9363);
   U32811 : OAI222_X1 port map( A1 => n40696, A2 => n40433, B1 => n41080, B2 =>
                           n40426, C1 => n40417, C2 => n38814, ZN => n9362);
   U32812 : OAI222_X1 port map( A1 => n40702, A2 => n40433, B1 => n41086, B2 =>
                           n40426, C1 => n40417, C2 => n38815, ZN => n9361);
   U32813 : OAI222_X1 port map( A1 => n40708, A2 => n40433, B1 => n41092, B2 =>
                           n40426, C1 => n40417, C2 => n38816, ZN => n9360);
   U32814 : OAI222_X1 port map( A1 => n40714, A2 => n40433, B1 => n41098, B2 =>
                           n40426, C1 => n40417, C2 => n38817, ZN => n9359);
   U32815 : OAI222_X1 port map( A1 => n40720, A2 => n40433, B1 => n41104, B2 =>
                           n40426, C1 => n40417, C2 => n38818, ZN => n9358);
   U32816 : OAI222_X1 port map( A1 => n40726, A2 => n40433, B1 => n41110, B2 =>
                           n40426, C1 => n40417, C2 => n38819, ZN => n9357);
   U32817 : OAI222_X1 port map( A1 => n40732, A2 => n40433, B1 => n41116, B2 =>
                           n40426, C1 => n40417, C2 => n38820, ZN => n9356);
   U32818 : OAI222_X1 port map( A1 => n40738, A2 => n40433, B1 => n41122, B2 =>
                           n40426, C1 => n40417, C2 => n38821, ZN => n9355);
   U32819 : OAI222_X1 port map( A1 => n40744, A2 => n40433, B1 => n41128, B2 =>
                           n40426, C1 => n40417, C2 => n38822, ZN => n9354);
   U32820 : OAI222_X1 port map( A1 => n40750, A2 => n40433, B1 => n41134, B2 =>
                           n40426, C1 => n40418, C2 => n38823, ZN => n9353);
   U32821 : OAI222_X1 port map( A1 => n40756, A2 => n40433, B1 => n41140, B2 =>
                           n40426, C1 => n40418, C2 => n38824, ZN => n9352);
   U32822 : OAI222_X1 port map( A1 => n40762, A2 => n40433, B1 => n41146, B2 =>
                           n40426, C1 => n40418, C2 => n38825, ZN => n9351);
   U32823 : OAI222_X1 port map( A1 => n40768, A2 => n40432, B1 => n41152, B2 =>
                           n40425, C1 => n40418, C2 => n38826, ZN => n9350);
   U32824 : OAI222_X1 port map( A1 => n40774, A2 => n40432, B1 => n41158, B2 =>
                           n40425, C1 => n40418, C2 => n38827, ZN => n9349);
   U32825 : OAI222_X1 port map( A1 => n40780, A2 => n40432, B1 => n41164, B2 =>
                           n40425, C1 => n40418, C2 => n38828, ZN => n9348);
   U32826 : OAI222_X1 port map( A1 => n40786, A2 => n40432, B1 => n41170, B2 =>
                           n40425, C1 => n40418, C2 => n38829, ZN => n9347);
   U32827 : OAI222_X1 port map( A1 => n40792, A2 => n40432, B1 => n41176, B2 =>
                           n40425, C1 => n40418, C2 => n38830, ZN => n9346);
   U32828 : OAI222_X1 port map( A1 => n40798, A2 => n40432, B1 => n41182, B2 =>
                           n40425, C1 => n40418, C2 => n38831, ZN => n9345);
   U32829 : OAI222_X1 port map( A1 => n40804, A2 => n40432, B1 => n41188, B2 =>
                           n40425, C1 => n40418, C2 => n38832, ZN => n9344);
   U32830 : OAI222_X1 port map( A1 => n40810, A2 => n40432, B1 => n41194, B2 =>
                           n40425, C1 => n40418, C2 => n38833, ZN => n9343);
   U32831 : OAI222_X1 port map( A1 => n40816, A2 => n40432, B1 => n41200, B2 =>
                           n40425, C1 => n40419, C2 => n38834, ZN => n9342);
   U32832 : OAI222_X1 port map( A1 => n40822, A2 => n40432, B1 => n41206, B2 =>
                           n40425, C1 => n40419, C2 => n38835, ZN => n9341);
   U32833 : OAI222_X1 port map( A1 => n40828, A2 => n40432, B1 => n41212, B2 =>
                           n40425, C1 => n40419, C2 => n38836, ZN => n9340);
   U32834 : OAI222_X1 port map( A1 => n40834, A2 => n40432, B1 => n41218, B2 =>
                           n40425, C1 => n40419, C2 => n38837, ZN => n9339);
   U32835 : OAI222_X1 port map( A1 => n40840, A2 => n40431, B1 => n41224, B2 =>
                           n40424, C1 => n40419, C2 => n38838, ZN => n9338);
   U32836 : OAI222_X1 port map( A1 => n40846, A2 => n40431, B1 => n41230, B2 =>
                           n40424, C1 => n40419, C2 => n38839, ZN => n9337);
   U32837 : OAI222_X1 port map( A1 => n40852, A2 => n40431, B1 => n41236, B2 =>
                           n40424, C1 => n40419, C2 => n38840, ZN => n9336);
   U32838 : OAI222_X1 port map( A1 => n40858, A2 => n40431, B1 => n41242, B2 =>
                           n40424, C1 => n40419, C2 => n38841, ZN => n9335);
   U32839 : OAI222_X1 port map( A1 => n40864, A2 => n40431, B1 => n41248, B2 =>
                           n40424, C1 => n40419, C2 => n38842, ZN => n9334);
   U32840 : OAI222_X1 port map( A1 => n40870, A2 => n40431, B1 => n41254, B2 =>
                           n40424, C1 => n40419, C2 => n38843, ZN => n9333);
   U32841 : OAI222_X1 port map( A1 => n40876, A2 => n40431, B1 => n41260, B2 =>
                           n40424, C1 => n40419, C2 => n38844, ZN => n9332);
   U32842 : OAI222_X1 port map( A1 => n40882, A2 => n40431, B1 => n41266, B2 =>
                           n40424, C1 => n40419, C2 => n38845, ZN => n9331);
   U32843 : OAI222_X1 port map( A1 => n40888, A2 => n40431, B1 => n41272, B2 =>
                           n40424, C1 => n40420, C2 => n38846, ZN => n9330);
   U32844 : OAI222_X1 port map( A1 => n40894, A2 => n40431, B1 => n41278, B2 =>
                           n40424, C1 => n40420, C2 => n38847, ZN => n9329);
   U32845 : OAI222_X1 port map( A1 => n40900, A2 => n40431, B1 => n41284, B2 =>
                           n40424, C1 => n40420, C2 => n38848, ZN => n9328);
   U32846 : OAI222_X1 port map( A1 => n40906, A2 => n40431, B1 => n41290, B2 =>
                           n40424, C1 => n40420, C2 => n38849, ZN => n9327);
   U32847 : OAI222_X1 port map( A1 => n40912, A2 => n40410, B1 => n41296, B2 =>
                           n40403, C1 => n40400, C2 => n38927, ZN => n9262);
   U32848 : OAI222_X1 port map( A1 => n40918, A2 => n40410, B1 => n41302, B2 =>
                           n40403, C1 => n40400, C2 => n38928, ZN => n9261);
   U32849 : OAI222_X1 port map( A1 => n40924, A2 => n40410, B1 => n41308, B2 =>
                           n40403, C1 => n40400, C2 => n38929, ZN => n9260);
   U32850 : OAI222_X1 port map( A1 => n40930, A2 => n40410, B1 => n41314, B2 =>
                           n40403, C1 => n40400, C2 => n38930, ZN => n9259);
   U32851 : OAI222_X1 port map( A1 => n40936, A2 => n40410, B1 => n41320, B2 =>
                           n40403, C1 => n40400, C2 => n38931, ZN => n9258);
   U32852 : OAI222_X1 port map( A1 => n40942, A2 => n40410, B1 => n41326, B2 =>
                           n40403, C1 => n40400, C2 => n38932, ZN => n9257);
   U32853 : OAI222_X1 port map( A1 => n40948, A2 => n40410, B1 => n41332, B2 =>
                           n40403, C1 => n40400, C2 => n38933, ZN => n9256);
   U32854 : OAI222_X1 port map( A1 => n40960, A2 => n40410, B1 => n41344, B2 =>
                           n40403, C1 => n40400, C2 => n38934, ZN => n9254);
   U32855 : OAI222_X1 port map( A1 => n40911, A2 => n40210, B1 => n41295, B2 =>
                           n40203, C1 => n40200, C2 => n33110, ZN => n8622);
   U32856 : OAI222_X1 port map( A1 => n40917, A2 => n40210, B1 => n41301, B2 =>
                           n40203, C1 => n40200, C2 => n33109, ZN => n8621);
   U32857 : OAI222_X1 port map( A1 => n40923, A2 => n40210, B1 => n41307, B2 =>
                           n40203, C1 => n40200, C2 => n33108, ZN => n8620);
   U32858 : OAI222_X1 port map( A1 => n40929, A2 => n40210, B1 => n41313, B2 =>
                           n40203, C1 => n40200, C2 => n33107, ZN => n8619);
   U32859 : OAI222_X1 port map( A1 => n40935, A2 => n40210, B1 => n41319, B2 =>
                           n40203, C1 => n40200, C2 => n33106, ZN => n8618);
   U32860 : OAI222_X1 port map( A1 => n40941, A2 => n40210, B1 => n41325, B2 =>
                           n40203, C1 => n40200, C2 => n33105, ZN => n8617);
   U32861 : OAI222_X1 port map( A1 => n40947, A2 => n40210, B1 => n41331, B2 =>
                           n40203, C1 => n40200, C2 => n33104, ZN => n8616);
   U32862 : OAI222_X1 port map( A1 => n40959, A2 => n40210, B1 => n41343, B2 =>
                           n40203, C1 => n40200, C2 => n33102, ZN => n8614);
   U32863 : OAI222_X1 port map( A1 => n40911, A2 => n40230, B1 => n41295, B2 =>
                           n40223, C1 => n40220, C2 => n33098, ZN => n8686);
   U32864 : OAI222_X1 port map( A1 => n40917, A2 => n40230, B1 => n41301, B2 =>
                           n40223, C1 => n40220, C2 => n33097, ZN => n8685);
   U32865 : OAI222_X1 port map( A1 => n40923, A2 => n40230, B1 => n41307, B2 =>
                           n40223, C1 => n40220, C2 => n33096, ZN => n8684);
   U32866 : OAI222_X1 port map( A1 => n40929, A2 => n40230, B1 => n41313, B2 =>
                           n40223, C1 => n40220, C2 => n33095, ZN => n8683);
   U32867 : OAI222_X1 port map( A1 => n40935, A2 => n40230, B1 => n41319, B2 =>
                           n40223, C1 => n40220, C2 => n33094, ZN => n8682);
   U32868 : OAI222_X1 port map( A1 => n40941, A2 => n40230, B1 => n41325, B2 =>
                           n40223, C1 => n40220, C2 => n33093, ZN => n8681);
   U32869 : OAI222_X1 port map( A1 => n40947, A2 => n40230, B1 => n41331, B2 =>
                           n40223, C1 => n40220, C2 => n33092, ZN => n8680);
   U32870 : OAI222_X1 port map( A1 => n40959, A2 => n40230, B1 => n41343, B2 =>
                           n40223, C1 => n40220, C2 => n33090, ZN => n8678);
   U32871 : OAI222_X1 port map( A1 => n40624, A2 => n40414, B1 => n41008, B2 =>
                           n40407, C1 => n40396, C2 => n38935, ZN => n9310);
   U32872 : OAI222_X1 port map( A1 => n40630, A2 => n40414, B1 => n41014, B2 =>
                           n40407, C1 => n40396, C2 => n38936, ZN => n9309);
   U32873 : OAI222_X1 port map( A1 => n40636, A2 => n40414, B1 => n41020, B2 =>
                           n40407, C1 => n40396, C2 => n38937, ZN => n9308);
   U32874 : OAI222_X1 port map( A1 => n40642, A2 => n40414, B1 => n41026, B2 =>
                           n40407, C1 => n40396, C2 => n38938, ZN => n9307);
   U32875 : OAI222_X1 port map( A1 => n40648, A2 => n40414, B1 => n41032, B2 =>
                           n40407, C1 => n40396, C2 => n38939, ZN => n9306);
   U32876 : OAI222_X1 port map( A1 => n40654, A2 => n40414, B1 => n41038, B2 =>
                           n40407, C1 => n40396, C2 => n38940, ZN => n9305);
   U32877 : OAI222_X1 port map( A1 => n40660, A2 => n40414, B1 => n41044, B2 =>
                           n40407, C1 => n40396, C2 => n38941, ZN => n9304);
   U32878 : OAI222_X1 port map( A1 => n40666, A2 => n40414, B1 => n41050, B2 =>
                           n40407, C1 => n40396, C2 => n38942, ZN => n9303);
   U32879 : OAI222_X1 port map( A1 => n40672, A2 => n40414, B1 => n41056, B2 =>
                           n40407, C1 => n40397, C2 => n38943, ZN => n9302);
   U32880 : OAI222_X1 port map( A1 => n40678, A2 => n40414, B1 => n41062, B2 =>
                           n40407, C1 => n40397, C2 => n38944, ZN => n9301);
   U32881 : OAI222_X1 port map( A1 => n40684, A2 => n40414, B1 => n41068, B2 =>
                           n40407, C1 => n40397, C2 => n38945, ZN => n9300);
   U32882 : OAI222_X1 port map( A1 => n40690, A2 => n40414, B1 => n41074, B2 =>
                           n40407, C1 => n40398, C2 => n38946, ZN => n9299);
   U32883 : OAI222_X1 port map( A1 => n40696, A2 => n40413, B1 => n41080, B2 =>
                           n40406, C1 => n40397, C2 => n38947, ZN => n9298);
   U32884 : OAI222_X1 port map( A1 => n40702, A2 => n40413, B1 => n41086, B2 =>
                           n40406, C1 => n40397, C2 => n38948, ZN => n9297);
   U32885 : OAI222_X1 port map( A1 => n40708, A2 => n40413, B1 => n41092, B2 =>
                           n40406, C1 => n40397, C2 => n38949, ZN => n9296);
   U32886 : OAI222_X1 port map( A1 => n40714, A2 => n40413, B1 => n41098, B2 =>
                           n40406, C1 => n40397, C2 => n38950, ZN => n9295);
   U32887 : OAI222_X1 port map( A1 => n40720, A2 => n40413, B1 => n41104, B2 =>
                           n40406, C1 => n40397, C2 => n38951, ZN => n9294);
   U32888 : OAI222_X1 port map( A1 => n40726, A2 => n40413, B1 => n41110, B2 =>
                           n40406, C1 => n40397, C2 => n38952, ZN => n9293);
   U32889 : OAI222_X1 port map( A1 => n40732, A2 => n40413, B1 => n41116, B2 =>
                           n40406, C1 => n40397, C2 => n38953, ZN => n9292);
   U32890 : OAI222_X1 port map( A1 => n40738, A2 => n40413, B1 => n41122, B2 =>
                           n40406, C1 => n40397, C2 => n38954, ZN => n9291);
   U32891 : OAI222_X1 port map( A1 => n40744, A2 => n40413, B1 => n41128, B2 =>
                           n40406, C1 => n40397, C2 => n38955, ZN => n9290);
   U32892 : OAI222_X1 port map( A1 => n40750, A2 => n40413, B1 => n41134, B2 =>
                           n40406, C1 => n40398, C2 => n38956, ZN => n9289);
   U32893 : OAI222_X1 port map( A1 => n40756, A2 => n40413, B1 => n41140, B2 =>
                           n40406, C1 => n40398, C2 => n38957, ZN => n9288);
   U32894 : OAI222_X1 port map( A1 => n40762, A2 => n40413, B1 => n41146, B2 =>
                           n40406, C1 => n40398, C2 => n38958, ZN => n9287);
   U32895 : OAI222_X1 port map( A1 => n40768, A2 => n40412, B1 => n41152, B2 =>
                           n40405, C1 => n40398, C2 => n38959, ZN => n9286);
   U32896 : OAI222_X1 port map( A1 => n40774, A2 => n40412, B1 => n41158, B2 =>
                           n40405, C1 => n40398, C2 => n38960, ZN => n9285);
   U32897 : OAI222_X1 port map( A1 => n40780, A2 => n40412, B1 => n41164, B2 =>
                           n40405, C1 => n40398, C2 => n38961, ZN => n9284);
   U32898 : OAI222_X1 port map( A1 => n40786, A2 => n40412, B1 => n41170, B2 =>
                           n40405, C1 => n40398, C2 => n38962, ZN => n9283);
   U32899 : OAI222_X1 port map( A1 => n40792, A2 => n40412, B1 => n41176, B2 =>
                           n40405, C1 => n40398, C2 => n38963, ZN => n9282);
   U32900 : OAI222_X1 port map( A1 => n40798, A2 => n40412, B1 => n41182, B2 =>
                           n40405, C1 => n40398, C2 => n38964, ZN => n9281);
   U32901 : OAI222_X1 port map( A1 => n40804, A2 => n40412, B1 => n41188, B2 =>
                           n40405, C1 => n40398, C2 => n38965, ZN => n9280);
   U32902 : OAI222_X1 port map( A1 => n40810, A2 => n40412, B1 => n41194, B2 =>
                           n40405, C1 => n40398, C2 => n38966, ZN => n9279);
   U32903 : OAI222_X1 port map( A1 => n40816, A2 => n40412, B1 => n41200, B2 =>
                           n40405, C1 => n40399, C2 => n38967, ZN => n9278);
   U32904 : OAI222_X1 port map( A1 => n40822, A2 => n40412, B1 => n41206, B2 =>
                           n40405, C1 => n40399, C2 => n38968, ZN => n9277);
   U32905 : OAI222_X1 port map( A1 => n40828, A2 => n40412, B1 => n41212, B2 =>
                           n40405, C1 => n40399, C2 => n38969, ZN => n9276);
   U32906 : OAI222_X1 port map( A1 => n40834, A2 => n40412, B1 => n41218, B2 =>
                           n40405, C1 => n40399, C2 => n38970, ZN => n9275);
   U32907 : OAI222_X1 port map( A1 => n40840, A2 => n40411, B1 => n41224, B2 =>
                           n40404, C1 => n40399, C2 => n38971, ZN => n9274);
   U32908 : OAI222_X1 port map( A1 => n40846, A2 => n40411, B1 => n41230, B2 =>
                           n40404, C1 => n40399, C2 => n38972, ZN => n9273);
   U32909 : OAI222_X1 port map( A1 => n40852, A2 => n40411, B1 => n41236, B2 =>
                           n40404, C1 => n40399, C2 => n38973, ZN => n9272);
   U32910 : OAI222_X1 port map( A1 => n40858, A2 => n40411, B1 => n41242, B2 =>
                           n40404, C1 => n40399, C2 => n38974, ZN => n9271);
   U32911 : OAI222_X1 port map( A1 => n40864, A2 => n40411, B1 => n41248, B2 =>
                           n40404, C1 => n40399, C2 => n38975, ZN => n9270);
   U32912 : OAI222_X1 port map( A1 => n40870, A2 => n40411, B1 => n41254, B2 =>
                           n40404, C1 => n40399, C2 => n38976, ZN => n9269);
   U32913 : OAI222_X1 port map( A1 => n40876, A2 => n40411, B1 => n41260, B2 =>
                           n40404, C1 => n40399, C2 => n38977, ZN => n9268);
   U32914 : OAI222_X1 port map( A1 => n40882, A2 => n40411, B1 => n41266, B2 =>
                           n40404, C1 => n40399, C2 => n38978, ZN => n9267);
   U32915 : OAI222_X1 port map( A1 => n40888, A2 => n40411, B1 => n41272, B2 =>
                           n40404, C1 => n40400, C2 => n38979, ZN => n9266);
   U32916 : OAI222_X1 port map( A1 => n40894, A2 => n40411, B1 => n41278, B2 =>
                           n40404, C1 => n40400, C2 => n38980, ZN => n9265);
   U32917 : OAI222_X1 port map( A1 => n40900, A2 => n40411, B1 => n41284, B2 =>
                           n40404, C1 => n40400, C2 => n38981, ZN => n9264);
   U32918 : OAI222_X1 port map( A1 => n40906, A2 => n40411, B1 => n41290, B2 =>
                           n40404, C1 => n40400, C2 => n38982, ZN => n9263);
   U32919 : OAI222_X1 port map( A1 => n40623, A2 => n40214, B1 => n41007, B2 =>
                           n40207, C1 => n40196, C2 => n32942, ZN => n8670);
   U32920 : OAI222_X1 port map( A1 => n40629, A2 => n40214, B1 => n41013, B2 =>
                           n40207, C1 => n40196, C2 => n32941, ZN => n8669);
   U32921 : OAI222_X1 port map( A1 => n40635, A2 => n40214, B1 => n41019, B2 =>
                           n40207, C1 => n40196, C2 => n32940, ZN => n8668);
   U32922 : OAI222_X1 port map( A1 => n40641, A2 => n40214, B1 => n41025, B2 =>
                           n40207, C1 => n40196, C2 => n32939, ZN => n8667);
   U32923 : OAI222_X1 port map( A1 => n40647, A2 => n40214, B1 => n41031, B2 =>
                           n40207, C1 => n40196, C2 => n32938, ZN => n8666);
   U32924 : OAI222_X1 port map( A1 => n40653, A2 => n40214, B1 => n41037, B2 =>
                           n40207, C1 => n40196, C2 => n32937, ZN => n8665);
   U32925 : OAI222_X1 port map( A1 => n40659, A2 => n40214, B1 => n41043, B2 =>
                           n40207, C1 => n40196, C2 => n32936, ZN => n8664);
   U32926 : OAI222_X1 port map( A1 => n40665, A2 => n40214, B1 => n41049, B2 =>
                           n40207, C1 => n40196, C2 => n32935, ZN => n8663);
   U32927 : OAI222_X1 port map( A1 => n40671, A2 => n40214, B1 => n41055, B2 =>
                           n40207, C1 => n40197, C2 => n32934, ZN => n8662);
   U32928 : OAI222_X1 port map( A1 => n40677, A2 => n40214, B1 => n41061, B2 =>
                           n40207, C1 => n40197, C2 => n32933, ZN => n8661);
   U32929 : OAI222_X1 port map( A1 => n40683, A2 => n40214, B1 => n41067, B2 =>
                           n40207, C1 => n40197, C2 => n32932, ZN => n8660);
   U32930 : OAI222_X1 port map( A1 => n40689, A2 => n40214, B1 => n41073, B2 =>
                           n40207, C1 => n40198, C2 => n32931, ZN => n8659);
   U32931 : OAI222_X1 port map( A1 => n40695, A2 => n40213, B1 => n41079, B2 =>
                           n40206, C1 => n40197, C2 => n32930, ZN => n8658);
   U32932 : OAI222_X1 port map( A1 => n40701, A2 => n40213, B1 => n41085, B2 =>
                           n40206, C1 => n40197, C2 => n32929, ZN => n8657);
   U32933 : OAI222_X1 port map( A1 => n40707, A2 => n40213, B1 => n41091, B2 =>
                           n40206, C1 => n40197, C2 => n32928, ZN => n8656);
   U32934 : OAI222_X1 port map( A1 => n40713, A2 => n40213, B1 => n41097, B2 =>
                           n40206, C1 => n40197, C2 => n32927, ZN => n8655);
   U32935 : OAI222_X1 port map( A1 => n40719, A2 => n40213, B1 => n41103, B2 =>
                           n40206, C1 => n40197, C2 => n32926, ZN => n8654);
   U32936 : OAI222_X1 port map( A1 => n40725, A2 => n40213, B1 => n41109, B2 =>
                           n40206, C1 => n40197, C2 => n32925, ZN => n8653);
   U32937 : OAI222_X1 port map( A1 => n40731, A2 => n40213, B1 => n41115, B2 =>
                           n40206, C1 => n40197, C2 => n32924, ZN => n8652);
   U32938 : OAI222_X1 port map( A1 => n40737, A2 => n40213, B1 => n41121, B2 =>
                           n40206, C1 => n40197, C2 => n32923, ZN => n8651);
   U32939 : OAI222_X1 port map( A1 => n40743, A2 => n40213, B1 => n41127, B2 =>
                           n40206, C1 => n40197, C2 => n32922, ZN => n8650);
   U32940 : OAI222_X1 port map( A1 => n40749, A2 => n40213, B1 => n41133, B2 =>
                           n40206, C1 => n40198, C2 => n32921, ZN => n8649);
   U32941 : OAI222_X1 port map( A1 => n40755, A2 => n40213, B1 => n41139, B2 =>
                           n40206, C1 => n40198, C2 => n32920, ZN => n8648);
   U32942 : OAI222_X1 port map( A1 => n40761, A2 => n40213, B1 => n41145, B2 =>
                           n40206, C1 => n40198, C2 => n32919, ZN => n8647);
   U32943 : OAI222_X1 port map( A1 => n40767, A2 => n40212, B1 => n41151, B2 =>
                           n40205, C1 => n40198, C2 => n32918, ZN => n8646);
   U32944 : OAI222_X1 port map( A1 => n40773, A2 => n40212, B1 => n41157, B2 =>
                           n40205, C1 => n40198, C2 => n32917, ZN => n8645);
   U32945 : OAI222_X1 port map( A1 => n40779, A2 => n40212, B1 => n41163, B2 =>
                           n40205, C1 => n40198, C2 => n32916, ZN => n8644);
   U32946 : OAI222_X1 port map( A1 => n40785, A2 => n40212, B1 => n41169, B2 =>
                           n40205, C1 => n40198, C2 => n32915, ZN => n8643);
   U32947 : OAI222_X1 port map( A1 => n40791, A2 => n40212, B1 => n41175, B2 =>
                           n40205, C1 => n40198, C2 => n32914, ZN => n8642);
   U32948 : OAI222_X1 port map( A1 => n40797, A2 => n40212, B1 => n41181, B2 =>
                           n40205, C1 => n40198, C2 => n32913, ZN => n8641);
   U32949 : OAI222_X1 port map( A1 => n40803, A2 => n40212, B1 => n41187, B2 =>
                           n40205, C1 => n40198, C2 => n32912, ZN => n8640);
   U32950 : OAI222_X1 port map( A1 => n40809, A2 => n40212, B1 => n41193, B2 =>
                           n40205, C1 => n40198, C2 => n32911, ZN => n8639);
   U32951 : OAI222_X1 port map( A1 => n40815, A2 => n40212, B1 => n41199, B2 =>
                           n40205, C1 => n40199, C2 => n32910, ZN => n8638);
   U32952 : OAI222_X1 port map( A1 => n40821, A2 => n40212, B1 => n41205, B2 =>
                           n40205, C1 => n40199, C2 => n32909, ZN => n8637);
   U32953 : OAI222_X1 port map( A1 => n40827, A2 => n40212, B1 => n41211, B2 =>
                           n40205, C1 => n40199, C2 => n32908, ZN => n8636);
   U32954 : OAI222_X1 port map( A1 => n40833, A2 => n40212, B1 => n41217, B2 =>
                           n40205, C1 => n40199, C2 => n32907, ZN => n8635);
   U32955 : OAI222_X1 port map( A1 => n40839, A2 => n40211, B1 => n41223, B2 =>
                           n40204, C1 => n40199, C2 => n32906, ZN => n8634);
   U32956 : OAI222_X1 port map( A1 => n40845, A2 => n40211, B1 => n41229, B2 =>
                           n40204, C1 => n40199, C2 => n32905, ZN => n8633);
   U32957 : OAI222_X1 port map( A1 => n40851, A2 => n40211, B1 => n41235, B2 =>
                           n40204, C1 => n40199, C2 => n32904, ZN => n8632);
   U32958 : OAI222_X1 port map( A1 => n40857, A2 => n40211, B1 => n41241, B2 =>
                           n40204, C1 => n40199, C2 => n32903, ZN => n8631);
   U32959 : OAI222_X1 port map( A1 => n40863, A2 => n40211, B1 => n41247, B2 =>
                           n40204, C1 => n40199, C2 => n32902, ZN => n8630);
   U32960 : OAI222_X1 port map( A1 => n40869, A2 => n40211, B1 => n41253, B2 =>
                           n40204, C1 => n40199, C2 => n32901, ZN => n8629);
   U32961 : OAI222_X1 port map( A1 => n40875, A2 => n40211, B1 => n41259, B2 =>
                           n40204, C1 => n40199, C2 => n32900, ZN => n8628);
   U32962 : OAI222_X1 port map( A1 => n40881, A2 => n40211, B1 => n41265, B2 =>
                           n40204, C1 => n40199, C2 => n32899, ZN => n8627);
   U32963 : OAI222_X1 port map( A1 => n40887, A2 => n40211, B1 => n41271, B2 =>
                           n40204, C1 => n40200, C2 => n32898, ZN => n8626);
   U32964 : OAI222_X1 port map( A1 => n40893, A2 => n40211, B1 => n41277, B2 =>
                           n40204, C1 => n40200, C2 => n32897, ZN => n8625);
   U32965 : OAI222_X1 port map( A1 => n40899, A2 => n40211, B1 => n41283, B2 =>
                           n40204, C1 => n40200, C2 => n32896, ZN => n8624);
   U32966 : OAI222_X1 port map( A1 => n40905, A2 => n40211, B1 => n41289, B2 =>
                           n40204, C1 => n40200, C2 => n32895, ZN => n8623);
   U32967 : OAI222_X1 port map( A1 => n40623, A2 => n40234, B1 => n41007, B2 =>
                           n40227, C1 => n40216, C2 => n32894, ZN => n8734);
   U32968 : OAI222_X1 port map( A1 => n40629, A2 => n40234, B1 => n41013, B2 =>
                           n40227, C1 => n40216, C2 => n32893, ZN => n8733);
   U32969 : OAI222_X1 port map( A1 => n40635, A2 => n40234, B1 => n41019, B2 =>
                           n40227, C1 => n40216, C2 => n32892, ZN => n8732);
   U32970 : OAI222_X1 port map( A1 => n40641, A2 => n40234, B1 => n41025, B2 =>
                           n40227, C1 => n40216, C2 => n32891, ZN => n8731);
   U32971 : OAI222_X1 port map( A1 => n40647, A2 => n40234, B1 => n41031, B2 =>
                           n40227, C1 => n40216, C2 => n32890, ZN => n8730);
   U32972 : OAI222_X1 port map( A1 => n40653, A2 => n40234, B1 => n41037, B2 =>
                           n40227, C1 => n40216, C2 => n32889, ZN => n8729);
   U32973 : OAI222_X1 port map( A1 => n40659, A2 => n40234, B1 => n41043, B2 =>
                           n40227, C1 => n40216, C2 => n32888, ZN => n8728);
   U32974 : OAI222_X1 port map( A1 => n40665, A2 => n40234, B1 => n41049, B2 =>
                           n40227, C1 => n40216, C2 => n32887, ZN => n8727);
   U32975 : OAI222_X1 port map( A1 => n40671, A2 => n40234, B1 => n41055, B2 =>
                           n40227, C1 => n40217, C2 => n32886, ZN => n8726);
   U32976 : OAI222_X1 port map( A1 => n40677, A2 => n40234, B1 => n41061, B2 =>
                           n40227, C1 => n40217, C2 => n32885, ZN => n8725);
   U32977 : OAI222_X1 port map( A1 => n40683, A2 => n40234, B1 => n41067, B2 =>
                           n40227, C1 => n40217, C2 => n32884, ZN => n8724);
   U32978 : OAI222_X1 port map( A1 => n40689, A2 => n40234, B1 => n41073, B2 =>
                           n40227, C1 => n40218, C2 => n32883, ZN => n8723);
   U32979 : OAI222_X1 port map( A1 => n40695, A2 => n40233, B1 => n41079, B2 =>
                           n40226, C1 => n40217, C2 => n32882, ZN => n8722);
   U32980 : OAI222_X1 port map( A1 => n40701, A2 => n40233, B1 => n41085, B2 =>
                           n40226, C1 => n40217, C2 => n32881, ZN => n8721);
   U32981 : OAI222_X1 port map( A1 => n40707, A2 => n40233, B1 => n41091, B2 =>
                           n40226, C1 => n40217, C2 => n32880, ZN => n8720);
   U32982 : OAI222_X1 port map( A1 => n40713, A2 => n40233, B1 => n41097, B2 =>
                           n40226, C1 => n40217, C2 => n32879, ZN => n8719);
   U32983 : OAI222_X1 port map( A1 => n40719, A2 => n40233, B1 => n41103, B2 =>
                           n40226, C1 => n40217, C2 => n32878, ZN => n8718);
   U32984 : OAI222_X1 port map( A1 => n40725, A2 => n40233, B1 => n41109, B2 =>
                           n40226, C1 => n40217, C2 => n32877, ZN => n8717);
   U32985 : OAI222_X1 port map( A1 => n40731, A2 => n40233, B1 => n41115, B2 =>
                           n40226, C1 => n40217, C2 => n32876, ZN => n8716);
   U32986 : OAI222_X1 port map( A1 => n40737, A2 => n40233, B1 => n41121, B2 =>
                           n40226, C1 => n40217, C2 => n32875, ZN => n8715);
   U32987 : OAI222_X1 port map( A1 => n40743, A2 => n40233, B1 => n41127, B2 =>
                           n40226, C1 => n40217, C2 => n32874, ZN => n8714);
   U32988 : OAI222_X1 port map( A1 => n40749, A2 => n40233, B1 => n41133, B2 =>
                           n40226, C1 => n40218, C2 => n32873, ZN => n8713);
   U32989 : OAI222_X1 port map( A1 => n40755, A2 => n40233, B1 => n41139, B2 =>
                           n40226, C1 => n40218, C2 => n32872, ZN => n8712);
   U32990 : OAI222_X1 port map( A1 => n40761, A2 => n40233, B1 => n41145, B2 =>
                           n40226, C1 => n40218, C2 => n32871, ZN => n8711);
   U32991 : OAI222_X1 port map( A1 => n40767, A2 => n40232, B1 => n41151, B2 =>
                           n40225, C1 => n40218, C2 => n32870, ZN => n8710);
   U32992 : OAI222_X1 port map( A1 => n40773, A2 => n40232, B1 => n41157, B2 =>
                           n40225, C1 => n40218, C2 => n32869, ZN => n8709);
   U32993 : OAI222_X1 port map( A1 => n40779, A2 => n40232, B1 => n41163, B2 =>
                           n40225, C1 => n40218, C2 => n32868, ZN => n8708);
   U32994 : OAI222_X1 port map( A1 => n40785, A2 => n40232, B1 => n41169, B2 =>
                           n40225, C1 => n40218, C2 => n32867, ZN => n8707);
   U32995 : OAI222_X1 port map( A1 => n40791, A2 => n40232, B1 => n41175, B2 =>
                           n40225, C1 => n40218, C2 => n32866, ZN => n8706);
   U32996 : OAI222_X1 port map( A1 => n40797, A2 => n40232, B1 => n41181, B2 =>
                           n40225, C1 => n40218, C2 => n32865, ZN => n8705);
   U32997 : OAI222_X1 port map( A1 => n40803, A2 => n40232, B1 => n41187, B2 =>
                           n40225, C1 => n40218, C2 => n32864, ZN => n8704);
   U32998 : OAI222_X1 port map( A1 => n40809, A2 => n40232, B1 => n41193, B2 =>
                           n40225, C1 => n40218, C2 => n32863, ZN => n8703);
   U32999 : OAI222_X1 port map( A1 => n40815, A2 => n40232, B1 => n41199, B2 =>
                           n40225, C1 => n40219, C2 => n32862, ZN => n8702);
   U33000 : OAI222_X1 port map( A1 => n40821, A2 => n40232, B1 => n41205, B2 =>
                           n40225, C1 => n40219, C2 => n32861, ZN => n8701);
   U33001 : OAI222_X1 port map( A1 => n40827, A2 => n40232, B1 => n41211, B2 =>
                           n40225, C1 => n40219, C2 => n32860, ZN => n8700);
   U33002 : OAI222_X1 port map( A1 => n40833, A2 => n40232, B1 => n41217, B2 =>
                           n40225, C1 => n40219, C2 => n32859, ZN => n8699);
   U33003 : OAI222_X1 port map( A1 => n40839, A2 => n40231, B1 => n41223, B2 =>
                           n40224, C1 => n40219, C2 => n32858, ZN => n8698);
   U33004 : OAI222_X1 port map( A1 => n40845, A2 => n40231, B1 => n41229, B2 =>
                           n40224, C1 => n40219, C2 => n32857, ZN => n8697);
   U33005 : OAI222_X1 port map( A1 => n40851, A2 => n40231, B1 => n41235, B2 =>
                           n40224, C1 => n40219, C2 => n32856, ZN => n8696);
   U33006 : OAI222_X1 port map( A1 => n40857, A2 => n40231, B1 => n41241, B2 =>
                           n40224, C1 => n40219, C2 => n32855, ZN => n8695);
   U33007 : OAI222_X1 port map( A1 => n40863, A2 => n40231, B1 => n41247, B2 =>
                           n40224, C1 => n40219, C2 => n32854, ZN => n8694);
   U33008 : OAI222_X1 port map( A1 => n40869, A2 => n40231, B1 => n41253, B2 =>
                           n40224, C1 => n40219, C2 => n32853, ZN => n8693);
   U33009 : OAI222_X1 port map( A1 => n40875, A2 => n40231, B1 => n41259, B2 =>
                           n40224, C1 => n40219, C2 => n32852, ZN => n8692);
   U33010 : OAI222_X1 port map( A1 => n40881, A2 => n40231, B1 => n41265, B2 =>
                           n40224, C1 => n40219, C2 => n32851, ZN => n8691);
   U33011 : OAI222_X1 port map( A1 => n40887, A2 => n40231, B1 => n41271, B2 =>
                           n40224, C1 => n40220, C2 => n32850, ZN => n8690);
   U33012 : OAI222_X1 port map( A1 => n40893, A2 => n40231, B1 => n41277, B2 =>
                           n40224, C1 => n40220, C2 => n32849, ZN => n8689);
   U33013 : OAI222_X1 port map( A1 => n40899, A2 => n40231, B1 => n41283, B2 =>
                           n40224, C1 => n40220, C2 => n32848, ZN => n8688);
   U33014 : OAI222_X1 port map( A1 => n40905, A2 => n40231, B1 => n41289, B2 =>
                           n40224, C1 => n40220, C2 => n32847, ZN => n8687);
   U33015 : OAI222_X1 port map( A1 => n40912, A2 => n40310, B1 => n41296, B2 =>
                           n40303, C1 => n40300, C2 => n32726, ZN => n8942);
   U33016 : OAI222_X1 port map( A1 => n40918, A2 => n40310, B1 => n41302, B2 =>
                           n40303, C1 => n40300, C2 => n32725, ZN => n8941);
   U33017 : OAI222_X1 port map( A1 => n40924, A2 => n40310, B1 => n41308, B2 =>
                           n40303, C1 => n40300, C2 => n32724, ZN => n8940);
   U33018 : OAI222_X1 port map( A1 => n40930, A2 => n40310, B1 => n41314, B2 =>
                           n40303, C1 => n40300, C2 => n32723, ZN => n8939);
   U33019 : OAI222_X1 port map( A1 => n40936, A2 => n40310, B1 => n41320, B2 =>
                           n40303, C1 => n40300, C2 => n32722, ZN => n8938);
   U33020 : OAI222_X1 port map( A1 => n40942, A2 => n40310, B1 => n41326, B2 =>
                           n40303, C1 => n40300, C2 => n32721, ZN => n8937);
   U33021 : OAI222_X1 port map( A1 => n40948, A2 => n40310, B1 => n41332, B2 =>
                           n40303, C1 => n40300, C2 => n32720, ZN => n8936);
   U33022 : OAI222_X1 port map( A1 => n40960, A2 => n40310, B1 => n41344, B2 =>
                           n40303, C1 => n40300, C2 => n32718, ZN => n8934);
   U33023 : OAI222_X1 port map( A1 => n40912, A2 => n40330, B1 => n41296, B2 =>
                           n40323, C1 => n40320, C2 => n32714, ZN => n9006);
   U33024 : OAI222_X1 port map( A1 => n40918, A2 => n40330, B1 => n41302, B2 =>
                           n40323, C1 => n40320, C2 => n32713, ZN => n9005);
   U33025 : OAI222_X1 port map( A1 => n40924, A2 => n40330, B1 => n41308, B2 =>
                           n40323, C1 => n40320, C2 => n32712, ZN => n9004);
   U33026 : OAI222_X1 port map( A1 => n40930, A2 => n40330, B1 => n41314, B2 =>
                           n40323, C1 => n40320, C2 => n32711, ZN => n9003);
   U33027 : OAI222_X1 port map( A1 => n40936, A2 => n40330, B1 => n41320, B2 =>
                           n40323, C1 => n40320, C2 => n32710, ZN => n9002);
   U33028 : OAI222_X1 port map( A1 => n40942, A2 => n40330, B1 => n41326, B2 =>
                           n40323, C1 => n40320, C2 => n32709, ZN => n9001);
   U33029 : OAI222_X1 port map( A1 => n40948, A2 => n40330, B1 => n41332, B2 =>
                           n40323, C1 => n40320, C2 => n32708, ZN => n9000);
   U33030 : OAI222_X1 port map( A1 => n40960, A2 => n40330, B1 => n41344, B2 =>
                           n40323, C1 => n40320, C2 => n32706, ZN => n8998);
   U33031 : OAI222_X1 port map( A1 => n40910, A2 => n39835, B1 => n41294, B2 =>
                           n39828, C1 => n39825, C2 => n32702, ZN => n7406);
   U33032 : OAI222_X1 port map( A1 => n40916, A2 => n39835, B1 => n41300, B2 =>
                           n39828, C1 => n39825, C2 => n32701, ZN => n7405);
   U33033 : OAI222_X1 port map( A1 => n40922, A2 => n39835, B1 => n41306, B2 =>
                           n39828, C1 => n39825, C2 => n32700, ZN => n7404);
   U33034 : OAI222_X1 port map( A1 => n40928, A2 => n39835, B1 => n41312, B2 =>
                           n39828, C1 => n39825, C2 => n32699, ZN => n7403);
   U33035 : OAI222_X1 port map( A1 => n40934, A2 => n39835, B1 => n41318, B2 =>
                           n39828, C1 => n39825, C2 => n32698, ZN => n7402);
   U33036 : OAI222_X1 port map( A1 => n40940, A2 => n39835, B1 => n41324, B2 =>
                           n39828, C1 => n39825, C2 => n32697, ZN => n7401);
   U33037 : OAI222_X1 port map( A1 => n40946, A2 => n39835, B1 => n41330, B2 =>
                           n39828, C1 => n39825, C2 => n32696, ZN => n7400);
   U33038 : OAI222_X1 port map( A1 => n40958, A2 => n39835, B1 => n41342, B2 =>
                           n39828, C1 => n39825, C2 => n32694, ZN => n7398);
   U33039 : OAI222_X1 port map( A1 => n40624, A2 => n40314, B1 => n41008, B2 =>
                           n40307, C1 => n40296, C2 => n32690, ZN => n8990);
   U33040 : OAI222_X1 port map( A1 => n40630, A2 => n40314, B1 => n41014, B2 =>
                           n40307, C1 => n40296, C2 => n32689, ZN => n8989);
   U33041 : OAI222_X1 port map( A1 => n40636, A2 => n40314, B1 => n41020, B2 =>
                           n40307, C1 => n40296, C2 => n32688, ZN => n8988);
   U33042 : OAI222_X1 port map( A1 => n40642, A2 => n40314, B1 => n41026, B2 =>
                           n40307, C1 => n40296, C2 => n32687, ZN => n8987);
   U33043 : OAI222_X1 port map( A1 => n40648, A2 => n40314, B1 => n41032, B2 =>
                           n40307, C1 => n40296, C2 => n32686, ZN => n8986);
   U33044 : OAI222_X1 port map( A1 => n40654, A2 => n40314, B1 => n41038, B2 =>
                           n40307, C1 => n40296, C2 => n32685, ZN => n8985);
   U33045 : OAI222_X1 port map( A1 => n40660, A2 => n40314, B1 => n41044, B2 =>
                           n40307, C1 => n40296, C2 => n32684, ZN => n8984);
   U33046 : OAI222_X1 port map( A1 => n40666, A2 => n40314, B1 => n41050, B2 =>
                           n40307, C1 => n40296, C2 => n32683, ZN => n8983);
   U33047 : OAI222_X1 port map( A1 => n40672, A2 => n40314, B1 => n41056, B2 =>
                           n40307, C1 => n40297, C2 => n32682, ZN => n8982);
   U33048 : OAI222_X1 port map( A1 => n40678, A2 => n40314, B1 => n41062, B2 =>
                           n40307, C1 => n40297, C2 => n32681, ZN => n8981);
   U33049 : OAI222_X1 port map( A1 => n40684, A2 => n40314, B1 => n41068, B2 =>
                           n40307, C1 => n40297, C2 => n32680, ZN => n8980);
   U33050 : OAI222_X1 port map( A1 => n40690, A2 => n40314, B1 => n41074, B2 =>
                           n40307, C1 => n40298, C2 => n32679, ZN => n8979);
   U33051 : OAI222_X1 port map( A1 => n40696, A2 => n40313, B1 => n41080, B2 =>
                           n40306, C1 => n40297, C2 => n32678, ZN => n8978);
   U33052 : OAI222_X1 port map( A1 => n40702, A2 => n40313, B1 => n41086, B2 =>
                           n40306, C1 => n40297, C2 => n32677, ZN => n8977);
   U33053 : OAI222_X1 port map( A1 => n40708, A2 => n40313, B1 => n41092, B2 =>
                           n40306, C1 => n40297, C2 => n32676, ZN => n8976);
   U33054 : OAI222_X1 port map( A1 => n40714, A2 => n40313, B1 => n41098, B2 =>
                           n40306, C1 => n40297, C2 => n32675, ZN => n8975);
   U33055 : OAI222_X1 port map( A1 => n40720, A2 => n40313, B1 => n41104, B2 =>
                           n40306, C1 => n40297, C2 => n32674, ZN => n8974);
   U33056 : OAI222_X1 port map( A1 => n40726, A2 => n40313, B1 => n41110, B2 =>
                           n40306, C1 => n40297, C2 => n32673, ZN => n8973);
   U33057 : OAI222_X1 port map( A1 => n40732, A2 => n40313, B1 => n41116, B2 =>
                           n40306, C1 => n40297, C2 => n32672, ZN => n8972);
   U33058 : OAI222_X1 port map( A1 => n40738, A2 => n40313, B1 => n41122, B2 =>
                           n40306, C1 => n40297, C2 => n32671, ZN => n8971);
   U33059 : OAI222_X1 port map( A1 => n40744, A2 => n40313, B1 => n41128, B2 =>
                           n40306, C1 => n40297, C2 => n32670, ZN => n8970);
   U33060 : OAI222_X1 port map( A1 => n40750, A2 => n40313, B1 => n41134, B2 =>
                           n40306, C1 => n40298, C2 => n32669, ZN => n8969);
   U33061 : OAI222_X1 port map( A1 => n40756, A2 => n40313, B1 => n41140, B2 =>
                           n40306, C1 => n40298, C2 => n32668, ZN => n8968);
   U33062 : OAI222_X1 port map( A1 => n40762, A2 => n40313, B1 => n41146, B2 =>
                           n40306, C1 => n40298, C2 => n32667, ZN => n8967);
   U33063 : OAI222_X1 port map( A1 => n40768, A2 => n40312, B1 => n41152, B2 =>
                           n40305, C1 => n40298, C2 => n32666, ZN => n8966);
   U33064 : OAI222_X1 port map( A1 => n40774, A2 => n40312, B1 => n41158, B2 =>
                           n40305, C1 => n40298, C2 => n32665, ZN => n8965);
   U33065 : OAI222_X1 port map( A1 => n40780, A2 => n40312, B1 => n41164, B2 =>
                           n40305, C1 => n40298, C2 => n32664, ZN => n8964);
   U33066 : OAI222_X1 port map( A1 => n40786, A2 => n40312, B1 => n41170, B2 =>
                           n40305, C1 => n40298, C2 => n32663, ZN => n8963);
   U33067 : OAI222_X1 port map( A1 => n40792, A2 => n40312, B1 => n41176, B2 =>
                           n40305, C1 => n40298, C2 => n32662, ZN => n8962);
   U33068 : OAI222_X1 port map( A1 => n40798, A2 => n40312, B1 => n41182, B2 =>
                           n40305, C1 => n40298, C2 => n32661, ZN => n8961);
   U33069 : OAI222_X1 port map( A1 => n40804, A2 => n40312, B1 => n41188, B2 =>
                           n40305, C1 => n40298, C2 => n32660, ZN => n8960);
   U33070 : OAI222_X1 port map( A1 => n40810, A2 => n40312, B1 => n41194, B2 =>
                           n40305, C1 => n40298, C2 => n32659, ZN => n8959);
   U33071 : OAI222_X1 port map( A1 => n40816, A2 => n40312, B1 => n41200, B2 =>
                           n40305, C1 => n40299, C2 => n32658, ZN => n8958);
   U33072 : OAI222_X1 port map( A1 => n40822, A2 => n40312, B1 => n41206, B2 =>
                           n40305, C1 => n40299, C2 => n32657, ZN => n8957);
   U33073 : OAI222_X1 port map( A1 => n40828, A2 => n40312, B1 => n41212, B2 =>
                           n40305, C1 => n40299, C2 => n32656, ZN => n8956);
   U33074 : OAI222_X1 port map( A1 => n40834, A2 => n40312, B1 => n41218, B2 =>
                           n40305, C1 => n40299, C2 => n32655, ZN => n8955);
   U33075 : OAI222_X1 port map( A1 => n40840, A2 => n40311, B1 => n41224, B2 =>
                           n40304, C1 => n40299, C2 => n32654, ZN => n8954);
   U33076 : OAI222_X1 port map( A1 => n40846, A2 => n40311, B1 => n41230, B2 =>
                           n40304, C1 => n40299, C2 => n32653, ZN => n8953);
   U33077 : OAI222_X1 port map( A1 => n40852, A2 => n40311, B1 => n41236, B2 =>
                           n40304, C1 => n40299, C2 => n32652, ZN => n8952);
   U33078 : OAI222_X1 port map( A1 => n40858, A2 => n40311, B1 => n41242, B2 =>
                           n40304, C1 => n40299, C2 => n32651, ZN => n8951);
   U33079 : OAI222_X1 port map( A1 => n40864, A2 => n40311, B1 => n41248, B2 =>
                           n40304, C1 => n40299, C2 => n32650, ZN => n8950);
   U33080 : OAI222_X1 port map( A1 => n40870, A2 => n40311, B1 => n41254, B2 =>
                           n40304, C1 => n40299, C2 => n32649, ZN => n8949);
   U33081 : OAI222_X1 port map( A1 => n40876, A2 => n40311, B1 => n41260, B2 =>
                           n40304, C1 => n40299, C2 => n32648, ZN => n8948);
   U33082 : OAI222_X1 port map( A1 => n40882, A2 => n40311, B1 => n41266, B2 =>
                           n40304, C1 => n40299, C2 => n32647, ZN => n8947);
   U33083 : OAI222_X1 port map( A1 => n40888, A2 => n40311, B1 => n41272, B2 =>
                           n40304, C1 => n40300, C2 => n32646, ZN => n8946);
   U33084 : OAI222_X1 port map( A1 => n40894, A2 => n40311, B1 => n41278, B2 =>
                           n40304, C1 => n40300, C2 => n32645, ZN => n8945);
   U33085 : OAI222_X1 port map( A1 => n40900, A2 => n40311, B1 => n41284, B2 =>
                           n40304, C1 => n40300, C2 => n32644, ZN => n8944);
   U33086 : OAI222_X1 port map( A1 => n40906, A2 => n40311, B1 => n41290, B2 =>
                           n40304, C1 => n40300, C2 => n32643, ZN => n8943);
   U33087 : OAI222_X1 port map( A1 => n40624, A2 => n40334, B1 => n41008, B2 =>
                           n40327, C1 => n40316, C2 => n32642, ZN => n9054);
   U33088 : OAI222_X1 port map( A1 => n40630, A2 => n40334, B1 => n41014, B2 =>
                           n40327, C1 => n40316, C2 => n32641, ZN => n9053);
   U33089 : OAI222_X1 port map( A1 => n40636, A2 => n40334, B1 => n41020, B2 =>
                           n40327, C1 => n40316, C2 => n32640, ZN => n9052);
   U33090 : OAI222_X1 port map( A1 => n40642, A2 => n40334, B1 => n41026, B2 =>
                           n40327, C1 => n40316, C2 => n32639, ZN => n9051);
   U33091 : OAI222_X1 port map( A1 => n40648, A2 => n40334, B1 => n41032, B2 =>
                           n40327, C1 => n40316, C2 => n32638, ZN => n9050);
   U33092 : OAI222_X1 port map( A1 => n40654, A2 => n40334, B1 => n41038, B2 =>
                           n40327, C1 => n40316, C2 => n32637, ZN => n9049);
   U33093 : OAI222_X1 port map( A1 => n40660, A2 => n40334, B1 => n41044, B2 =>
                           n40327, C1 => n40316, C2 => n32636, ZN => n9048);
   U33094 : OAI222_X1 port map( A1 => n40666, A2 => n40334, B1 => n41050, B2 =>
                           n40327, C1 => n40316, C2 => n32635, ZN => n9047);
   U33095 : OAI222_X1 port map( A1 => n40672, A2 => n40334, B1 => n41056, B2 =>
                           n40327, C1 => n40317, C2 => n32634, ZN => n9046);
   U33096 : OAI222_X1 port map( A1 => n40678, A2 => n40334, B1 => n41062, B2 =>
                           n40327, C1 => n40317, C2 => n32633, ZN => n9045);
   U33097 : OAI222_X1 port map( A1 => n40684, A2 => n40334, B1 => n41068, B2 =>
                           n40327, C1 => n40317, C2 => n32632, ZN => n9044);
   U33098 : OAI222_X1 port map( A1 => n40690, A2 => n40334, B1 => n41074, B2 =>
                           n40327, C1 => n40318, C2 => n32631, ZN => n9043);
   U33099 : OAI222_X1 port map( A1 => n40696, A2 => n40333, B1 => n41080, B2 =>
                           n40326, C1 => n40317, C2 => n32630, ZN => n9042);
   U33100 : OAI222_X1 port map( A1 => n40702, A2 => n40333, B1 => n41086, B2 =>
                           n40326, C1 => n40317, C2 => n32629, ZN => n9041);
   U33101 : OAI222_X1 port map( A1 => n40708, A2 => n40333, B1 => n41092, B2 =>
                           n40326, C1 => n40317, C2 => n32628, ZN => n9040);
   U33102 : OAI222_X1 port map( A1 => n40714, A2 => n40333, B1 => n41098, B2 =>
                           n40326, C1 => n40317, C2 => n32627, ZN => n9039);
   U33103 : OAI222_X1 port map( A1 => n40720, A2 => n40333, B1 => n41104, B2 =>
                           n40326, C1 => n40317, C2 => n32626, ZN => n9038);
   U33104 : OAI222_X1 port map( A1 => n40726, A2 => n40333, B1 => n41110, B2 =>
                           n40326, C1 => n40317, C2 => n32625, ZN => n9037);
   U33105 : OAI222_X1 port map( A1 => n40732, A2 => n40333, B1 => n41116, B2 =>
                           n40326, C1 => n40317, C2 => n32624, ZN => n9036);
   U33106 : OAI222_X1 port map( A1 => n40738, A2 => n40333, B1 => n41122, B2 =>
                           n40326, C1 => n40317, C2 => n32623, ZN => n9035);
   U33107 : OAI222_X1 port map( A1 => n40744, A2 => n40333, B1 => n41128, B2 =>
                           n40326, C1 => n40317, C2 => n32622, ZN => n9034);
   U33108 : OAI222_X1 port map( A1 => n40750, A2 => n40333, B1 => n41134, B2 =>
                           n40326, C1 => n40318, C2 => n32621, ZN => n9033);
   U33109 : OAI222_X1 port map( A1 => n40756, A2 => n40333, B1 => n41140, B2 =>
                           n40326, C1 => n40318, C2 => n32620, ZN => n9032);
   U33110 : OAI222_X1 port map( A1 => n40762, A2 => n40333, B1 => n41146, B2 =>
                           n40326, C1 => n40318, C2 => n32619, ZN => n9031);
   U33111 : OAI222_X1 port map( A1 => n40768, A2 => n40332, B1 => n41152, B2 =>
                           n40325, C1 => n40318, C2 => n32618, ZN => n9030);
   U33112 : OAI222_X1 port map( A1 => n40774, A2 => n40332, B1 => n41158, B2 =>
                           n40325, C1 => n40318, C2 => n32617, ZN => n9029);
   U33113 : OAI222_X1 port map( A1 => n40780, A2 => n40332, B1 => n41164, B2 =>
                           n40325, C1 => n40318, C2 => n32616, ZN => n9028);
   U33114 : OAI222_X1 port map( A1 => n40786, A2 => n40332, B1 => n41170, B2 =>
                           n40325, C1 => n40318, C2 => n32615, ZN => n9027);
   U33115 : OAI222_X1 port map( A1 => n40792, A2 => n40332, B1 => n41176, B2 =>
                           n40325, C1 => n40318, C2 => n32614, ZN => n9026);
   U33116 : OAI222_X1 port map( A1 => n40798, A2 => n40332, B1 => n41182, B2 =>
                           n40325, C1 => n40318, C2 => n32613, ZN => n9025);
   U33117 : OAI222_X1 port map( A1 => n40804, A2 => n40332, B1 => n41188, B2 =>
                           n40325, C1 => n40318, C2 => n32612, ZN => n9024);
   U33118 : OAI222_X1 port map( A1 => n40810, A2 => n40332, B1 => n41194, B2 =>
                           n40325, C1 => n40318, C2 => n32611, ZN => n9023);
   U33119 : OAI222_X1 port map( A1 => n40816, A2 => n40332, B1 => n41200, B2 =>
                           n40325, C1 => n40319, C2 => n32610, ZN => n9022);
   U33120 : OAI222_X1 port map( A1 => n40822, A2 => n40332, B1 => n41206, B2 =>
                           n40325, C1 => n40319, C2 => n32609, ZN => n9021);
   U33121 : OAI222_X1 port map( A1 => n40828, A2 => n40332, B1 => n41212, B2 =>
                           n40325, C1 => n40319, C2 => n32608, ZN => n9020);
   U33122 : OAI222_X1 port map( A1 => n40834, A2 => n40332, B1 => n41218, B2 =>
                           n40325, C1 => n40319, C2 => n32607, ZN => n9019);
   U33123 : OAI222_X1 port map( A1 => n40840, A2 => n40331, B1 => n41224, B2 =>
                           n40324, C1 => n40319, C2 => n32606, ZN => n9018);
   U33124 : OAI222_X1 port map( A1 => n40846, A2 => n40331, B1 => n41230, B2 =>
                           n40324, C1 => n40319, C2 => n32605, ZN => n9017);
   U33125 : OAI222_X1 port map( A1 => n40852, A2 => n40331, B1 => n41236, B2 =>
                           n40324, C1 => n40319, C2 => n32604, ZN => n9016);
   U33126 : OAI222_X1 port map( A1 => n40858, A2 => n40331, B1 => n41242, B2 =>
                           n40324, C1 => n40319, C2 => n32603, ZN => n9015);
   U33127 : OAI222_X1 port map( A1 => n40864, A2 => n40331, B1 => n41248, B2 =>
                           n40324, C1 => n40319, C2 => n32602, ZN => n9014);
   U33128 : OAI222_X1 port map( A1 => n40870, A2 => n40331, B1 => n41254, B2 =>
                           n40324, C1 => n40319, C2 => n32601, ZN => n9013);
   U33129 : OAI222_X1 port map( A1 => n40876, A2 => n40331, B1 => n41260, B2 =>
                           n40324, C1 => n40319, C2 => n32600, ZN => n9012);
   U33130 : OAI222_X1 port map( A1 => n40882, A2 => n40331, B1 => n41266, B2 =>
                           n40324, C1 => n40319, C2 => n32599, ZN => n9011);
   U33131 : OAI222_X1 port map( A1 => n40888, A2 => n40331, B1 => n41272, B2 =>
                           n40324, C1 => n40320, C2 => n32598, ZN => n9010);
   U33132 : OAI222_X1 port map( A1 => n40894, A2 => n40331, B1 => n41278, B2 =>
                           n40324, C1 => n40320, C2 => n32597, ZN => n9009);
   U33133 : OAI222_X1 port map( A1 => n40900, A2 => n40331, B1 => n41284, B2 =>
                           n40324, C1 => n40320, C2 => n32596, ZN => n9008);
   U33134 : OAI222_X1 port map( A1 => n40906, A2 => n40331, B1 => n41290, B2 =>
                           n40324, C1 => n40320, C2 => n32595, ZN => n9007);
   U33135 : OAI222_X1 port map( A1 => n40622, A2 => n39839, B1 => n41006, B2 =>
                           n39832, C1 => n39821, C2 => n32594, ZN => n7454);
   U33136 : OAI222_X1 port map( A1 => n40628, A2 => n39839, B1 => n41012, B2 =>
                           n39832, C1 => n39821, C2 => n32593, ZN => n7453);
   U33137 : OAI222_X1 port map( A1 => n40634, A2 => n39839, B1 => n41018, B2 =>
                           n39832, C1 => n39821, C2 => n32592, ZN => n7452);
   U33138 : OAI222_X1 port map( A1 => n40640, A2 => n39839, B1 => n41024, B2 =>
                           n39832, C1 => n39821, C2 => n32591, ZN => n7451);
   U33139 : OAI222_X1 port map( A1 => n40646, A2 => n39839, B1 => n41030, B2 =>
                           n39832, C1 => n39821, C2 => n32590, ZN => n7450);
   U33140 : OAI222_X1 port map( A1 => n40652, A2 => n39839, B1 => n41036, B2 =>
                           n39832, C1 => n39821, C2 => n32589, ZN => n7449);
   U33141 : OAI222_X1 port map( A1 => n40658, A2 => n39839, B1 => n41042, B2 =>
                           n39832, C1 => n39821, C2 => n32588, ZN => n7448);
   U33142 : OAI222_X1 port map( A1 => n40664, A2 => n39839, B1 => n41048, B2 =>
                           n39832, C1 => n39821, C2 => n32587, ZN => n7447);
   U33143 : OAI222_X1 port map( A1 => n40670, A2 => n39839, B1 => n41054, B2 =>
                           n39832, C1 => n39822, C2 => n32586, ZN => n7446);
   U33144 : OAI222_X1 port map( A1 => n40676, A2 => n39839, B1 => n41060, B2 =>
                           n39832, C1 => n39822, C2 => n32585, ZN => n7445);
   U33145 : OAI222_X1 port map( A1 => n40682, A2 => n39839, B1 => n41066, B2 =>
                           n39832, C1 => n39822, C2 => n32584, ZN => n7444);
   U33146 : OAI222_X1 port map( A1 => n40688, A2 => n39839, B1 => n41072, B2 =>
                           n39832, C1 => n39823, C2 => n32583, ZN => n7443);
   U33147 : OAI222_X1 port map( A1 => n40694, A2 => n39838, B1 => n41078, B2 =>
                           n39831, C1 => n39822, C2 => n32582, ZN => n7442);
   U33148 : OAI222_X1 port map( A1 => n40700, A2 => n39838, B1 => n41084, B2 =>
                           n39831, C1 => n39822, C2 => n32581, ZN => n7441);
   U33149 : OAI222_X1 port map( A1 => n40706, A2 => n39838, B1 => n41090, B2 =>
                           n39831, C1 => n39822, C2 => n32580, ZN => n7440);
   U33150 : OAI222_X1 port map( A1 => n40712, A2 => n39838, B1 => n41096, B2 =>
                           n39831, C1 => n39822, C2 => n32579, ZN => n7439);
   U33151 : OAI222_X1 port map( A1 => n40718, A2 => n39838, B1 => n41102, B2 =>
                           n39831, C1 => n39822, C2 => n32578, ZN => n7438);
   U33152 : OAI222_X1 port map( A1 => n40724, A2 => n39838, B1 => n41108, B2 =>
                           n39831, C1 => n39822, C2 => n32577, ZN => n7437);
   U33153 : OAI222_X1 port map( A1 => n40730, A2 => n39838, B1 => n41114, B2 =>
                           n39831, C1 => n39822, C2 => n32576, ZN => n7436);
   U33154 : OAI222_X1 port map( A1 => n40736, A2 => n39838, B1 => n41120, B2 =>
                           n39831, C1 => n39822, C2 => n32575, ZN => n7435);
   U33155 : OAI222_X1 port map( A1 => n40742, A2 => n39838, B1 => n41126, B2 =>
                           n39831, C1 => n39822, C2 => n32574, ZN => n7434);
   U33156 : OAI222_X1 port map( A1 => n40748, A2 => n39838, B1 => n41132, B2 =>
                           n39831, C1 => n39823, C2 => n32573, ZN => n7433);
   U33157 : OAI222_X1 port map( A1 => n40754, A2 => n39838, B1 => n41138, B2 =>
                           n39831, C1 => n39823, C2 => n32572, ZN => n7432);
   U33158 : OAI222_X1 port map( A1 => n40760, A2 => n39838, B1 => n41144, B2 =>
                           n39831, C1 => n39823, C2 => n32571, ZN => n7431);
   U33159 : OAI222_X1 port map( A1 => n40766, A2 => n39837, B1 => n41150, B2 =>
                           n39830, C1 => n39823, C2 => n32570, ZN => n7430);
   U33160 : OAI222_X1 port map( A1 => n40772, A2 => n39837, B1 => n41156, B2 =>
                           n39830, C1 => n39823, C2 => n32569, ZN => n7429);
   U33161 : OAI222_X1 port map( A1 => n40778, A2 => n39837, B1 => n41162, B2 =>
                           n39830, C1 => n39823, C2 => n32568, ZN => n7428);
   U33162 : OAI222_X1 port map( A1 => n40784, A2 => n39837, B1 => n41168, B2 =>
                           n39830, C1 => n39823, C2 => n32567, ZN => n7427);
   U33163 : OAI222_X1 port map( A1 => n40790, A2 => n39837, B1 => n41174, B2 =>
                           n39830, C1 => n39823, C2 => n32566, ZN => n7426);
   U33164 : OAI222_X1 port map( A1 => n40796, A2 => n39837, B1 => n41180, B2 =>
                           n39830, C1 => n39823, C2 => n32565, ZN => n7425);
   U33165 : OAI222_X1 port map( A1 => n40802, A2 => n39837, B1 => n41186, B2 =>
                           n39830, C1 => n39823, C2 => n32564, ZN => n7424);
   U33166 : OAI222_X1 port map( A1 => n40808, A2 => n39837, B1 => n41192, B2 =>
                           n39830, C1 => n39823, C2 => n32563, ZN => n7423);
   U33167 : OAI222_X1 port map( A1 => n40814, A2 => n39837, B1 => n41198, B2 =>
                           n39830, C1 => n39824, C2 => n32562, ZN => n7422);
   U33168 : OAI222_X1 port map( A1 => n40820, A2 => n39837, B1 => n41204, B2 =>
                           n39830, C1 => n39824, C2 => n32561, ZN => n7421);
   U33169 : OAI222_X1 port map( A1 => n40826, A2 => n39837, B1 => n41210, B2 =>
                           n39830, C1 => n39824, C2 => n32560, ZN => n7420);
   U33170 : OAI222_X1 port map( A1 => n40832, A2 => n39837, B1 => n41216, B2 =>
                           n39830, C1 => n39824, C2 => n32559, ZN => n7419);
   U33171 : OAI222_X1 port map( A1 => n40838, A2 => n39836, B1 => n41222, B2 =>
                           n39829, C1 => n39824, C2 => n32558, ZN => n7418);
   U33172 : OAI222_X1 port map( A1 => n40844, A2 => n39836, B1 => n41228, B2 =>
                           n39829, C1 => n39824, C2 => n32557, ZN => n7417);
   U33173 : OAI222_X1 port map( A1 => n40850, A2 => n39836, B1 => n41234, B2 =>
                           n39829, C1 => n39824, C2 => n32556, ZN => n7416);
   U33174 : OAI222_X1 port map( A1 => n40856, A2 => n39836, B1 => n41240, B2 =>
                           n39829, C1 => n39824, C2 => n32555, ZN => n7415);
   U33175 : OAI222_X1 port map( A1 => n40862, A2 => n39836, B1 => n41246, B2 =>
                           n39829, C1 => n39824, C2 => n32554, ZN => n7414);
   U33176 : OAI222_X1 port map( A1 => n40868, A2 => n39836, B1 => n41252, B2 =>
                           n39829, C1 => n39824, C2 => n32553, ZN => n7413);
   U33177 : OAI222_X1 port map( A1 => n40874, A2 => n39836, B1 => n41258, B2 =>
                           n39829, C1 => n39824, C2 => n32552, ZN => n7412);
   U33178 : OAI222_X1 port map( A1 => n40880, A2 => n39836, B1 => n41264, B2 =>
                           n39829, C1 => n39824, C2 => n32551, ZN => n7411);
   U33179 : OAI222_X1 port map( A1 => n40886, A2 => n39836, B1 => n41270, B2 =>
                           n39829, C1 => n39825, C2 => n32550, ZN => n7410);
   U33180 : OAI222_X1 port map( A1 => n40892, A2 => n39836, B1 => n41276, B2 =>
                           n39829, C1 => n39825, C2 => n32549, ZN => n7409);
   U33181 : OAI222_X1 port map( A1 => n40898, A2 => n39836, B1 => n41282, B2 =>
                           n39829, C1 => n39825, C2 => n32548, ZN => n7408);
   U33182 : OAI222_X1 port map( A1 => n40904, A2 => n39836, B1 => n41288, B2 =>
                           n39829, C1 => n39825, C2 => n32547, ZN => n7407);
   U33183 : OAI222_X1 port map( A1 => n40635, A2 => n40134, B1 => n41019, B2 =>
                           n40127, C1 => n40116, C2 => n38850, ZN => n8412);
   U33184 : OAI222_X1 port map( A1 => n40623, A2 => n40134, B1 => n41007, B2 =>
                           n40127, C1 => n40116, C2 => n38851, ZN => n8414);
   U33185 : OAI222_X1 port map( A1 => n40629, A2 => n40134, B1 => n41013, B2 =>
                           n40127, C1 => n40116, C2 => n38852, ZN => n8413);
   U33186 : OAI222_X1 port map( A1 => n40641, A2 => n40134, B1 => n41025, B2 =>
                           n40127, C1 => n40116, C2 => n38853, ZN => n8411);
   U33187 : OAI222_X1 port map( A1 => n40647, A2 => n40134, B1 => n41031, B2 =>
                           n40127, C1 => n40116, C2 => n38854, ZN => n8410);
   U33188 : OAI222_X1 port map( A1 => n40653, A2 => n40134, B1 => n41037, B2 =>
                           n40127, C1 => n40116, C2 => n38855, ZN => n8409);
   U33189 : OAI222_X1 port map( A1 => n40600, A2 => n40435, B1 => n40984, B2 =>
                           n40428, C1 => n40416, C2 => n38856, ZN => n9378);
   U33190 : OAI222_X1 port map( A1 => n40606, A2 => n40435, B1 => n40990, B2 =>
                           n40428, C1 => n40416, C2 => n38857, ZN => n9377);
   U33191 : OAI222_X1 port map( A1 => n40612, A2 => n40435, B1 => n40996, B2 =>
                           n40428, C1 => n40416, C2 => n38858, ZN => n9376);
   U33192 : OAI222_X1 port map( A1 => n40618, A2 => n40435, B1 => n41002, B2 =>
                           n40428, C1 => n40416, C2 => n38859, ZN => n9375);
   U33193 : OAI222_X1 port map( A1 => n40600, A2 => n40415, B1 => n40984, B2 =>
                           n40408, C1 => n40396, C2 => n38983, ZN => n9314);
   U33194 : OAI222_X1 port map( A1 => n40606, A2 => n40415, B1 => n40990, B2 =>
                           n40408, C1 => n40396, C2 => n38984, ZN => n9313);
   U33195 : OAI222_X1 port map( A1 => n40612, A2 => n40415, B1 => n40996, B2 =>
                           n40408, C1 => n40396, C2 => n38985, ZN => n9312);
   U33196 : OAI222_X1 port map( A1 => n40618, A2 => n40415, B1 => n41002, B2 =>
                           n40408, C1 => n40396, C2 => n38986, ZN => n9311);
   U33197 : OAI222_X1 port map( A1 => n40599, A2 => n40215, B1 => n40983, B2 =>
                           n40208, C1 => n40196, C2 => n32483, ZN => n8674);
   U33198 : OAI222_X1 port map( A1 => n40605, A2 => n40215, B1 => n40989, B2 =>
                           n40208, C1 => n40196, C2 => n32482, ZN => n8673);
   U33199 : OAI222_X1 port map( A1 => n40611, A2 => n40215, B1 => n40995, B2 =>
                           n40208, C1 => n40196, C2 => n32481, ZN => n8672);
   U33200 : OAI222_X1 port map( A1 => n40617, A2 => n40215, B1 => n41001, B2 =>
                           n40208, C1 => n40196, C2 => n32480, ZN => n8671);
   U33201 : OAI222_X1 port map( A1 => n40599, A2 => n40235, B1 => n40983, B2 =>
                           n40228, C1 => n40216, C2 => n32479, ZN => n8738);
   U33202 : OAI222_X1 port map( A1 => n40605, A2 => n40235, B1 => n40989, B2 =>
                           n40228, C1 => n40216, C2 => n32478, ZN => n8737);
   U33203 : OAI222_X1 port map( A1 => n40611, A2 => n40235, B1 => n40995, B2 =>
                           n40228, C1 => n40216, C2 => n32477, ZN => n8736);
   U33204 : OAI222_X1 port map( A1 => n40617, A2 => n40235, B1 => n41001, B2 =>
                           n40228, C1 => n40216, C2 => n32476, ZN => n8735);
   U33205 : OAI222_X1 port map( A1 => n40600, A2 => n40315, B1 => n40984, B2 =>
                           n40308, C1 => n40296, C2 => n32467, ZN => n8994);
   U33206 : OAI222_X1 port map( A1 => n40606, A2 => n40315, B1 => n40990, B2 =>
                           n40308, C1 => n40296, C2 => n32466, ZN => n8993);
   U33207 : OAI222_X1 port map( A1 => n40612, A2 => n40315, B1 => n40996, B2 =>
                           n40308, C1 => n40296, C2 => n32465, ZN => n8992);
   U33208 : OAI222_X1 port map( A1 => n40618, A2 => n40315, B1 => n41002, B2 =>
                           n40308, C1 => n40296, C2 => n32464, ZN => n8991);
   U33209 : OAI222_X1 port map( A1 => n40600, A2 => n40335, B1 => n40984, B2 =>
                           n40328, C1 => n40316, C2 => n32463, ZN => n9058);
   U33210 : OAI222_X1 port map( A1 => n40606, A2 => n40335, B1 => n40990, B2 =>
                           n40328, C1 => n40316, C2 => n32462, ZN => n9057);
   U33211 : OAI222_X1 port map( A1 => n40612, A2 => n40335, B1 => n40996, B2 =>
                           n40328, C1 => n40316, C2 => n32461, ZN => n9056);
   U33212 : OAI222_X1 port map( A1 => n40618, A2 => n40335, B1 => n41002, B2 =>
                           n40328, C1 => n40316, C2 => n32460, ZN => n9055);
   U33213 : OAI222_X1 port map( A1 => n40598, A2 => n39840, B1 => n40982, B2 =>
                           n39833, C1 => n39821, C2 => n32459, ZN => n7458);
   U33214 : OAI222_X1 port map( A1 => n40604, A2 => n39840, B1 => n40988, B2 =>
                           n39833, C1 => n39821, C2 => n32458, ZN => n7457);
   U33215 : OAI222_X1 port map( A1 => n40610, A2 => n39840, B1 => n40994, B2 =>
                           n39833, C1 => n39821, C2 => n32457, ZN => n7456);
   U33216 : OAI222_X1 port map( A1 => n40616, A2 => n39840, B1 => n41000, B2 =>
                           n39833, C1 => n39821, C2 => n32456, ZN => n7455);
   U33217 : OAI222_X1 port map( A1 => n40599, A2 => n40135, B1 => n40983, B2 =>
                           n40128, C1 => n40116, C2 => n38860, ZN => n8418);
   U33218 : OAI222_X1 port map( A1 => n40605, A2 => n40135, B1 => n40989, B2 =>
                           n40128, C1 => n40116, C2 => n38861, ZN => n8417);
   U33219 : OAI222_X1 port map( A1 => n40611, A2 => n40135, B1 => n40995, B2 =>
                           n40128, C1 => n40116, C2 => n38862, ZN => n8416);
   U33220 : OAI222_X1 port map( A1 => n40617, A2 => n40135, B1 => n41001, B2 =>
                           n40128, C1 => n40116, C2 => n38863, ZN => n8415);
   U33221 : OAI222_X1 port map( A1 => n40913, A2 => n40530, B1 => n41297, B2 =>
                           n40523, C1 => n40520, C2 => n38864, ZN => n9646);
   U33222 : OAI222_X1 port map( A1 => n40919, A2 => n40530, B1 => n41303, B2 =>
                           n40523, C1 => n40520, C2 => n38865, ZN => n9645);
   U33223 : OAI222_X1 port map( A1 => n40925, A2 => n40530, B1 => n41309, B2 =>
                           n40523, C1 => n40520, C2 => n38866, ZN => n9644);
   U33224 : OAI222_X1 port map( A1 => n40931, A2 => n40530, B1 => n41315, B2 =>
                           n40523, C1 => n40520, C2 => n38867, ZN => n9643);
   U33225 : OAI222_X1 port map( A1 => n40937, A2 => n40530, B1 => n41321, B2 =>
                           n40523, C1 => n40520, C2 => n38868, ZN => n9642);
   U33226 : OAI222_X1 port map( A1 => n40943, A2 => n40530, B1 => n41327, B2 =>
                           n40523, C1 => n40520, C2 => n38869, ZN => n9641);
   U33227 : OAI222_X1 port map( A1 => n40949, A2 => n40530, B1 => n41333, B2 =>
                           n40523, C1 => n40520, C2 => n38870, ZN => n9640);
   U33228 : OAI222_X1 port map( A1 => n40961, A2 => n40530, B1 => n41345, B2 =>
                           n40523, C1 => n40520, C2 => n38871, ZN => n9638);
   U33229 : OAI222_X1 port map( A1 => n40625, A2 => n40534, B1 => n41009, B2 =>
                           n40527, C1 => n40516, C2 => n38872, ZN => n9694);
   U33230 : OAI222_X1 port map( A1 => n40631, A2 => n40534, B1 => n41015, B2 =>
                           n40527, C1 => n40516, C2 => n38873, ZN => n9693);
   U33231 : OAI222_X1 port map( A1 => n40637, A2 => n40534, B1 => n41021, B2 =>
                           n40527, C1 => n40516, C2 => n38874, ZN => n9692);
   U33232 : OAI222_X1 port map( A1 => n40643, A2 => n40534, B1 => n41027, B2 =>
                           n40527, C1 => n40516, C2 => n38875, ZN => n9691);
   U33233 : OAI222_X1 port map( A1 => n40649, A2 => n40534, B1 => n41033, B2 =>
                           n40527, C1 => n40516, C2 => n38876, ZN => n9690);
   U33234 : OAI222_X1 port map( A1 => n40655, A2 => n40534, B1 => n41039, B2 =>
                           n40527, C1 => n40516, C2 => n38877, ZN => n9689);
   U33235 : OAI222_X1 port map( A1 => n40661, A2 => n40534, B1 => n41045, B2 =>
                           n40527, C1 => n40516, C2 => n38878, ZN => n9688);
   U33236 : OAI222_X1 port map( A1 => n40667, A2 => n40534, B1 => n41051, B2 =>
                           n40527, C1 => n40516, C2 => n38879, ZN => n9687);
   U33237 : OAI222_X1 port map( A1 => n40673, A2 => n40534, B1 => n41057, B2 =>
                           n40527, C1 => n40517, C2 => n38880, ZN => n9686);
   U33238 : OAI222_X1 port map( A1 => n40679, A2 => n40534, B1 => n41063, B2 =>
                           n40527, C1 => n40517, C2 => n38881, ZN => n9685);
   U33239 : OAI222_X1 port map( A1 => n40685, A2 => n40534, B1 => n41069, B2 =>
                           n40527, C1 => n40517, C2 => n38882, ZN => n9684);
   U33240 : OAI222_X1 port map( A1 => n40691, A2 => n40534, B1 => n41075, B2 =>
                           n40527, C1 => n40518, C2 => n38883, ZN => n9683);
   U33241 : OAI222_X1 port map( A1 => n40697, A2 => n40533, B1 => n41081, B2 =>
                           n40526, C1 => n40517, C2 => n38884, ZN => n9682);
   U33242 : OAI222_X1 port map( A1 => n40703, A2 => n40533, B1 => n41087, B2 =>
                           n40526, C1 => n40517, C2 => n38885, ZN => n9681);
   U33243 : OAI222_X1 port map( A1 => n40709, A2 => n40533, B1 => n41093, B2 =>
                           n40526, C1 => n40517, C2 => n38886, ZN => n9680);
   U33244 : OAI222_X1 port map( A1 => n40715, A2 => n40533, B1 => n41099, B2 =>
                           n40526, C1 => n40517, C2 => n38887, ZN => n9679);
   U33245 : OAI222_X1 port map( A1 => n40721, A2 => n40533, B1 => n41105, B2 =>
                           n40526, C1 => n40517, C2 => n38888, ZN => n9678);
   U33246 : OAI222_X1 port map( A1 => n40727, A2 => n40533, B1 => n41111, B2 =>
                           n40526, C1 => n40517, C2 => n38889, ZN => n9677);
   U33247 : OAI222_X1 port map( A1 => n40733, A2 => n40533, B1 => n41117, B2 =>
                           n40526, C1 => n40517, C2 => n38890, ZN => n9676);
   U33248 : OAI222_X1 port map( A1 => n40739, A2 => n40533, B1 => n41123, B2 =>
                           n40526, C1 => n40517, C2 => n38891, ZN => n9675);
   U33249 : OAI222_X1 port map( A1 => n40745, A2 => n40533, B1 => n41129, B2 =>
                           n40526, C1 => n40517, C2 => n38892, ZN => n9674);
   U33250 : OAI222_X1 port map( A1 => n40751, A2 => n40533, B1 => n41135, B2 =>
                           n40526, C1 => n40518, C2 => n38893, ZN => n9673);
   U33251 : OAI222_X1 port map( A1 => n40757, A2 => n40533, B1 => n41141, B2 =>
                           n40526, C1 => n40518, C2 => n38894, ZN => n9672);
   U33252 : OAI222_X1 port map( A1 => n40763, A2 => n40533, B1 => n41147, B2 =>
                           n40526, C1 => n40518, C2 => n38895, ZN => n9671);
   U33253 : OAI222_X1 port map( A1 => n40769, A2 => n40532, B1 => n41153, B2 =>
                           n40525, C1 => n40518, C2 => n38896, ZN => n9670);
   U33254 : OAI222_X1 port map( A1 => n40775, A2 => n40532, B1 => n41159, B2 =>
                           n40525, C1 => n40518, C2 => n38897, ZN => n9669);
   U33255 : OAI222_X1 port map( A1 => n40781, A2 => n40532, B1 => n41165, B2 =>
                           n40525, C1 => n40518, C2 => n38898, ZN => n9668);
   U33256 : OAI222_X1 port map( A1 => n40787, A2 => n40532, B1 => n41171, B2 =>
                           n40525, C1 => n40518, C2 => n38899, ZN => n9667);
   U33257 : OAI222_X1 port map( A1 => n40793, A2 => n40532, B1 => n41177, B2 =>
                           n40525, C1 => n40518, C2 => n38900, ZN => n9666);
   U33258 : OAI222_X1 port map( A1 => n40799, A2 => n40532, B1 => n41183, B2 =>
                           n40525, C1 => n40518, C2 => n38901, ZN => n9665);
   U33259 : OAI222_X1 port map( A1 => n40805, A2 => n40532, B1 => n41189, B2 =>
                           n40525, C1 => n40518, C2 => n38902, ZN => n9664);
   U33260 : OAI222_X1 port map( A1 => n40811, A2 => n40532, B1 => n41195, B2 =>
                           n40525, C1 => n40518, C2 => n38903, ZN => n9663);
   U33261 : OAI222_X1 port map( A1 => n40817, A2 => n40532, B1 => n41201, B2 =>
                           n40525, C1 => n40519, C2 => n38904, ZN => n9662);
   U33262 : OAI222_X1 port map( A1 => n40823, A2 => n40532, B1 => n41207, B2 =>
                           n40525, C1 => n40519, C2 => n38905, ZN => n9661);
   U33263 : OAI222_X1 port map( A1 => n40829, A2 => n40532, B1 => n41213, B2 =>
                           n40525, C1 => n40519, C2 => n38906, ZN => n9660);
   U33264 : OAI222_X1 port map( A1 => n40835, A2 => n40532, B1 => n41219, B2 =>
                           n40525, C1 => n40519, C2 => n38907, ZN => n9659);
   U33265 : OAI222_X1 port map( A1 => n40841, A2 => n40531, B1 => n41225, B2 =>
                           n40524, C1 => n40519, C2 => n38908, ZN => n9658);
   U33266 : OAI222_X1 port map( A1 => n40847, A2 => n40531, B1 => n41231, B2 =>
                           n40524, C1 => n40519, C2 => n38909, ZN => n9657);
   U33267 : OAI222_X1 port map( A1 => n40853, A2 => n40531, B1 => n41237, B2 =>
                           n40524, C1 => n40519, C2 => n38910, ZN => n9656);
   U33268 : OAI222_X1 port map( A1 => n40859, A2 => n40531, B1 => n41243, B2 =>
                           n40524, C1 => n40519, C2 => n38911, ZN => n9655);
   U33269 : OAI222_X1 port map( A1 => n40865, A2 => n40531, B1 => n41249, B2 =>
                           n40524, C1 => n40519, C2 => n38912, ZN => n9654);
   U33270 : OAI222_X1 port map( A1 => n40871, A2 => n40531, B1 => n41255, B2 =>
                           n40524, C1 => n40519, C2 => n38913, ZN => n9653);
   U33271 : OAI222_X1 port map( A1 => n40877, A2 => n40531, B1 => n41261, B2 =>
                           n40524, C1 => n40519, C2 => n38914, ZN => n9652);
   U33272 : OAI222_X1 port map( A1 => n40883, A2 => n40531, B1 => n41267, B2 =>
                           n40524, C1 => n40519, C2 => n38915, ZN => n9651);
   U33273 : OAI222_X1 port map( A1 => n40889, A2 => n40531, B1 => n41273, B2 =>
                           n40524, C1 => n40520, C2 => n38916, ZN => n9650);
   U33274 : OAI222_X1 port map( A1 => n40895, A2 => n40531, B1 => n41279, B2 =>
                           n40524, C1 => n40520, C2 => n38917, ZN => n9649);
   U33275 : OAI222_X1 port map( A1 => n40901, A2 => n40531, B1 => n41285, B2 =>
                           n40524, C1 => n40520, C2 => n38918, ZN => n9648);
   U33276 : OAI222_X1 port map( A1 => n40907, A2 => n40531, B1 => n41291, B2 =>
                           n40524, C1 => n40520, C2 => n38919, ZN => n9647);
   U33277 : OAI222_X1 port map( A1 => n40912, A2 => n40510, B1 => n41296, B2 =>
                           n40503, C1 => n40500, C2 => n38987, ZN => n9582);
   U33278 : OAI222_X1 port map( A1 => n40918, A2 => n40510, B1 => n41302, B2 =>
                           n40503, C1 => n40500, C2 => n38988, ZN => n9581);
   U33279 : OAI222_X1 port map( A1 => n40924, A2 => n40510, B1 => n41308, B2 =>
                           n40503, C1 => n40500, C2 => n38989, ZN => n9580);
   U33280 : OAI222_X1 port map( A1 => n40930, A2 => n40510, B1 => n41314, B2 =>
                           n40503, C1 => n40500, C2 => n38990, ZN => n9579);
   U33281 : OAI222_X1 port map( A1 => n40936, A2 => n40510, B1 => n41320, B2 =>
                           n40503, C1 => n40500, C2 => n38991, ZN => n9578);
   U33282 : OAI222_X1 port map( A1 => n40942, A2 => n40510, B1 => n41326, B2 =>
                           n40503, C1 => n40500, C2 => n38992, ZN => n9577);
   U33283 : OAI222_X1 port map( A1 => n40948, A2 => n40510, B1 => n41332, B2 =>
                           n40503, C1 => n40500, C2 => n38993, ZN => n9576);
   U33284 : OAI222_X1 port map( A1 => n40960, A2 => n40510, B1 => n41344, B2 =>
                           n40503, C1 => n40500, C2 => n38994, ZN => n9574);
   U33285 : OAI222_X1 port map( A1 => n40624, A2 => n40514, B1 => n41008, B2 =>
                           n40507, C1 => n40496, C2 => n38995, ZN => n9630);
   U33286 : OAI222_X1 port map( A1 => n40630, A2 => n40514, B1 => n41014, B2 =>
                           n40507, C1 => n40496, C2 => n38996, ZN => n9629);
   U33287 : OAI222_X1 port map( A1 => n40636, A2 => n40514, B1 => n41020, B2 =>
                           n40507, C1 => n40496, C2 => n38997, ZN => n9628);
   U33288 : OAI222_X1 port map( A1 => n40642, A2 => n40514, B1 => n41026, B2 =>
                           n40507, C1 => n40496, C2 => n38998, ZN => n9627);
   U33289 : OAI222_X1 port map( A1 => n40648, A2 => n40514, B1 => n41032, B2 =>
                           n40507, C1 => n40496, C2 => n38999, ZN => n9626);
   U33290 : OAI222_X1 port map( A1 => n40654, A2 => n40514, B1 => n41038, B2 =>
                           n40507, C1 => n40496, C2 => n39000, ZN => n9625);
   U33291 : OAI222_X1 port map( A1 => n40660, A2 => n40514, B1 => n41044, B2 =>
                           n40507, C1 => n40496, C2 => n39001, ZN => n9624);
   U33292 : OAI222_X1 port map( A1 => n40666, A2 => n40514, B1 => n41050, B2 =>
                           n40507, C1 => n40496, C2 => n39002, ZN => n9623);
   U33293 : OAI222_X1 port map( A1 => n40672, A2 => n40514, B1 => n41056, B2 =>
                           n40507, C1 => n40497, C2 => n39003, ZN => n9622);
   U33294 : OAI222_X1 port map( A1 => n40678, A2 => n40514, B1 => n41062, B2 =>
                           n40507, C1 => n40497, C2 => n39004, ZN => n9621);
   U33295 : OAI222_X1 port map( A1 => n40684, A2 => n40514, B1 => n41068, B2 =>
                           n40507, C1 => n40497, C2 => n39005, ZN => n9620);
   U33296 : OAI222_X1 port map( A1 => n40690, A2 => n40514, B1 => n41074, B2 =>
                           n40507, C1 => n40498, C2 => n39006, ZN => n9619);
   U33297 : OAI222_X1 port map( A1 => n40696, A2 => n40513, B1 => n41080, B2 =>
                           n40506, C1 => n40497, C2 => n39007, ZN => n9618);
   U33298 : OAI222_X1 port map( A1 => n40702, A2 => n40513, B1 => n41086, B2 =>
                           n40506, C1 => n40497, C2 => n39008, ZN => n9617);
   U33299 : OAI222_X1 port map( A1 => n40708, A2 => n40513, B1 => n41092, B2 =>
                           n40506, C1 => n40497, C2 => n39009, ZN => n9616);
   U33300 : OAI222_X1 port map( A1 => n40714, A2 => n40513, B1 => n41098, B2 =>
                           n40506, C1 => n40497, C2 => n39010, ZN => n9615);
   U33301 : OAI222_X1 port map( A1 => n40720, A2 => n40513, B1 => n41104, B2 =>
                           n40506, C1 => n40497, C2 => n39011, ZN => n9614);
   U33302 : OAI222_X1 port map( A1 => n40726, A2 => n40513, B1 => n41110, B2 =>
                           n40506, C1 => n40497, C2 => n39012, ZN => n9613);
   U33303 : OAI222_X1 port map( A1 => n40732, A2 => n40513, B1 => n41116, B2 =>
                           n40506, C1 => n40497, C2 => n39013, ZN => n9612);
   U33304 : OAI222_X1 port map( A1 => n40738, A2 => n40513, B1 => n41122, B2 =>
                           n40506, C1 => n40497, C2 => n39014, ZN => n9611);
   U33305 : OAI222_X1 port map( A1 => n40744, A2 => n40513, B1 => n41128, B2 =>
                           n40506, C1 => n40497, C2 => n39015, ZN => n9610);
   U33306 : OAI222_X1 port map( A1 => n40750, A2 => n40513, B1 => n41134, B2 =>
                           n40506, C1 => n40498, C2 => n39016, ZN => n9609);
   U33307 : OAI222_X1 port map( A1 => n40756, A2 => n40513, B1 => n41140, B2 =>
                           n40506, C1 => n40498, C2 => n39017, ZN => n9608);
   U33308 : OAI222_X1 port map( A1 => n40762, A2 => n40513, B1 => n41146, B2 =>
                           n40506, C1 => n40498, C2 => n39018, ZN => n9607);
   U33309 : OAI222_X1 port map( A1 => n40768, A2 => n40512, B1 => n41152, B2 =>
                           n40505, C1 => n40498, C2 => n39019, ZN => n9606);
   U33310 : OAI222_X1 port map( A1 => n40774, A2 => n40512, B1 => n41158, B2 =>
                           n40505, C1 => n40498, C2 => n39020, ZN => n9605);
   U33311 : OAI222_X1 port map( A1 => n40780, A2 => n40512, B1 => n41164, B2 =>
                           n40505, C1 => n40498, C2 => n39021, ZN => n9604);
   U33312 : OAI222_X1 port map( A1 => n40786, A2 => n40512, B1 => n41170, B2 =>
                           n40505, C1 => n40498, C2 => n39022, ZN => n9603);
   U33313 : OAI222_X1 port map( A1 => n40792, A2 => n40512, B1 => n41176, B2 =>
                           n40505, C1 => n40498, C2 => n39023, ZN => n9602);
   U33314 : OAI222_X1 port map( A1 => n40798, A2 => n40512, B1 => n41182, B2 =>
                           n40505, C1 => n40498, C2 => n39024, ZN => n9601);
   U33315 : OAI222_X1 port map( A1 => n40804, A2 => n40512, B1 => n41188, B2 =>
                           n40505, C1 => n40498, C2 => n39025, ZN => n9600);
   U33316 : OAI222_X1 port map( A1 => n40810, A2 => n40512, B1 => n41194, B2 =>
                           n40505, C1 => n40498, C2 => n39026, ZN => n9599);
   U33317 : OAI222_X1 port map( A1 => n40816, A2 => n40512, B1 => n41200, B2 =>
                           n40505, C1 => n40499, C2 => n39027, ZN => n9598);
   U33318 : OAI222_X1 port map( A1 => n40822, A2 => n40512, B1 => n41206, B2 =>
                           n40505, C1 => n40499, C2 => n39028, ZN => n9597);
   U33319 : OAI222_X1 port map( A1 => n40828, A2 => n40512, B1 => n41212, B2 =>
                           n40505, C1 => n40499, C2 => n39029, ZN => n9596);
   U33320 : OAI222_X1 port map( A1 => n40834, A2 => n40512, B1 => n41218, B2 =>
                           n40505, C1 => n40499, C2 => n39030, ZN => n9595);
   U33321 : OAI222_X1 port map( A1 => n40840, A2 => n40511, B1 => n41224, B2 =>
                           n40504, C1 => n40499, C2 => n39031, ZN => n9594);
   U33322 : OAI222_X1 port map( A1 => n40846, A2 => n40511, B1 => n41230, B2 =>
                           n40504, C1 => n40499, C2 => n39032, ZN => n9593);
   U33323 : OAI222_X1 port map( A1 => n40852, A2 => n40511, B1 => n41236, B2 =>
                           n40504, C1 => n40499, C2 => n39033, ZN => n9592);
   U33324 : OAI222_X1 port map( A1 => n40858, A2 => n40511, B1 => n41242, B2 =>
                           n40504, C1 => n40499, C2 => n39034, ZN => n9591);
   U33325 : OAI222_X1 port map( A1 => n40864, A2 => n40511, B1 => n41248, B2 =>
                           n40504, C1 => n40499, C2 => n39035, ZN => n9590);
   U33326 : OAI222_X1 port map( A1 => n40870, A2 => n40511, B1 => n41254, B2 =>
                           n40504, C1 => n40499, C2 => n39036, ZN => n9589);
   U33327 : OAI222_X1 port map( A1 => n40876, A2 => n40511, B1 => n41260, B2 =>
                           n40504, C1 => n40499, C2 => n39037, ZN => n9588);
   U33328 : OAI222_X1 port map( A1 => n40882, A2 => n40511, B1 => n41266, B2 =>
                           n40504, C1 => n40499, C2 => n39038, ZN => n9587);
   U33329 : OAI222_X1 port map( A1 => n40888, A2 => n40511, B1 => n41272, B2 =>
                           n40504, C1 => n40500, C2 => n39039, ZN => n9586);
   U33330 : OAI222_X1 port map( A1 => n40894, A2 => n40511, B1 => n41278, B2 =>
                           n40504, C1 => n40500, C2 => n39040, ZN => n9585);
   U33331 : OAI222_X1 port map( A1 => n40900, A2 => n40511, B1 => n41284, B2 =>
                           n40504, C1 => n40500, C2 => n39041, ZN => n9584);
   U33332 : OAI222_X1 port map( A1 => n40906, A2 => n40511, B1 => n41290, B2 =>
                           n40504, C1 => n40500, C2 => n39042, ZN => n9583);
   U33333 : OAI222_X1 port map( A1 => n40601, A2 => n40535, B1 => n40985, B2 =>
                           n40528, C1 => n40516, C2 => n38920, ZN => n9698);
   U33334 : OAI222_X1 port map( A1 => n40607, A2 => n40535, B1 => n40991, B2 =>
                           n40528, C1 => n40516, C2 => n38921, ZN => n9697);
   U33335 : OAI222_X1 port map( A1 => n40613, A2 => n40535, B1 => n40997, B2 =>
                           n40528, C1 => n40516, C2 => n38922, ZN => n9696);
   U33336 : OAI222_X1 port map( A1 => n40619, A2 => n40535, B1 => n41003, B2 =>
                           n40528, C1 => n40516, C2 => n38923, ZN => n9695);
   U33337 : OAI222_X1 port map( A1 => n40600, A2 => n40515, B1 => n40984, B2 =>
                           n40508, C1 => n40496, C2 => n39043, ZN => n9634);
   U33338 : OAI222_X1 port map( A1 => n40606, A2 => n40515, B1 => n40990, B2 =>
                           n40508, C1 => n40496, C2 => n39044, ZN => n9633);
   U33339 : OAI222_X1 port map( A1 => n40612, A2 => n40515, B1 => n40996, B2 =>
                           n40508, C1 => n40496, C2 => n39045, ZN => n9632);
   U33340 : OAI222_X1 port map( A1 => n40618, A2 => n40515, B1 => n41002, B2 =>
                           n40508, C1 => n40496, C2 => n39046, ZN => n9631);
   U33341 : AOI221_X1 port map( B1 => n39222, B2 => n29415, C1 => n39216, C2 =>
                           n29479, A => n37018, ZN => n37013);
   U33342 : OAI222_X1 port map( A1 => n31675, A2 => n39210, B1 => n31739, B2 =>
                           n39204, C1 => n31611, C2 => n39198, ZN => n37018);
   U33343 : AOI221_X1 port map( B1 => n39223, B2 => n29414, C1 => n39217, C2 =>
                           n29478, A => n36999, ZN => n36994);
   U33344 : OAI222_X1 port map( A1 => n31674, A2 => n39211, B1 => n31738, B2 =>
                           n39205, C1 => n31610, C2 => n39199, ZN => n36999);
   U33345 : AOI221_X1 port map( B1 => n39223, B2 => n29413, C1 => n39217, C2 =>
                           n29477, A => n36980, ZN => n36975);
   U33346 : OAI222_X1 port map( A1 => n31673, A2 => n39211, B1 => n31737, B2 =>
                           n39205, C1 => n31609, C2 => n39199, ZN => n36980);
   U33347 : AOI221_X1 port map( B1 => n39223, B2 => n29412, C1 => n39217, C2 =>
                           n29476, A => n36961, ZN => n36956);
   U33348 : OAI222_X1 port map( A1 => n31672, A2 => n39211, B1 => n31736, B2 =>
                           n39205, C1 => n31608, C2 => n39199, ZN => n36961);
   U33349 : AOI221_X1 port map( B1 => n39223, B2 => n29411, C1 => n39217, C2 =>
                           n29475, A => n36942, ZN => n36937);
   U33350 : OAI222_X1 port map( A1 => n31671, A2 => n39211, B1 => n31735, B2 =>
                           n39205, C1 => n31607, C2 => n39199, ZN => n36942);
   U33351 : AOI221_X1 port map( B1 => n39223, B2 => n29410, C1 => n39217, C2 =>
                           n29474, A => n36923, ZN => n36918);
   U33352 : OAI222_X1 port map( A1 => n31670, A2 => n39211, B1 => n31734, B2 =>
                           n39205, C1 => n31606, C2 => n39199, ZN => n36923);
   U33353 : AOI221_X1 port map( B1 => n39223, B2 => n29409, C1 => n39217, C2 =>
                           n29473, A => n36904, ZN => n36899);
   U33354 : OAI222_X1 port map( A1 => n31669, A2 => n39211, B1 => n31733, B2 =>
                           n39205, C1 => n31605, C2 => n39199, ZN => n36904);
   U33355 : AOI221_X1 port map( B1 => n39223, B2 => n29408, C1 => n39217, C2 =>
                           n29472, A => n36885, ZN => n36880);
   U33356 : OAI222_X1 port map( A1 => n31668, A2 => n39211, B1 => n31732, B2 =>
                           n39205, C1 => n31604, C2 => n39199, ZN => n36885);
   U33357 : AOI221_X1 port map( B1 => n39223, B2 => n29407, C1 => n39217, C2 =>
                           n29471, A => n36866, ZN => n36861);
   U33358 : OAI222_X1 port map( A1 => n31667, A2 => n39211, B1 => n31731, B2 =>
                           n39205, C1 => n31603, C2 => n39199, ZN => n36866);
   U33359 : AOI221_X1 port map( B1 => n39223, B2 => n29406, C1 => n39217, C2 =>
                           n29470, A => n36847, ZN => n36842);
   U33360 : OAI222_X1 port map( A1 => n31666, A2 => n39211, B1 => n31730, B2 =>
                           n39205, C1 => n31602, C2 => n39199, ZN => n36847);
   U33361 : AOI221_X1 port map( B1 => n39223, B2 => n29405, C1 => n39217, C2 =>
                           n29469, A => n36828, ZN => n36823);
   U33362 : OAI222_X1 port map( A1 => n31665, A2 => n39211, B1 => n31729, B2 =>
                           n39205, C1 => n31601, C2 => n39199, ZN => n36828);
   U33363 : AOI221_X1 port map( B1 => n39223, B2 => n29404, C1 => n39217, C2 =>
                           n29468, A => n36809, ZN => n36804);
   U33364 : OAI222_X1 port map( A1 => n31664, A2 => n39211, B1 => n31728, B2 =>
                           n39205, C1 => n31600, C2 => n39199, ZN => n36809);
   U33365 : AOI221_X1 port map( B1 => n39223, B2 => n29403, C1 => n39217, C2 =>
                           n29467, A => n36790, ZN => n36785);
   U33366 : OAI222_X1 port map( A1 => n31663, A2 => n39211, B1 => n31727, B2 =>
                           n39205, C1 => n31599, C2 => n39199, ZN => n36790);
   U33367 : AOI221_X1 port map( B1 => n39224, B2 => n29402, C1 => n39218, C2 =>
                           n29466, A => n36771, ZN => n36766);
   U33368 : OAI222_X1 port map( A1 => n31662, A2 => n39212, B1 => n31726, B2 =>
                           n39206, C1 => n31598, C2 => n39200, ZN => n36771);
   U33369 : AOI221_X1 port map( B1 => n39224, B2 => n29401, C1 => n39218, C2 =>
                           n29465, A => n36752, ZN => n36747);
   U33370 : OAI222_X1 port map( A1 => n31661, A2 => n39212, B1 => n31725, B2 =>
                           n39206, C1 => n31597, C2 => n39200, ZN => n36752);
   U33371 : AOI221_X1 port map( B1 => n39224, B2 => n29400, C1 => n39218, C2 =>
                           n29464, A => n36733, ZN => n36728);
   U33372 : OAI222_X1 port map( A1 => n31660, A2 => n39212, B1 => n31724, B2 =>
                           n39206, C1 => n31596, C2 => n39200, ZN => n36733);
   U33373 : AOI221_X1 port map( B1 => n39224, B2 => n29399, C1 => n39218, C2 =>
                           n29463, A => n36714, ZN => n36709);
   U33374 : OAI222_X1 port map( A1 => n31659, A2 => n39212, B1 => n31723, B2 =>
                           n39206, C1 => n31595, C2 => n39200, ZN => n36714);
   U33375 : AOI221_X1 port map( B1 => n39224, B2 => n29398, C1 => n39218, C2 =>
                           n29462, A => n36695, ZN => n36690);
   U33376 : OAI222_X1 port map( A1 => n31658, A2 => n39212, B1 => n31722, B2 =>
                           n39206, C1 => n31594, C2 => n39200, ZN => n36695);
   U33377 : AOI221_X1 port map( B1 => n39224, B2 => n29397, C1 => n39218, C2 =>
                           n29461, A => n36676, ZN => n36671);
   U33378 : OAI222_X1 port map( A1 => n31657, A2 => n39212, B1 => n31721, B2 =>
                           n39206, C1 => n31593, C2 => n39200, ZN => n36676);
   U33379 : AOI221_X1 port map( B1 => n39224, B2 => n29396, C1 => n39218, C2 =>
                           n29460, A => n36657, ZN => n36652);
   U33380 : OAI222_X1 port map( A1 => n31656, A2 => n39212, B1 => n31720, B2 =>
                           n39206, C1 => n31592, C2 => n39200, ZN => n36657);
   U33381 : AOI221_X1 port map( B1 => n39224, B2 => n29395, C1 => n39218, C2 =>
                           n29459, A => n36638, ZN => n36633);
   U33382 : OAI222_X1 port map( A1 => n31655, A2 => n39212, B1 => n31719, B2 =>
                           n39206, C1 => n31591, C2 => n39200, ZN => n36638);
   U33383 : AOI221_X1 port map( B1 => n39224, B2 => n29394, C1 => n39218, C2 =>
                           n29458, A => n36619, ZN => n36614);
   U33384 : OAI222_X1 port map( A1 => n31654, A2 => n39212, B1 => n31718, B2 =>
                           n39206, C1 => n31590, C2 => n39200, ZN => n36619);
   U33385 : AOI221_X1 port map( B1 => n39224, B2 => n29393, C1 => n39218, C2 =>
                           n29457, A => n36600, ZN => n36595);
   U33386 : OAI222_X1 port map( A1 => n31653, A2 => n39212, B1 => n31717, B2 =>
                           n39206, C1 => n31589, C2 => n39200, ZN => n36600);
   U33387 : AOI221_X1 port map( B1 => n39224, B2 => n29392, C1 => n39218, C2 =>
                           n29456, A => n36581, ZN => n36576);
   U33388 : OAI222_X1 port map( A1 => n31652, A2 => n39212, B1 => n31716, B2 =>
                           n39206, C1 => n31588, C2 => n39200, ZN => n36581);
   U33389 : AOI221_X1 port map( B1 => n39224, B2 => n29391, C1 => n39218, C2 =>
                           n29455, A => n36562, ZN => n36557);
   U33390 : OAI222_X1 port map( A1 => n31651, A2 => n39212, B1 => n31715, B2 =>
                           n39206, C1 => n31587, C2 => n39200, ZN => n36562);
   U33391 : AOI221_X1 port map( B1 => n39225, B2 => n29390, C1 => n39219, C2 =>
                           n29454, A => n36543, ZN => n36538);
   U33392 : OAI222_X1 port map( A1 => n31650, A2 => n39213, B1 => n31714, B2 =>
                           n39207, C1 => n31586, C2 => n39201, ZN => n36543);
   U33393 : AOI221_X1 port map( B1 => n39225, B2 => n29389, C1 => n39219, C2 =>
                           n29453, A => n36524, ZN => n36519);
   U33394 : OAI222_X1 port map( A1 => n31649, A2 => n39213, B1 => n31713, B2 =>
                           n39207, C1 => n31585, C2 => n39201, ZN => n36524);
   U33395 : AOI221_X1 port map( B1 => n39225, B2 => n29388, C1 => n39219, C2 =>
                           n29452, A => n36505, ZN => n36500);
   U33396 : OAI222_X1 port map( A1 => n31648, A2 => n39213, B1 => n31712, B2 =>
                           n39207, C1 => n31584, C2 => n39201, ZN => n36505);
   U33397 : AOI221_X1 port map( B1 => n39225, B2 => n29387, C1 => n39219, C2 =>
                           n29451, A => n36486, ZN => n36481);
   U33398 : OAI222_X1 port map( A1 => n31647, A2 => n39213, B1 => n31711, B2 =>
                           n39207, C1 => n31583, C2 => n39201, ZN => n36486);
   U33399 : AOI221_X1 port map( B1 => n39225, B2 => n29386, C1 => n39219, C2 =>
                           n29450, A => n36467, ZN => n36462);
   U33400 : OAI222_X1 port map( A1 => n31646, A2 => n39213, B1 => n31710, B2 =>
                           n39207, C1 => n31582, C2 => n39201, ZN => n36467);
   U33401 : AOI221_X1 port map( B1 => n39225, B2 => n29385, C1 => n39219, C2 =>
                           n29449, A => n36448, ZN => n36443);
   U33402 : OAI222_X1 port map( A1 => n31645, A2 => n39213, B1 => n31709, B2 =>
                           n39207, C1 => n31581, C2 => n39201, ZN => n36448);
   U33403 : AOI221_X1 port map( B1 => n39225, B2 => n29384, C1 => n39219, C2 =>
                           n29448, A => n36429, ZN => n36424);
   U33404 : OAI222_X1 port map( A1 => n31644, A2 => n39213, B1 => n31708, B2 =>
                           n39207, C1 => n31580, C2 => n39201, ZN => n36429);
   U33405 : AOI221_X1 port map( B1 => n39225, B2 => n29383, C1 => n39219, C2 =>
                           n29447, A => n36410, ZN => n36405);
   U33406 : OAI222_X1 port map( A1 => n31643, A2 => n39213, B1 => n31707, B2 =>
                           n39207, C1 => n31579, C2 => n39201, ZN => n36410);
   U33407 : AOI221_X1 port map( B1 => n39225, B2 => n29382, C1 => n39219, C2 =>
                           n29446, A => n36391, ZN => n36386);
   U33408 : OAI222_X1 port map( A1 => n31642, A2 => n39213, B1 => n31706, B2 =>
                           n39207, C1 => n31578, C2 => n39201, ZN => n36391);
   U33409 : AOI221_X1 port map( B1 => n39225, B2 => n29381, C1 => n39219, C2 =>
                           n29445, A => n36372, ZN => n36367);
   U33410 : OAI222_X1 port map( A1 => n31641, A2 => n39213, B1 => n31705, B2 =>
                           n39207, C1 => n31577, C2 => n39201, ZN => n36372);
   U33411 : AOI221_X1 port map( B1 => n39225, B2 => n29380, C1 => n39219, C2 =>
                           n29444, A => n36353, ZN => n36348);
   U33412 : OAI222_X1 port map( A1 => n31640, A2 => n39213, B1 => n31704, B2 =>
                           n39207, C1 => n31576, C2 => n39201, ZN => n36353);
   U33413 : AOI221_X1 port map( B1 => n39225, B2 => n29379, C1 => n39219, C2 =>
                           n29443, A => n36334, ZN => n36329);
   U33414 : OAI222_X1 port map( A1 => n31639, A2 => n39213, B1 => n31703, B2 =>
                           n39207, C1 => n31575, C2 => n39201, ZN => n36334);
   U33415 : AOI221_X1 port map( B1 => n39226, B2 => n29378, C1 => n39220, C2 =>
                           n29442, A => n36315, ZN => n36310);
   U33416 : OAI222_X1 port map( A1 => n31638, A2 => n39214, B1 => n31702, B2 =>
                           n39208, C1 => n31574, C2 => n39202, ZN => n36315);
   U33417 : AOI221_X1 port map( B1 => n39226, B2 => n29377, C1 => n39220, C2 =>
                           n29441, A => n36296, ZN => n36291);
   U33418 : OAI222_X1 port map( A1 => n31637, A2 => n39214, B1 => n31701, B2 =>
                           n39208, C1 => n31573, C2 => n39202, ZN => n36296);
   U33419 : AOI221_X1 port map( B1 => n39226, B2 => n29376, C1 => n39220, C2 =>
                           n29440, A => n36277, ZN => n36272);
   U33420 : OAI222_X1 port map( A1 => n31636, A2 => n39214, B1 => n31700, B2 =>
                           n39208, C1 => n31572, C2 => n39202, ZN => n36277);
   U33421 : AOI221_X1 port map( B1 => n39226, B2 => n29375, C1 => n39220, C2 =>
                           n29439, A => n36258, ZN => n36253);
   U33422 : OAI222_X1 port map( A1 => n31635, A2 => n39214, B1 => n31699, B2 =>
                           n39208, C1 => n31571, C2 => n39202, ZN => n36258);
   U33423 : AOI221_X1 port map( B1 => n39226, B2 => n29374, C1 => n39220, C2 =>
                           n29438, A => n36239, ZN => n36234);
   U33424 : OAI222_X1 port map( A1 => n31634, A2 => n39214, B1 => n31698, B2 =>
                           n39208, C1 => n31570, C2 => n39202, ZN => n36239);
   U33425 : AOI221_X1 port map( B1 => n39226, B2 => n29373, C1 => n39220, C2 =>
                           n29437, A => n36220, ZN => n36215);
   U33426 : OAI222_X1 port map( A1 => n31633, A2 => n39214, B1 => n31697, B2 =>
                           n39208, C1 => n31569, C2 => n39202, ZN => n36220);
   U33427 : AOI221_X1 port map( B1 => n39222, B2 => n29425, C1 => n39216, C2 =>
                           n29489, A => n37208, ZN => n37203);
   U33428 : OAI222_X1 port map( A1 => n31685, A2 => n39210, B1 => n31749, B2 =>
                           n39204, C1 => n31621, C2 => n39198, ZN => n37208);
   U33429 : AOI221_X1 port map( B1 => n39222, B2 => n29424, C1 => n39216, C2 =>
                           n29488, A => n37189, ZN => n37184);
   U33430 : OAI222_X1 port map( A1 => n31684, A2 => n39210, B1 => n31748, B2 =>
                           n39204, C1 => n31620, C2 => n39198, ZN => n37189);
   U33431 : AOI221_X1 port map( B1 => n39222, B2 => n29423, C1 => n39216, C2 =>
                           n29487, A => n37170, ZN => n37165);
   U33432 : OAI222_X1 port map( A1 => n31683, A2 => n39210, B1 => n31747, B2 =>
                           n39204, C1 => n31619, C2 => n39198, ZN => n37170);
   U33433 : AOI221_X1 port map( B1 => n39222, B2 => n29422, C1 => n39216, C2 =>
                           n29486, A => n37151, ZN => n37146);
   U33434 : OAI222_X1 port map( A1 => n31682, A2 => n39210, B1 => n31746, B2 =>
                           n39204, C1 => n31618, C2 => n39198, ZN => n37151);
   U33435 : AOI221_X1 port map( B1 => n39222, B2 => n29421, C1 => n39216, C2 =>
                           n29485, A => n37132, ZN => n37127);
   U33436 : OAI222_X1 port map( A1 => n31681, A2 => n39210, B1 => n31745, B2 =>
                           n39204, C1 => n31617, C2 => n39198, ZN => n37132);
   U33437 : AOI221_X1 port map( B1 => n39227, B2 => n29366, C1 => n39221, C2 =>
                           n29430, A => n36087, ZN => n36082);
   U33438 : OAI222_X1 port map( A1 => n31626, A2 => n39215, B1 => n31690, B2 =>
                           n39209, C1 => n31562, C2 => n39203, ZN => n36087);
   U33439 : AOI221_X1 port map( B1 => n39227, B2 => n29365, C1 => n39221, C2 =>
                           n29429, A => n36068, ZN => n36063);
   U33440 : OAI222_X1 port map( A1 => n31625, A2 => n39215, B1 => n31689, B2 =>
                           n39209, C1 => n31561, C2 => n39203, ZN => n36068);
   U33441 : AOI221_X1 port map( B1 => n39227, B2 => n29364, C1 => n39221, C2 =>
                           n29428, A => n36049, ZN => n36044);
   U33442 : OAI222_X1 port map( A1 => n31624, A2 => n39215, B1 => n31688, B2 =>
                           n39209, C1 => n31560, C2 => n39203, ZN => n36049);
   U33443 : AOI221_X1 port map( B1 => n39227, B2 => n29363, C1 => n39221, C2 =>
                           n29427, A => n36002, ZN => n35985);
   U33444 : OAI222_X1 port map( A1 => n31623, A2 => n39215, B1 => n31687, B2 =>
                           n39209, C1 => n31559, C2 => n39203, ZN => n36002);
   U33445 : AOI221_X1 port map( B1 => n39222, B2 => n29426, C1 => n39216, C2 =>
                           n29490, A => n37237, ZN => n37222);
   U33446 : OAI222_X1 port map( A1 => n31686, A2 => n39210, B1 => n31750, B2 =>
                           n39204, C1 => n31622, C2 => n39198, ZN => n37237);
   U33447 : AOI221_X1 port map( B1 => n39222, B2 => n29420, C1 => n39216, C2 =>
                           n29484, A => n37113, ZN => n37108);
   U33448 : OAI222_X1 port map( A1 => n31680, A2 => n39210, B1 => n31744, B2 =>
                           n39204, C1 => n31616, C2 => n39198, ZN => n37113);
   U33449 : AOI221_X1 port map( B1 => n39222, B2 => n29419, C1 => n39216, C2 =>
                           n29483, A => n37094, ZN => n37089);
   U33450 : OAI222_X1 port map( A1 => n31679, A2 => n39210, B1 => n31743, B2 =>
                           n39204, C1 => n31615, C2 => n39198, ZN => n37094);
   U33451 : AOI221_X1 port map( B1 => n39222, B2 => n29418, C1 => n39216, C2 =>
                           n29482, A => n37075, ZN => n37070);
   U33452 : OAI222_X1 port map( A1 => n31678, A2 => n39210, B1 => n31742, B2 =>
                           n39204, C1 => n31614, C2 => n39198, ZN => n37075);
   U33453 : AOI221_X1 port map( B1 => n39222, B2 => n29417, C1 => n39216, C2 =>
                           n29481, A => n37056, ZN => n37051);
   U33454 : OAI222_X1 port map( A1 => n31677, A2 => n39210, B1 => n31741, B2 =>
                           n39204, C1 => n31613, C2 => n39198, ZN => n37056);
   U33455 : AOI221_X1 port map( B1 => n39222, B2 => n29416, C1 => n39216, C2 =>
                           n29480, A => n37037, ZN => n37032);
   U33456 : OAI222_X1 port map( A1 => n31676, A2 => n39210, B1 => n31740, B2 =>
                           n39204, C1 => n31612, C2 => n39198, ZN => n37037);
   U33457 : AOI221_X1 port map( B1 => n39226, B2 => n29372, C1 => n39220, C2 =>
                           n29436, A => n36201, ZN => n36196);
   U33458 : OAI222_X1 port map( A1 => n31632, A2 => n39214, B1 => n31696, B2 =>
                           n39208, C1 => n31568, C2 => n39202, ZN => n36201);
   U33459 : AOI221_X1 port map( B1 => n39226, B2 => n29371, C1 => n39220, C2 =>
                           n29435, A => n36182, ZN => n36177);
   U33460 : OAI222_X1 port map( A1 => n31631, A2 => n39214, B1 => n31695, B2 =>
                           n39208, C1 => n31567, C2 => n39202, ZN => n36182);
   U33461 : AOI221_X1 port map( B1 => n39226, B2 => n29370, C1 => n39220, C2 =>
                           n29434, A => n36163, ZN => n36158);
   U33462 : OAI222_X1 port map( A1 => n31630, A2 => n39214, B1 => n31694, B2 =>
                           n39208, C1 => n31566, C2 => n39202, ZN => n36163);
   U33463 : AOI221_X1 port map( B1 => n39226, B2 => n29369, C1 => n39220, C2 =>
                           n29433, A => n36144, ZN => n36139);
   U33464 : OAI222_X1 port map( A1 => n31629, A2 => n39214, B1 => n31693, B2 =>
                           n39208, C1 => n31565, C2 => n39202, ZN => n36144);
   U33465 : AOI221_X1 port map( B1 => n39226, B2 => n29368, C1 => n39220, C2 =>
                           n29432, A => n36125, ZN => n36120);
   U33466 : OAI222_X1 port map( A1 => n31628, A2 => n39214, B1 => n31692, B2 =>
                           n39208, C1 => n31564, C2 => n39202, ZN => n36125);
   U33467 : AOI221_X1 port map( B1 => n39226, B2 => n29367, C1 => n39220, C2 =>
                           n29431, A => n36106, ZN => n36101);
   U33468 : OAI222_X1 port map( A1 => n31627, A2 => n39214, B1 => n31691, B2 =>
                           n39208, C1 => n31563, C2 => n39202, ZN => n36106);
   U33469 : AOI221_X1 port map( B1 => n39729, B2 => n29426, C1 => n39723, C2 =>
                           n29490, A => n33447, ZN => n33430);
   U33470 : OAI222_X1 port map( A1 => n31686, A2 => n39717, B1 => n31750, B2 =>
                           n39711, C1 => n31622, C2 => n39705, ZN => n33447);
   U33471 : AOI221_X1 port map( B1 => n39477, B2 => n29426, C1 => n39471, C2 =>
                           n29490, A => n34721, ZN => n34704);
   U33472 : OAI222_X1 port map( A1 => n31686, A2 => n39465, B1 => n31750, B2 =>
                           n39459, C1 => n31622, C2 => n39453, ZN => n34721);
   U33473 : AOI221_X1 port map( B1 => n39729, B2 => n29425, C1 => n39723, C2 =>
                           n29489, A => n33494, ZN => n33489);
   U33474 : OAI222_X1 port map( A1 => n31685, A2 => n39717, B1 => n31749, B2 =>
                           n39711, C1 => n31621, C2 => n39705, ZN => n33494);
   U33475 : AOI221_X1 port map( B1 => n39477, B2 => n29425, C1 => n39471, C2 =>
                           n29489, A => n34768, ZN => n34763);
   U33476 : OAI222_X1 port map( A1 => n31685, A2 => n39465, B1 => n31749, B2 =>
                           n39459, C1 => n31621, C2 => n39453, ZN => n34768);
   U33477 : AOI221_X1 port map( B1 => n39729, B2 => n29424, C1 => n39723, C2 =>
                           n29488, A => n33513, ZN => n33508);
   U33478 : OAI222_X1 port map( A1 => n31684, A2 => n39717, B1 => n31748, B2 =>
                           n39711, C1 => n31620, C2 => n39705, ZN => n33513);
   U33479 : AOI221_X1 port map( B1 => n39477, B2 => n29424, C1 => n39471, C2 =>
                           n29488, A => n34787, ZN => n34782);
   U33480 : OAI222_X1 port map( A1 => n31684, A2 => n39465, B1 => n31748, B2 =>
                           n39459, C1 => n31620, C2 => n39453, ZN => n34787);
   U33481 : AOI221_X1 port map( B1 => n39729, B2 => n29423, C1 => n39723, C2 =>
                           n29487, A => n33532, ZN => n33527);
   U33482 : OAI222_X1 port map( A1 => n31683, A2 => n39717, B1 => n31747, B2 =>
                           n39711, C1 => n31619, C2 => n39705, ZN => n33532);
   U33483 : AOI221_X1 port map( B1 => n39477, B2 => n29423, C1 => n39471, C2 =>
                           n29487, A => n34806, ZN => n34801);
   U33484 : OAI222_X1 port map( A1 => n31683, A2 => n39465, B1 => n31747, B2 =>
                           n39459, C1 => n31619, C2 => n39453, ZN => n34806);
   U33485 : AOI221_X1 port map( B1 => n39728, B2 => n29422, C1 => n39722, C2 =>
                           n29486, A => n33551, ZN => n33546);
   U33486 : OAI222_X1 port map( A1 => n31682, A2 => n39716, B1 => n31746, B2 =>
                           n39710, C1 => n31618, C2 => n39704, ZN => n33551);
   U33487 : AOI221_X1 port map( B1 => n39476, B2 => n29422, C1 => n39470, C2 =>
                           n29486, A => n34825, ZN => n34820);
   U33488 : OAI222_X1 port map( A1 => n31682, A2 => n39464, B1 => n31746, B2 =>
                           n39458, C1 => n31618, C2 => n39452, ZN => n34825);
   U33489 : AOI221_X1 port map( B1 => n39728, B2 => n29421, C1 => n39722, C2 =>
                           n29485, A => n33570, ZN => n33565);
   U33490 : OAI222_X1 port map( A1 => n31681, A2 => n39716, B1 => n31745, B2 =>
                           n39710, C1 => n31617, C2 => n39704, ZN => n33570);
   U33491 : AOI221_X1 port map( B1 => n39476, B2 => n29421, C1 => n39470, C2 =>
                           n29485, A => n34844, ZN => n34839);
   U33492 : OAI222_X1 port map( A1 => n31681, A2 => n39464, B1 => n31745, B2 =>
                           n39458, C1 => n31617, C2 => n39452, ZN => n34844);
   U33493 : AOI221_X1 port map( B1 => n39728, B2 => n29420, C1 => n39722, C2 =>
                           n29484, A => n33589, ZN => n33584);
   U33494 : OAI222_X1 port map( A1 => n31680, A2 => n39716, B1 => n31744, B2 =>
                           n39710, C1 => n31616, C2 => n39704, ZN => n33589);
   U33495 : AOI221_X1 port map( B1 => n39476, B2 => n29420, C1 => n39470, C2 =>
                           n29484, A => n34863, ZN => n34858);
   U33496 : OAI222_X1 port map( A1 => n31680, A2 => n39464, B1 => n31744, B2 =>
                           n39458, C1 => n31616, C2 => n39452, ZN => n34863);
   U33497 : AOI221_X1 port map( B1 => n39728, B2 => n29419, C1 => n39722, C2 =>
                           n29483, A => n33608, ZN => n33603);
   U33498 : OAI222_X1 port map( A1 => n31679, A2 => n39716, B1 => n31743, B2 =>
                           n39710, C1 => n31615, C2 => n39704, ZN => n33608);
   U33499 : AOI221_X1 port map( B1 => n39476, B2 => n29419, C1 => n39470, C2 =>
                           n29483, A => n34882, ZN => n34877);
   U33500 : OAI222_X1 port map( A1 => n31679, A2 => n39464, B1 => n31743, B2 =>
                           n39458, C1 => n31615, C2 => n39452, ZN => n34882);
   U33501 : AOI221_X1 port map( B1 => n39728, B2 => n29418, C1 => n39722, C2 =>
                           n29482, A => n33627, ZN => n33622);
   U33502 : OAI222_X1 port map( A1 => n31678, A2 => n39716, B1 => n31742, B2 =>
                           n39710, C1 => n31614, C2 => n39704, ZN => n33627);
   U33503 : AOI221_X1 port map( B1 => n39476, B2 => n29418, C1 => n39470, C2 =>
                           n29482, A => n34901, ZN => n34896);
   U33504 : OAI222_X1 port map( A1 => n31678, A2 => n39464, B1 => n31742, B2 =>
                           n39458, C1 => n31614, C2 => n39452, ZN => n34901);
   U33505 : AOI221_X1 port map( B1 => n39728, B2 => n29417, C1 => n39722, C2 =>
                           n29481, A => n33646, ZN => n33641);
   U33506 : OAI222_X1 port map( A1 => n31677, A2 => n39716, B1 => n31741, B2 =>
                           n39710, C1 => n31613, C2 => n39704, ZN => n33646);
   U33507 : AOI221_X1 port map( B1 => n39476, B2 => n29417, C1 => n39470, C2 =>
                           n29481, A => n34920, ZN => n34915);
   U33508 : OAI222_X1 port map( A1 => n31677, A2 => n39464, B1 => n31741, B2 =>
                           n39458, C1 => n31613, C2 => n39452, ZN => n34920);
   U33509 : AOI221_X1 port map( B1 => n39728, B2 => n29416, C1 => n39722, C2 =>
                           n29480, A => n33665, ZN => n33660);
   U33510 : OAI222_X1 port map( A1 => n31676, A2 => n39716, B1 => n31740, B2 =>
                           n39710, C1 => n31612, C2 => n39704, ZN => n33665);
   U33511 : AOI221_X1 port map( B1 => n39476, B2 => n29416, C1 => n39470, C2 =>
                           n29480, A => n34939, ZN => n34934);
   U33512 : OAI222_X1 port map( A1 => n31676, A2 => n39464, B1 => n31740, B2 =>
                           n39458, C1 => n31612, C2 => n39452, ZN => n34939);
   U33513 : AOI221_X1 port map( B1 => n39728, B2 => n29415, C1 => n39722, C2 =>
                           n29479, A => n33684, ZN => n33679);
   U33514 : OAI222_X1 port map( A1 => n31675, A2 => n39716, B1 => n31739, B2 =>
                           n39710, C1 => n31611, C2 => n39704, ZN => n33684);
   U33515 : AOI221_X1 port map( B1 => n39476, B2 => n29415, C1 => n39470, C2 =>
                           n29479, A => n34958, ZN => n34953);
   U33516 : OAI222_X1 port map( A1 => n31675, A2 => n39464, B1 => n31739, B2 =>
                           n39458, C1 => n31611, C2 => n39452, ZN => n34958);
   U33517 : AOI221_X1 port map( B1 => n39728, B2 => n29414, C1 => n39722, C2 =>
                           n29478, A => n33703, ZN => n33698);
   U33518 : OAI222_X1 port map( A1 => n31674, A2 => n39716, B1 => n31738, B2 =>
                           n39710, C1 => n31610, C2 => n39704, ZN => n33703);
   U33519 : AOI221_X1 port map( B1 => n39476, B2 => n29414, C1 => n39470, C2 =>
                           n29478, A => n34977, ZN => n34972);
   U33520 : OAI222_X1 port map( A1 => n31674, A2 => n39464, B1 => n31738, B2 =>
                           n39458, C1 => n31610, C2 => n39452, ZN => n34977);
   U33521 : AOI221_X1 port map( B1 => n39728, B2 => n29413, C1 => n39722, C2 =>
                           n29477, A => n33722, ZN => n33717);
   U33522 : OAI222_X1 port map( A1 => n31673, A2 => n39716, B1 => n31737, B2 =>
                           n39710, C1 => n31609, C2 => n39704, ZN => n33722);
   U33523 : AOI221_X1 port map( B1 => n39476, B2 => n29413, C1 => n39470, C2 =>
                           n29477, A => n34996, ZN => n34991);
   U33524 : OAI222_X1 port map( A1 => n31673, A2 => n39464, B1 => n31737, B2 =>
                           n39458, C1 => n31609, C2 => n39452, ZN => n34996);
   U33525 : AOI221_X1 port map( B1 => n39728, B2 => n29412, C1 => n39722, C2 =>
                           n29476, A => n33741, ZN => n33736);
   U33526 : OAI222_X1 port map( A1 => n31672, A2 => n39716, B1 => n31736, B2 =>
                           n39710, C1 => n31608, C2 => n39704, ZN => n33741);
   U33527 : AOI221_X1 port map( B1 => n39476, B2 => n29412, C1 => n39470, C2 =>
                           n29476, A => n35015, ZN => n35010);
   U33528 : OAI222_X1 port map( A1 => n31672, A2 => n39464, B1 => n31736, B2 =>
                           n39458, C1 => n31608, C2 => n39452, ZN => n35015);
   U33529 : AOI221_X1 port map( B1 => n39728, B2 => n29411, C1 => n39722, C2 =>
                           n29475, A => n33760, ZN => n33755);
   U33530 : OAI222_X1 port map( A1 => n31671, A2 => n39716, B1 => n31735, B2 =>
                           n39710, C1 => n31607, C2 => n39704, ZN => n33760);
   U33531 : AOI221_X1 port map( B1 => n39476, B2 => n29411, C1 => n39470, C2 =>
                           n29475, A => n35034, ZN => n35029);
   U33532 : OAI222_X1 port map( A1 => n31671, A2 => n39464, B1 => n31735, B2 =>
                           n39458, C1 => n31607, C2 => n39452, ZN => n35034);
   U33533 : AOI221_X1 port map( B1 => n39727, B2 => n29410, C1 => n39721, C2 =>
                           n29474, A => n33779, ZN => n33774);
   U33534 : OAI222_X1 port map( A1 => n31670, A2 => n39715, B1 => n31734, B2 =>
                           n39709, C1 => n31606, C2 => n39703, ZN => n33779);
   U33535 : AOI221_X1 port map( B1 => n39475, B2 => n29410, C1 => n39469, C2 =>
                           n29474, A => n35053, ZN => n35048);
   U33536 : OAI222_X1 port map( A1 => n31670, A2 => n39463, B1 => n31734, B2 =>
                           n39457, C1 => n31606, C2 => n39451, ZN => n35053);
   U33537 : AOI221_X1 port map( B1 => n39727, B2 => n29409, C1 => n39721, C2 =>
                           n29473, A => n33798, ZN => n33793);
   U33538 : OAI222_X1 port map( A1 => n31669, A2 => n39715, B1 => n31733, B2 =>
                           n39709, C1 => n31605, C2 => n39703, ZN => n33798);
   U33539 : AOI221_X1 port map( B1 => n39475, B2 => n29409, C1 => n39469, C2 =>
                           n29473, A => n35072, ZN => n35067);
   U33540 : OAI222_X1 port map( A1 => n31669, A2 => n39463, B1 => n31733, B2 =>
                           n39457, C1 => n31605, C2 => n39451, ZN => n35072);
   U33541 : AOI221_X1 port map( B1 => n39727, B2 => n29408, C1 => n39721, C2 =>
                           n29472, A => n33817, ZN => n33812);
   U33542 : OAI222_X1 port map( A1 => n31668, A2 => n39715, B1 => n31732, B2 =>
                           n39709, C1 => n31604, C2 => n39703, ZN => n33817);
   U33543 : AOI221_X1 port map( B1 => n39475, B2 => n29408, C1 => n39469, C2 =>
                           n29472, A => n35091, ZN => n35086);
   U33544 : OAI222_X1 port map( A1 => n31668, A2 => n39463, B1 => n31732, B2 =>
                           n39457, C1 => n31604, C2 => n39451, ZN => n35091);
   U33545 : AOI221_X1 port map( B1 => n39727, B2 => n29407, C1 => n39721, C2 =>
                           n29471, A => n33836, ZN => n33831);
   U33546 : OAI222_X1 port map( A1 => n31667, A2 => n39715, B1 => n31731, B2 =>
                           n39709, C1 => n31603, C2 => n39703, ZN => n33836);
   U33547 : AOI221_X1 port map( B1 => n39475, B2 => n29407, C1 => n39469, C2 =>
                           n29471, A => n35110, ZN => n35105);
   U33548 : OAI222_X1 port map( A1 => n31667, A2 => n39463, B1 => n31731, B2 =>
                           n39457, C1 => n31603, C2 => n39451, ZN => n35110);
   U33549 : AOI221_X1 port map( B1 => n39727, B2 => n29406, C1 => n39721, C2 =>
                           n29470, A => n33855, ZN => n33850);
   U33550 : OAI222_X1 port map( A1 => n31666, A2 => n39715, B1 => n31730, B2 =>
                           n39709, C1 => n31602, C2 => n39703, ZN => n33855);
   U33551 : AOI221_X1 port map( B1 => n39475, B2 => n29406, C1 => n39469, C2 =>
                           n29470, A => n35129, ZN => n35124);
   U33552 : OAI222_X1 port map( A1 => n31666, A2 => n39463, B1 => n31730, B2 =>
                           n39457, C1 => n31602, C2 => n39451, ZN => n35129);
   U33553 : AOI221_X1 port map( B1 => n39727, B2 => n29405, C1 => n39721, C2 =>
                           n29469, A => n33874, ZN => n33869);
   U33554 : OAI222_X1 port map( A1 => n31665, A2 => n39715, B1 => n31729, B2 =>
                           n39709, C1 => n31601, C2 => n39703, ZN => n33874);
   U33555 : AOI221_X1 port map( B1 => n39475, B2 => n29405, C1 => n39469, C2 =>
                           n29469, A => n35148, ZN => n35143);
   U33556 : OAI222_X1 port map( A1 => n31665, A2 => n39463, B1 => n31729, B2 =>
                           n39457, C1 => n31601, C2 => n39451, ZN => n35148);
   U33557 : AOI221_X1 port map( B1 => n39727, B2 => n29404, C1 => n39721, C2 =>
                           n29468, A => n33893, ZN => n33888);
   U33558 : OAI222_X1 port map( A1 => n31664, A2 => n39715, B1 => n31728, B2 =>
                           n39709, C1 => n31600, C2 => n39703, ZN => n33893);
   U33559 : AOI221_X1 port map( B1 => n39475, B2 => n29404, C1 => n39469, C2 =>
                           n29468, A => n35167, ZN => n35162);
   U33560 : OAI222_X1 port map( A1 => n31664, A2 => n39463, B1 => n31728, B2 =>
                           n39457, C1 => n31600, C2 => n39451, ZN => n35167);
   U33561 : AOI221_X1 port map( B1 => n39727, B2 => n29403, C1 => n39721, C2 =>
                           n29467, A => n33912, ZN => n33907);
   U33562 : OAI222_X1 port map( A1 => n31663, A2 => n39715, B1 => n31727, B2 =>
                           n39709, C1 => n31599, C2 => n39703, ZN => n33912);
   U33563 : AOI221_X1 port map( B1 => n39475, B2 => n29403, C1 => n39469, C2 =>
                           n29467, A => n35186, ZN => n35181);
   U33564 : OAI222_X1 port map( A1 => n31663, A2 => n39463, B1 => n31727, B2 =>
                           n39457, C1 => n31599, C2 => n39451, ZN => n35186);
   U33565 : AOI221_X1 port map( B1 => n39727, B2 => n29402, C1 => n39721, C2 =>
                           n29466, A => n33931, ZN => n33926);
   U33566 : OAI222_X1 port map( A1 => n31662, A2 => n39715, B1 => n31726, B2 =>
                           n39709, C1 => n31598, C2 => n39703, ZN => n33931);
   U33567 : AOI221_X1 port map( B1 => n39475, B2 => n29402, C1 => n39469, C2 =>
                           n29466, A => n35205, ZN => n35200);
   U33568 : OAI222_X1 port map( A1 => n31662, A2 => n39463, B1 => n31726, B2 =>
                           n39457, C1 => n31598, C2 => n39451, ZN => n35205);
   U33569 : AOI221_X1 port map( B1 => n39727, B2 => n29401, C1 => n39721, C2 =>
                           n29465, A => n33950, ZN => n33945);
   U33570 : OAI222_X1 port map( A1 => n31661, A2 => n39715, B1 => n31725, B2 =>
                           n39709, C1 => n31597, C2 => n39703, ZN => n33950);
   U33571 : AOI221_X1 port map( B1 => n39475, B2 => n29401, C1 => n39469, C2 =>
                           n29465, A => n35224, ZN => n35219);
   U33572 : OAI222_X1 port map( A1 => n31661, A2 => n39463, B1 => n31725, B2 =>
                           n39457, C1 => n31597, C2 => n39451, ZN => n35224);
   U33573 : AOI221_X1 port map( B1 => n39727, B2 => n29400, C1 => n39721, C2 =>
                           n29464, A => n33969, ZN => n33964);
   U33574 : OAI222_X1 port map( A1 => n31660, A2 => n39715, B1 => n31724, B2 =>
                           n39709, C1 => n31596, C2 => n39703, ZN => n33969);
   U33575 : AOI221_X1 port map( B1 => n39475, B2 => n29400, C1 => n39469, C2 =>
                           n29464, A => n35243, ZN => n35238);
   U33576 : OAI222_X1 port map( A1 => n31660, A2 => n39463, B1 => n31724, B2 =>
                           n39457, C1 => n31596, C2 => n39451, ZN => n35243);
   U33577 : AOI221_X1 port map( B1 => n39727, B2 => n29399, C1 => n39721, C2 =>
                           n29463, A => n33988, ZN => n33983);
   U33578 : OAI222_X1 port map( A1 => n31659, A2 => n39715, B1 => n31723, B2 =>
                           n39709, C1 => n31595, C2 => n39703, ZN => n33988);
   U33579 : AOI221_X1 port map( B1 => n39475, B2 => n29399, C1 => n39469, C2 =>
                           n29463, A => n35262, ZN => n35257);
   U33580 : OAI222_X1 port map( A1 => n31659, A2 => n39463, B1 => n31723, B2 =>
                           n39457, C1 => n31595, C2 => n39451, ZN => n35262);
   U33581 : AOI221_X1 port map( B1 => n39726, B2 => n29398, C1 => n39720, C2 =>
                           n29462, A => n34007, ZN => n34002);
   U33582 : OAI222_X1 port map( A1 => n31658, A2 => n39714, B1 => n31722, B2 =>
                           n39708, C1 => n31594, C2 => n39702, ZN => n34007);
   U33583 : AOI221_X1 port map( B1 => n39474, B2 => n29398, C1 => n39468, C2 =>
                           n29462, A => n35281, ZN => n35276);
   U33584 : OAI222_X1 port map( A1 => n31658, A2 => n39462, B1 => n31722, B2 =>
                           n39456, C1 => n31594, C2 => n39450, ZN => n35281);
   U33585 : AOI221_X1 port map( B1 => n39726, B2 => n29397, C1 => n39720, C2 =>
                           n29461, A => n34026, ZN => n34021);
   U33586 : OAI222_X1 port map( A1 => n31657, A2 => n39714, B1 => n31721, B2 =>
                           n39708, C1 => n31593, C2 => n39702, ZN => n34026);
   U33587 : AOI221_X1 port map( B1 => n39474, B2 => n29397, C1 => n39468, C2 =>
                           n29461, A => n35300, ZN => n35295);
   U33588 : OAI222_X1 port map( A1 => n31657, A2 => n39462, B1 => n31721, B2 =>
                           n39456, C1 => n31593, C2 => n39450, ZN => n35300);
   U33589 : AOI221_X1 port map( B1 => n39726, B2 => n29396, C1 => n39720, C2 =>
                           n29460, A => n34045, ZN => n34040);
   U33590 : OAI222_X1 port map( A1 => n31656, A2 => n39714, B1 => n31720, B2 =>
                           n39708, C1 => n31592, C2 => n39702, ZN => n34045);
   U33591 : AOI221_X1 port map( B1 => n39474, B2 => n29396, C1 => n39468, C2 =>
                           n29460, A => n35319, ZN => n35314);
   U33592 : OAI222_X1 port map( A1 => n31656, A2 => n39462, B1 => n31720, B2 =>
                           n39456, C1 => n31592, C2 => n39450, ZN => n35319);
   U33593 : AOI221_X1 port map( B1 => n39726, B2 => n29395, C1 => n39720, C2 =>
                           n29459, A => n34064, ZN => n34059);
   U33594 : OAI222_X1 port map( A1 => n31655, A2 => n39714, B1 => n31719, B2 =>
                           n39708, C1 => n31591, C2 => n39702, ZN => n34064);
   U33595 : AOI221_X1 port map( B1 => n39474, B2 => n29395, C1 => n39468, C2 =>
                           n29459, A => n35338, ZN => n35333);
   U33596 : OAI222_X1 port map( A1 => n31655, A2 => n39462, B1 => n31719, B2 =>
                           n39456, C1 => n31591, C2 => n39450, ZN => n35338);
   U33597 : AOI221_X1 port map( B1 => n39726, B2 => n29394, C1 => n39720, C2 =>
                           n29458, A => n34083, ZN => n34078);
   U33598 : OAI222_X1 port map( A1 => n31654, A2 => n39714, B1 => n31718, B2 =>
                           n39708, C1 => n31590, C2 => n39702, ZN => n34083);
   U33599 : AOI221_X1 port map( B1 => n39474, B2 => n29394, C1 => n39468, C2 =>
                           n29458, A => n35357, ZN => n35352);
   U33600 : OAI222_X1 port map( A1 => n31654, A2 => n39462, B1 => n31718, B2 =>
                           n39456, C1 => n31590, C2 => n39450, ZN => n35357);
   U33601 : AOI221_X1 port map( B1 => n39726, B2 => n29393, C1 => n39720, C2 =>
                           n29457, A => n34102, ZN => n34097);
   U33602 : OAI222_X1 port map( A1 => n31653, A2 => n39714, B1 => n31717, B2 =>
                           n39708, C1 => n31589, C2 => n39702, ZN => n34102);
   U33603 : AOI221_X1 port map( B1 => n39474, B2 => n29393, C1 => n39468, C2 =>
                           n29457, A => n35376, ZN => n35371);
   U33604 : OAI222_X1 port map( A1 => n31653, A2 => n39462, B1 => n31717, B2 =>
                           n39456, C1 => n31589, C2 => n39450, ZN => n35376);
   U33605 : AOI221_X1 port map( B1 => n39726, B2 => n29392, C1 => n39720, C2 =>
                           n29456, A => n34121, ZN => n34116);
   U33606 : OAI222_X1 port map( A1 => n31652, A2 => n39714, B1 => n31716, B2 =>
                           n39708, C1 => n31588, C2 => n39702, ZN => n34121);
   U33607 : AOI221_X1 port map( B1 => n39474, B2 => n29392, C1 => n39468, C2 =>
                           n29456, A => n35395, ZN => n35390);
   U33608 : OAI222_X1 port map( A1 => n31652, A2 => n39462, B1 => n31716, B2 =>
                           n39456, C1 => n31588, C2 => n39450, ZN => n35395);
   U33609 : AOI221_X1 port map( B1 => n39726, B2 => n29391, C1 => n39720, C2 =>
                           n29455, A => n34140, ZN => n34135);
   U33610 : OAI222_X1 port map( A1 => n31651, A2 => n39714, B1 => n31715, B2 =>
                           n39708, C1 => n31587, C2 => n39702, ZN => n34140);
   U33611 : AOI221_X1 port map( B1 => n39474, B2 => n29391, C1 => n39468, C2 =>
                           n29455, A => n35414, ZN => n35409);
   U33612 : OAI222_X1 port map( A1 => n31651, A2 => n39462, B1 => n31715, B2 =>
                           n39456, C1 => n31587, C2 => n39450, ZN => n35414);
   U33613 : AOI221_X1 port map( B1 => n39726, B2 => n29390, C1 => n39720, C2 =>
                           n29454, A => n34159, ZN => n34154);
   U33614 : OAI222_X1 port map( A1 => n31650, A2 => n39714, B1 => n31714, B2 =>
                           n39708, C1 => n31586, C2 => n39702, ZN => n34159);
   U33615 : AOI221_X1 port map( B1 => n39474, B2 => n29390, C1 => n39468, C2 =>
                           n29454, A => n35433, ZN => n35428);
   U33616 : OAI222_X1 port map( A1 => n31650, A2 => n39462, B1 => n31714, B2 =>
                           n39456, C1 => n31586, C2 => n39450, ZN => n35433);
   U33617 : AOI221_X1 port map( B1 => n39726, B2 => n29389, C1 => n39720, C2 =>
                           n29453, A => n34178, ZN => n34173);
   U33618 : OAI222_X1 port map( A1 => n31649, A2 => n39714, B1 => n31713, B2 =>
                           n39708, C1 => n31585, C2 => n39702, ZN => n34178);
   U33619 : AOI221_X1 port map( B1 => n39474, B2 => n29389, C1 => n39468, C2 =>
                           n29453, A => n35452, ZN => n35447);
   U33620 : OAI222_X1 port map( A1 => n31649, A2 => n39462, B1 => n31713, B2 =>
                           n39456, C1 => n31585, C2 => n39450, ZN => n35452);
   U33621 : AOI221_X1 port map( B1 => n39726, B2 => n29388, C1 => n39720, C2 =>
                           n29452, A => n34197, ZN => n34192);
   U33622 : OAI222_X1 port map( A1 => n31648, A2 => n39714, B1 => n31712, B2 =>
                           n39708, C1 => n31584, C2 => n39702, ZN => n34197);
   U33623 : AOI221_X1 port map( B1 => n39474, B2 => n29388, C1 => n39468, C2 =>
                           n29452, A => n35471, ZN => n35466);
   U33624 : OAI222_X1 port map( A1 => n31648, A2 => n39462, B1 => n31712, B2 =>
                           n39456, C1 => n31584, C2 => n39450, ZN => n35471);
   U33625 : AOI221_X1 port map( B1 => n39726, B2 => n29387, C1 => n39720, C2 =>
                           n29451, A => n34216, ZN => n34211);
   U33626 : OAI222_X1 port map( A1 => n31647, A2 => n39714, B1 => n31711, B2 =>
                           n39708, C1 => n31583, C2 => n39702, ZN => n34216);
   U33627 : AOI221_X1 port map( B1 => n39474, B2 => n29387, C1 => n39468, C2 =>
                           n29451, A => n35490, ZN => n35485);
   U33628 : OAI222_X1 port map( A1 => n31647, A2 => n39462, B1 => n31711, B2 =>
                           n39456, C1 => n31583, C2 => n39450, ZN => n35490);
   U33629 : AOI221_X1 port map( B1 => n39725, B2 => n29386, C1 => n39719, C2 =>
                           n29450, A => n34235, ZN => n34230);
   U33630 : OAI222_X1 port map( A1 => n31646, A2 => n39713, B1 => n31710, B2 =>
                           n39707, C1 => n31582, C2 => n39701, ZN => n34235);
   U33631 : AOI221_X1 port map( B1 => n39473, B2 => n29386, C1 => n39467, C2 =>
                           n29450, A => n35509, ZN => n35504);
   U33632 : OAI222_X1 port map( A1 => n31646, A2 => n39461, B1 => n31710, B2 =>
                           n39455, C1 => n31582, C2 => n39449, ZN => n35509);
   U33633 : AOI221_X1 port map( B1 => n39725, B2 => n29385, C1 => n39719, C2 =>
                           n29449, A => n34254, ZN => n34249);
   U33634 : OAI222_X1 port map( A1 => n31645, A2 => n39713, B1 => n31709, B2 =>
                           n39707, C1 => n31581, C2 => n39701, ZN => n34254);
   U33635 : AOI221_X1 port map( B1 => n39473, B2 => n29385, C1 => n39467, C2 =>
                           n29449, A => n35528, ZN => n35523);
   U33636 : OAI222_X1 port map( A1 => n31645, A2 => n39461, B1 => n31709, B2 =>
                           n39455, C1 => n31581, C2 => n39449, ZN => n35528);
   U33637 : AOI221_X1 port map( B1 => n39725, B2 => n29384, C1 => n39719, C2 =>
                           n29448, A => n34273, ZN => n34268);
   U33638 : OAI222_X1 port map( A1 => n31644, A2 => n39713, B1 => n31708, B2 =>
                           n39707, C1 => n31580, C2 => n39701, ZN => n34273);
   U33639 : AOI221_X1 port map( B1 => n39473, B2 => n29384, C1 => n39467, C2 =>
                           n29448, A => n35547, ZN => n35542);
   U33640 : OAI222_X1 port map( A1 => n31644, A2 => n39461, B1 => n31708, B2 =>
                           n39455, C1 => n31580, C2 => n39449, ZN => n35547);
   U33641 : AOI221_X1 port map( B1 => n39725, B2 => n29383, C1 => n39719, C2 =>
                           n29447, A => n34292, ZN => n34287);
   U33642 : OAI222_X1 port map( A1 => n31643, A2 => n39713, B1 => n31707, B2 =>
                           n39707, C1 => n31579, C2 => n39701, ZN => n34292);
   U33643 : AOI221_X1 port map( B1 => n39473, B2 => n29383, C1 => n39467, C2 =>
                           n29447, A => n35566, ZN => n35561);
   U33644 : OAI222_X1 port map( A1 => n31643, A2 => n39461, B1 => n31707, B2 =>
                           n39455, C1 => n31579, C2 => n39449, ZN => n35566);
   U33645 : AOI221_X1 port map( B1 => n39725, B2 => n29382, C1 => n39719, C2 =>
                           n29446, A => n34311, ZN => n34306);
   U33646 : OAI222_X1 port map( A1 => n31642, A2 => n39713, B1 => n31706, B2 =>
                           n39707, C1 => n31578, C2 => n39701, ZN => n34311);
   U33647 : AOI221_X1 port map( B1 => n39473, B2 => n29382, C1 => n39467, C2 =>
                           n29446, A => n35585, ZN => n35580);
   U33648 : OAI222_X1 port map( A1 => n31642, A2 => n39461, B1 => n31706, B2 =>
                           n39455, C1 => n31578, C2 => n39449, ZN => n35585);
   U33649 : AOI221_X1 port map( B1 => n39725, B2 => n29381, C1 => n39719, C2 =>
                           n29445, A => n34330, ZN => n34325);
   U33650 : OAI222_X1 port map( A1 => n31641, A2 => n39713, B1 => n31705, B2 =>
                           n39707, C1 => n31577, C2 => n39701, ZN => n34330);
   U33651 : AOI221_X1 port map( B1 => n39473, B2 => n29381, C1 => n39467, C2 =>
                           n29445, A => n35604, ZN => n35599);
   U33652 : OAI222_X1 port map( A1 => n31641, A2 => n39461, B1 => n31705, B2 =>
                           n39455, C1 => n31577, C2 => n39449, ZN => n35604);
   U33653 : AOI221_X1 port map( B1 => n39725, B2 => n29380, C1 => n39719, C2 =>
                           n29444, A => n34349, ZN => n34344);
   U33654 : OAI222_X1 port map( A1 => n31640, A2 => n39713, B1 => n31704, B2 =>
                           n39707, C1 => n31576, C2 => n39701, ZN => n34349);
   U33655 : AOI221_X1 port map( B1 => n39473, B2 => n29380, C1 => n39467, C2 =>
                           n29444, A => n35623, ZN => n35618);
   U33656 : OAI222_X1 port map( A1 => n31640, A2 => n39461, B1 => n31704, B2 =>
                           n39455, C1 => n31576, C2 => n39449, ZN => n35623);
   U33657 : AOI221_X1 port map( B1 => n39725, B2 => n29379, C1 => n39719, C2 =>
                           n29443, A => n34368, ZN => n34363);
   U33658 : OAI222_X1 port map( A1 => n31639, A2 => n39713, B1 => n31703, B2 =>
                           n39707, C1 => n31575, C2 => n39701, ZN => n34368);
   U33659 : AOI221_X1 port map( B1 => n39473, B2 => n29379, C1 => n39467, C2 =>
                           n29443, A => n35642, ZN => n35637);
   U33660 : OAI222_X1 port map( A1 => n31639, A2 => n39461, B1 => n31703, B2 =>
                           n39455, C1 => n31575, C2 => n39449, ZN => n35642);
   U33661 : AOI221_X1 port map( B1 => n39725, B2 => n29378, C1 => n39719, C2 =>
                           n29442, A => n34387, ZN => n34382);
   U33662 : OAI222_X1 port map( A1 => n31638, A2 => n39713, B1 => n31702, B2 =>
                           n39707, C1 => n31574, C2 => n39701, ZN => n34387);
   U33663 : AOI221_X1 port map( B1 => n39473, B2 => n29378, C1 => n39467, C2 =>
                           n29442, A => n35661, ZN => n35656);
   U33664 : OAI222_X1 port map( A1 => n31638, A2 => n39461, B1 => n31702, B2 =>
                           n39455, C1 => n31574, C2 => n39449, ZN => n35661);
   U33665 : AOI221_X1 port map( B1 => n39725, B2 => n29377, C1 => n39719, C2 =>
                           n29441, A => n34406, ZN => n34401);
   U33666 : OAI222_X1 port map( A1 => n31637, A2 => n39713, B1 => n31701, B2 =>
                           n39707, C1 => n31573, C2 => n39701, ZN => n34406);
   U33667 : AOI221_X1 port map( B1 => n39473, B2 => n29377, C1 => n39467, C2 =>
                           n29441, A => n35680, ZN => n35675);
   U33668 : OAI222_X1 port map( A1 => n31637, A2 => n39461, B1 => n31701, B2 =>
                           n39455, C1 => n31573, C2 => n39449, ZN => n35680);
   U33669 : AOI221_X1 port map( B1 => n39725, B2 => n29376, C1 => n39719, C2 =>
                           n29440, A => n34425, ZN => n34420);
   U33670 : OAI222_X1 port map( A1 => n31636, A2 => n39713, B1 => n31700, B2 =>
                           n39707, C1 => n31572, C2 => n39701, ZN => n34425);
   U33671 : AOI221_X1 port map( B1 => n39473, B2 => n29376, C1 => n39467, C2 =>
                           n29440, A => n35699, ZN => n35694);
   U33672 : OAI222_X1 port map( A1 => n31636, A2 => n39461, B1 => n31700, B2 =>
                           n39455, C1 => n31572, C2 => n39449, ZN => n35699);
   U33673 : AOI221_X1 port map( B1 => n39725, B2 => n29375, C1 => n39719, C2 =>
                           n29439, A => n34444, ZN => n34439);
   U33674 : OAI222_X1 port map( A1 => n31635, A2 => n39713, B1 => n31699, B2 =>
                           n39707, C1 => n31571, C2 => n39701, ZN => n34444);
   U33675 : AOI221_X1 port map( B1 => n39473, B2 => n29375, C1 => n39467, C2 =>
                           n29439, A => n35718, ZN => n35713);
   U33676 : OAI222_X1 port map( A1 => n31635, A2 => n39461, B1 => n31699, B2 =>
                           n39455, C1 => n31571, C2 => n39449, ZN => n35718);
   U33677 : AOI221_X1 port map( B1 => n39724, B2 => n29374, C1 => n39718, C2 =>
                           n29438, A => n34463, ZN => n34458);
   U33678 : OAI222_X1 port map( A1 => n31634, A2 => n39712, B1 => n31698, B2 =>
                           n39706, C1 => n31570, C2 => n39700, ZN => n34463);
   U33679 : AOI221_X1 port map( B1 => n39472, B2 => n29374, C1 => n39466, C2 =>
                           n29438, A => n35737, ZN => n35732);
   U33680 : OAI222_X1 port map( A1 => n31634, A2 => n39460, B1 => n31698, B2 =>
                           n39454, C1 => n31570, C2 => n39448, ZN => n35737);
   U33681 : AOI221_X1 port map( B1 => n39724, B2 => n29373, C1 => n39718, C2 =>
                           n29437, A => n34482, ZN => n34477);
   U33682 : OAI222_X1 port map( A1 => n31633, A2 => n39712, B1 => n31697, B2 =>
                           n39706, C1 => n31569, C2 => n39700, ZN => n34482);
   U33683 : AOI221_X1 port map( B1 => n39472, B2 => n29373, C1 => n39466, C2 =>
                           n29437, A => n35756, ZN => n35751);
   U33684 : OAI222_X1 port map( A1 => n31633, A2 => n39460, B1 => n31697, B2 =>
                           n39454, C1 => n31569, C2 => n39448, ZN => n35756);
   U33685 : AOI221_X1 port map( B1 => n39724, B2 => n29372, C1 => n39718, C2 =>
                           n29436, A => n34501, ZN => n34496);
   U33686 : OAI222_X1 port map( A1 => n31632, A2 => n39712, B1 => n31696, B2 =>
                           n39706, C1 => n31568, C2 => n39700, ZN => n34501);
   U33687 : AOI221_X1 port map( B1 => n39472, B2 => n29372, C1 => n39466, C2 =>
                           n29436, A => n35775, ZN => n35770);
   U33688 : OAI222_X1 port map( A1 => n31632, A2 => n39460, B1 => n31696, B2 =>
                           n39454, C1 => n31568, C2 => n39448, ZN => n35775);
   U33689 : AOI221_X1 port map( B1 => n39724, B2 => n29371, C1 => n39718, C2 =>
                           n29435, A => n34520, ZN => n34515);
   U33690 : OAI222_X1 port map( A1 => n31631, A2 => n39712, B1 => n31695, B2 =>
                           n39706, C1 => n31567, C2 => n39700, ZN => n34520);
   U33691 : AOI221_X1 port map( B1 => n39472, B2 => n29371, C1 => n39466, C2 =>
                           n29435, A => n35794, ZN => n35789);
   U33692 : OAI222_X1 port map( A1 => n31631, A2 => n39460, B1 => n31695, B2 =>
                           n39454, C1 => n31567, C2 => n39448, ZN => n35794);
   U33693 : AOI221_X1 port map( B1 => n39724, B2 => n29370, C1 => n39718, C2 =>
                           n29434, A => n34539, ZN => n34534);
   U33694 : OAI222_X1 port map( A1 => n31630, A2 => n39712, B1 => n31694, B2 =>
                           n39706, C1 => n31566, C2 => n39700, ZN => n34539);
   U33695 : AOI221_X1 port map( B1 => n39472, B2 => n29370, C1 => n39466, C2 =>
                           n29434, A => n35813, ZN => n35808);
   U33696 : OAI222_X1 port map( A1 => n31630, A2 => n39460, B1 => n31694, B2 =>
                           n39454, C1 => n31566, C2 => n39448, ZN => n35813);
   U33697 : AOI221_X1 port map( B1 => n39724, B2 => n29369, C1 => n39718, C2 =>
                           n29433, A => n34558, ZN => n34553);
   U33698 : OAI222_X1 port map( A1 => n31629, A2 => n39712, B1 => n31693, B2 =>
                           n39706, C1 => n31565, C2 => n39700, ZN => n34558);
   U33699 : AOI221_X1 port map( B1 => n39472, B2 => n29369, C1 => n39466, C2 =>
                           n29433, A => n35832, ZN => n35827);
   U33700 : OAI222_X1 port map( A1 => n31629, A2 => n39460, B1 => n31693, B2 =>
                           n39454, C1 => n31565, C2 => n39448, ZN => n35832);
   U33701 : AOI221_X1 port map( B1 => n39724, B2 => n29368, C1 => n39718, C2 =>
                           n29432, A => n34577, ZN => n34572);
   U33702 : OAI222_X1 port map( A1 => n31628, A2 => n39712, B1 => n31692, B2 =>
                           n39706, C1 => n31564, C2 => n39700, ZN => n34577);
   U33703 : AOI221_X1 port map( B1 => n39472, B2 => n29368, C1 => n39466, C2 =>
                           n29432, A => n35851, ZN => n35846);
   U33704 : OAI222_X1 port map( A1 => n31628, A2 => n39460, B1 => n31692, B2 =>
                           n39454, C1 => n31564, C2 => n39448, ZN => n35851);
   U33705 : AOI221_X1 port map( B1 => n39724, B2 => n29367, C1 => n39718, C2 =>
                           n29431, A => n34596, ZN => n34591);
   U33706 : OAI222_X1 port map( A1 => n31627, A2 => n39712, B1 => n31691, B2 =>
                           n39706, C1 => n31563, C2 => n39700, ZN => n34596);
   U33707 : AOI221_X1 port map( B1 => n39472, B2 => n29367, C1 => n39466, C2 =>
                           n29431, A => n35870, ZN => n35865);
   U33708 : OAI222_X1 port map( A1 => n31627, A2 => n39460, B1 => n31691, B2 =>
                           n39454, C1 => n31563, C2 => n39448, ZN => n35870);
   U33709 : AOI221_X1 port map( B1 => n39724, B2 => n29366, C1 => n39718, C2 =>
                           n29430, A => n34615, ZN => n34610);
   U33710 : OAI222_X1 port map( A1 => n31626, A2 => n39712, B1 => n31690, B2 =>
                           n39706, C1 => n31562, C2 => n39700, ZN => n34615);
   U33711 : AOI221_X1 port map( B1 => n39472, B2 => n29366, C1 => n39466, C2 =>
                           n29430, A => n35889, ZN => n35884);
   U33712 : OAI222_X1 port map( A1 => n31626, A2 => n39460, B1 => n31690, B2 =>
                           n39454, C1 => n31562, C2 => n39448, ZN => n35889);
   U33713 : AOI221_X1 port map( B1 => n39724, B2 => n29365, C1 => n39718, C2 =>
                           n29429, A => n34634, ZN => n34629);
   U33714 : OAI222_X1 port map( A1 => n31625, A2 => n39712, B1 => n31689, B2 =>
                           n39706, C1 => n31561, C2 => n39700, ZN => n34634);
   U33715 : AOI221_X1 port map( B1 => n39472, B2 => n29365, C1 => n39466, C2 =>
                           n29429, A => n35908, ZN => n35903);
   U33716 : OAI222_X1 port map( A1 => n31625, A2 => n39460, B1 => n31689, B2 =>
                           n39454, C1 => n31561, C2 => n39448, ZN => n35908);
   U33717 : AOI221_X1 port map( B1 => n39724, B2 => n29364, C1 => n39718, C2 =>
                           n29428, A => n34653, ZN => n34648);
   U33718 : OAI222_X1 port map( A1 => n31624, A2 => n39712, B1 => n31688, B2 =>
                           n39706, C1 => n31560, C2 => n39700, ZN => n34653);
   U33719 : AOI221_X1 port map( B1 => n39472, B2 => n29364, C1 => n39466, C2 =>
                           n29428, A => n35927, ZN => n35922);
   U33720 : OAI222_X1 port map( A1 => n31624, A2 => n39460, B1 => n31688, B2 =>
                           n39454, C1 => n31560, C2 => n39448, ZN => n35927);
   U33721 : AOI221_X1 port map( B1 => n39724, B2 => n29363, C1 => n39718, C2 =>
                           n29427, A => n34682, ZN => n34667);
   U33722 : OAI222_X1 port map( A1 => n31623, A2 => n39712, B1 => n31687, B2 =>
                           n39706, C1 => n31559, C2 => n39700, ZN => n34682);
   U33723 : AOI221_X1 port map( B1 => n39472, B2 => n29363, C1 => n39466, C2 =>
                           n29427, A => n35956, ZN => n35941);
   U33724 : OAI222_X1 port map( A1 => n31623, A2 => n39460, B1 => n31687, B2 =>
                           n39454, C1 => n31559, C2 => n39448, ZN => n35956);
   U33725 : AOI221_X1 port map( B1 => n39072, B2 => n30469, C1 => n39066, C2 =>
                           n27996, A => n37027, ZN => n37020);
   U33726 : OAI222_X1 port map( A1 => n30597, A2 => n39060, B1 => n30661, B2 =>
                           n39054, C1 => n30533, C2 => n39048, ZN => n37027);
   U33727 : AOI221_X1 port map( B1 => n39192, B2 => n29095, C1 => n39186, C2 =>
                           n29159, A => n37019, ZN => n37012);
   U33728 : OAI222_X1 port map( A1 => n31483, A2 => n39180, B1 => n31547, B2 =>
                           n39174, C1 => n31419, C2 => n39168, ZN => n37019);
   U33729 : AOI221_X1 port map( B1 => n39073, B2 => n30468, C1 => n39067, C2 =>
                           n27995, A => n37008, ZN => n37001);
   U33730 : OAI222_X1 port map( A1 => n30596, A2 => n39061, B1 => n30660, B2 =>
                           n39055, C1 => n30532, C2 => n39049, ZN => n37008);
   U33731 : AOI221_X1 port map( B1 => n39193, B2 => n29094, C1 => n39187, C2 =>
                           n29158, A => n37000, ZN => n36993);
   U33732 : OAI222_X1 port map( A1 => n31482, A2 => n39181, B1 => n31546, B2 =>
                           n39175, C1 => n31418, C2 => n39169, ZN => n37000);
   U33733 : AOI221_X1 port map( B1 => n39073, B2 => n30467, C1 => n39067, C2 =>
                           n27994, A => n36989, ZN => n36982);
   U33734 : OAI222_X1 port map( A1 => n30595, A2 => n39061, B1 => n30659, B2 =>
                           n39055, C1 => n30531, C2 => n39049, ZN => n36989);
   U33735 : AOI221_X1 port map( B1 => n39193, B2 => n29093, C1 => n39187, C2 =>
                           n29157, A => n36981, ZN => n36974);
   U33736 : OAI222_X1 port map( A1 => n31481, A2 => n39181, B1 => n31545, B2 =>
                           n39175, C1 => n31417, C2 => n39169, ZN => n36981);
   U33737 : AOI221_X1 port map( B1 => n39073, B2 => n30466, C1 => n39067, C2 =>
                           n27993, A => n36970, ZN => n36963);
   U33738 : OAI222_X1 port map( A1 => n30594, A2 => n39061, B1 => n30658, B2 =>
                           n39055, C1 => n30530, C2 => n39049, ZN => n36970);
   U33739 : AOI221_X1 port map( B1 => n39193, B2 => n29092, C1 => n39187, C2 =>
                           n29156, A => n36962, ZN => n36955);
   U33740 : OAI222_X1 port map( A1 => n31480, A2 => n39181, B1 => n31544, B2 =>
                           n39175, C1 => n31416, C2 => n39169, ZN => n36962);
   U33741 : AOI221_X1 port map( B1 => n39073, B2 => n30465, C1 => n39067, C2 =>
                           n27992, A => n36951, ZN => n36944);
   U33742 : OAI222_X1 port map( A1 => n30593, A2 => n39061, B1 => n30657, B2 =>
                           n39055, C1 => n30529, C2 => n39049, ZN => n36951);
   U33743 : AOI221_X1 port map( B1 => n39193, B2 => n29091, C1 => n39187, C2 =>
                           n29155, A => n36943, ZN => n36936);
   U33744 : OAI222_X1 port map( A1 => n31479, A2 => n39181, B1 => n31543, B2 =>
                           n39175, C1 => n31415, C2 => n39169, ZN => n36943);
   U33745 : AOI221_X1 port map( B1 => n39073, B2 => n30464, C1 => n39067, C2 =>
                           n27991, A => n36932, ZN => n36925);
   U33746 : OAI222_X1 port map( A1 => n30592, A2 => n39061, B1 => n30656, B2 =>
                           n39055, C1 => n30528, C2 => n39049, ZN => n36932);
   U33747 : AOI221_X1 port map( B1 => n39193, B2 => n29090, C1 => n39187, C2 =>
                           n29154, A => n36924, ZN => n36917);
   U33748 : OAI222_X1 port map( A1 => n31478, A2 => n39181, B1 => n31542, B2 =>
                           n39175, C1 => n31414, C2 => n39169, ZN => n36924);
   U33749 : AOI221_X1 port map( B1 => n39073, B2 => n30463, C1 => n39067, C2 =>
                           n27990, A => n36913, ZN => n36906);
   U33750 : OAI222_X1 port map( A1 => n30591, A2 => n39061, B1 => n30655, B2 =>
                           n39055, C1 => n30527, C2 => n39049, ZN => n36913);
   U33751 : AOI221_X1 port map( B1 => n39193, B2 => n29089, C1 => n39187, C2 =>
                           n29153, A => n36905, ZN => n36898);
   U33752 : OAI222_X1 port map( A1 => n31477, A2 => n39181, B1 => n31541, B2 =>
                           n39175, C1 => n31413, C2 => n39169, ZN => n36905);
   U33753 : AOI221_X1 port map( B1 => n39073, B2 => n30462, C1 => n39067, C2 =>
                           n27989, A => n36894, ZN => n36887);
   U33754 : OAI222_X1 port map( A1 => n30590, A2 => n39061, B1 => n30654, B2 =>
                           n39055, C1 => n30526, C2 => n39049, ZN => n36894);
   U33755 : AOI221_X1 port map( B1 => n39193, B2 => n29088, C1 => n39187, C2 =>
                           n29152, A => n36886, ZN => n36879);
   U33756 : OAI222_X1 port map( A1 => n31476, A2 => n39181, B1 => n31540, B2 =>
                           n39175, C1 => n31412, C2 => n39169, ZN => n36886);
   U33757 : AOI221_X1 port map( B1 => n39073, B2 => n30461, C1 => n39067, C2 =>
                           n27988, A => n36875, ZN => n36868);
   U33758 : OAI222_X1 port map( A1 => n30589, A2 => n39061, B1 => n30653, B2 =>
                           n39055, C1 => n30525, C2 => n39049, ZN => n36875);
   U33759 : AOI221_X1 port map( B1 => n39193, B2 => n29087, C1 => n39187, C2 =>
                           n29151, A => n36867, ZN => n36860);
   U33760 : OAI222_X1 port map( A1 => n31475, A2 => n39181, B1 => n31539, B2 =>
                           n39175, C1 => n31411, C2 => n39169, ZN => n36867);
   U33761 : AOI221_X1 port map( B1 => n39073, B2 => n30460, C1 => n39067, C2 =>
                           n27987, A => n36856, ZN => n36849);
   U33762 : OAI222_X1 port map( A1 => n30588, A2 => n39061, B1 => n30652, B2 =>
                           n39055, C1 => n30524, C2 => n39049, ZN => n36856);
   U33763 : AOI221_X1 port map( B1 => n39193, B2 => n29086, C1 => n39187, C2 =>
                           n29150, A => n36848, ZN => n36841);
   U33764 : OAI222_X1 port map( A1 => n31474, A2 => n39181, B1 => n31538, B2 =>
                           n39175, C1 => n31410, C2 => n39169, ZN => n36848);
   U33765 : AOI221_X1 port map( B1 => n39073, B2 => n30459, C1 => n39067, C2 =>
                           n27986, A => n36837, ZN => n36830);
   U33766 : OAI222_X1 port map( A1 => n30587, A2 => n39061, B1 => n30651, B2 =>
                           n39055, C1 => n30523, C2 => n39049, ZN => n36837);
   U33767 : AOI221_X1 port map( B1 => n39193, B2 => n29085, C1 => n39187, C2 =>
                           n29149, A => n36829, ZN => n36822);
   U33768 : OAI222_X1 port map( A1 => n31473, A2 => n39181, B1 => n31537, B2 =>
                           n39175, C1 => n31409, C2 => n39169, ZN => n36829);
   U33769 : AOI221_X1 port map( B1 => n39073, B2 => n30458, C1 => n39067, C2 =>
                           n27985, A => n36818, ZN => n36811);
   U33770 : OAI222_X1 port map( A1 => n30586, A2 => n39061, B1 => n30650, B2 =>
                           n39055, C1 => n30522, C2 => n39049, ZN => n36818);
   U33771 : AOI221_X1 port map( B1 => n39193, B2 => n29084, C1 => n39187, C2 =>
                           n29148, A => n36810, ZN => n36803);
   U33772 : OAI222_X1 port map( A1 => n31472, A2 => n39181, B1 => n31536, B2 =>
                           n39175, C1 => n31408, C2 => n39169, ZN => n36810);
   U33773 : AOI221_X1 port map( B1 => n39073, B2 => n32546, C1 => n39067, C2 =>
                           n27984, A => n36799, ZN => n36792);
   U33774 : OAI222_X1 port map( A1 => n30585, A2 => n39061, B1 => n30649, B2 =>
                           n39055, C1 => n30521, C2 => n39049, ZN => n36799);
   U33775 : AOI221_X1 port map( B1 => n39193, B2 => n29083, C1 => n39187, C2 =>
                           n29147, A => n36791, ZN => n36784);
   U33776 : OAI222_X1 port map( A1 => n31471, A2 => n39181, B1 => n31535, B2 =>
                           n39175, C1 => n31407, C2 => n39169, ZN => n36791);
   U33777 : AOI221_X1 port map( B1 => n39074, B2 => n32545, C1 => n39068, C2 =>
                           n27983, A => n36780, ZN => n36773);
   U33778 : OAI222_X1 port map( A1 => n30584, A2 => n39062, B1 => n30648, B2 =>
                           n39056, C1 => n30520, C2 => n39050, ZN => n36780);
   U33779 : AOI221_X1 port map( B1 => n39194, B2 => n29082, C1 => n39188, C2 =>
                           n29146, A => n36772, ZN => n36765);
   U33780 : OAI222_X1 port map( A1 => n31470, A2 => n39182, B1 => n31534, B2 =>
                           n39176, C1 => n31406, C2 => n39170, ZN => n36772);
   U33781 : AOI221_X1 port map( B1 => n39074, B2 => n32544, C1 => n39068, C2 =>
                           n27982, A => n36761, ZN => n36754);
   U33782 : OAI222_X1 port map( A1 => n30583, A2 => n39062, B1 => n30647, B2 =>
                           n39056, C1 => n30519, C2 => n39050, ZN => n36761);
   U33783 : AOI221_X1 port map( B1 => n39194, B2 => n29081, C1 => n39188, C2 =>
                           n29145, A => n36753, ZN => n36746);
   U33784 : OAI222_X1 port map( A1 => n31469, A2 => n39182, B1 => n31533, B2 =>
                           n39176, C1 => n31405, C2 => n39170, ZN => n36753);
   U33785 : AOI221_X1 port map( B1 => n39074, B2 => n32543, C1 => n39068, C2 =>
                           n27981, A => n36742, ZN => n36735);
   U33786 : OAI222_X1 port map( A1 => n30582, A2 => n39062, B1 => n30646, B2 =>
                           n39056, C1 => n30518, C2 => n39050, ZN => n36742);
   U33787 : AOI221_X1 port map( B1 => n39194, B2 => n29080, C1 => n39188, C2 =>
                           n29144, A => n36734, ZN => n36727);
   U33788 : OAI222_X1 port map( A1 => n31468, A2 => n39182, B1 => n31532, B2 =>
                           n39176, C1 => n31404, C2 => n39170, ZN => n36734);
   U33789 : AOI221_X1 port map( B1 => n39074, B2 => n32542, C1 => n39068, C2 =>
                           n27980, A => n36723, ZN => n36716);
   U33790 : OAI222_X1 port map( A1 => n30581, A2 => n39062, B1 => n30645, B2 =>
                           n39056, C1 => n30517, C2 => n39050, ZN => n36723);
   U33791 : AOI221_X1 port map( B1 => n39194, B2 => n29079, C1 => n39188, C2 =>
                           n29143, A => n36715, ZN => n36708);
   U33792 : OAI222_X1 port map( A1 => n31467, A2 => n39182, B1 => n31531, B2 =>
                           n39176, C1 => n31403, C2 => n39170, ZN => n36715);
   U33793 : AOI221_X1 port map( B1 => n39074, B2 => n32541, C1 => n39068, C2 =>
                           n27979, A => n36704, ZN => n36697);
   U33794 : OAI222_X1 port map( A1 => n30580, A2 => n39062, B1 => n30644, B2 =>
                           n39056, C1 => n30516, C2 => n39050, ZN => n36704);
   U33795 : AOI221_X1 port map( B1 => n39194, B2 => n29078, C1 => n39188, C2 =>
                           n29142, A => n36696, ZN => n36689);
   U33796 : OAI222_X1 port map( A1 => n31466, A2 => n39182, B1 => n31530, B2 =>
                           n39176, C1 => n31402, C2 => n39170, ZN => n36696);
   U33797 : AOI221_X1 port map( B1 => n39074, B2 => n32540, C1 => n39068, C2 =>
                           n27978, A => n36685, ZN => n36678);
   U33798 : OAI222_X1 port map( A1 => n30579, A2 => n39062, B1 => n30643, B2 =>
                           n39056, C1 => n30515, C2 => n39050, ZN => n36685);
   U33799 : AOI221_X1 port map( B1 => n39194, B2 => n29077, C1 => n39188, C2 =>
                           n29141, A => n36677, ZN => n36670);
   U33800 : OAI222_X1 port map( A1 => n31465, A2 => n39182, B1 => n31529, B2 =>
                           n39176, C1 => n31401, C2 => n39170, ZN => n36677);
   U33801 : AOI221_X1 port map( B1 => n39074, B2 => n32539, C1 => n39068, C2 =>
                           n27977, A => n36666, ZN => n36659);
   U33802 : OAI222_X1 port map( A1 => n30578, A2 => n39062, B1 => n30642, B2 =>
                           n39056, C1 => n30514, C2 => n39050, ZN => n36666);
   U33803 : AOI221_X1 port map( B1 => n39194, B2 => n29076, C1 => n39188, C2 =>
                           n29140, A => n36658, ZN => n36651);
   U33804 : OAI222_X1 port map( A1 => n31464, A2 => n39182, B1 => n31528, B2 =>
                           n39176, C1 => n31400, C2 => n39170, ZN => n36658);
   U33805 : AOI221_X1 port map( B1 => n39074, B2 => n32538, C1 => n39068, C2 =>
                           n27976, A => n36647, ZN => n36640);
   U33806 : OAI222_X1 port map( A1 => n30577, A2 => n39062, B1 => n30641, B2 =>
                           n39056, C1 => n30513, C2 => n39050, ZN => n36647);
   U33807 : AOI221_X1 port map( B1 => n39194, B2 => n29075, C1 => n39188, C2 =>
                           n29139, A => n36639, ZN => n36632);
   U33808 : OAI222_X1 port map( A1 => n31463, A2 => n39182, B1 => n31527, B2 =>
                           n39176, C1 => n31399, C2 => n39170, ZN => n36639);
   U33809 : AOI221_X1 port map( B1 => n39074, B2 => n32537, C1 => n39068, C2 =>
                           n27975, A => n36628, ZN => n36621);
   U33810 : OAI222_X1 port map( A1 => n30576, A2 => n39062, B1 => n30640, B2 =>
                           n39056, C1 => n30512, C2 => n39050, ZN => n36628);
   U33811 : AOI221_X1 port map( B1 => n39194, B2 => n29074, C1 => n39188, C2 =>
                           n29138, A => n36620, ZN => n36613);
   U33812 : OAI222_X1 port map( A1 => n31462, A2 => n39182, B1 => n31526, B2 =>
                           n39176, C1 => n31398, C2 => n39170, ZN => n36620);
   U33813 : AOI221_X1 port map( B1 => n39074, B2 => n32536, C1 => n39068, C2 =>
                           n27974, A => n36609, ZN => n36602);
   U33814 : OAI222_X1 port map( A1 => n30575, A2 => n39062, B1 => n30639, B2 =>
                           n39056, C1 => n30511, C2 => n39050, ZN => n36609);
   U33815 : AOI221_X1 port map( B1 => n39194, B2 => n29073, C1 => n39188, C2 =>
                           n29137, A => n36601, ZN => n36594);
   U33816 : OAI222_X1 port map( A1 => n31461, A2 => n39182, B1 => n31525, B2 =>
                           n39176, C1 => n31397, C2 => n39170, ZN => n36601);
   U33817 : AOI221_X1 port map( B1 => n39074, B2 => n32535, C1 => n39068, C2 =>
                           n27973, A => n36590, ZN => n36583);
   U33818 : OAI222_X1 port map( A1 => n30574, A2 => n39062, B1 => n30638, B2 =>
                           n39056, C1 => n30510, C2 => n39050, ZN => n36590);
   U33819 : AOI221_X1 port map( B1 => n39194, B2 => n29072, C1 => n39188, C2 =>
                           n29136, A => n36582, ZN => n36575);
   U33820 : OAI222_X1 port map( A1 => n31460, A2 => n39182, B1 => n31524, B2 =>
                           n39176, C1 => n31396, C2 => n39170, ZN => n36582);
   U33821 : AOI221_X1 port map( B1 => n39074, B2 => n32534, C1 => n39068, C2 =>
                           n27972, A => n36571, ZN => n36564);
   U33822 : OAI222_X1 port map( A1 => n30573, A2 => n39062, B1 => n30637, B2 =>
                           n39056, C1 => n30509, C2 => n39050, ZN => n36571);
   U33823 : AOI221_X1 port map( B1 => n39194, B2 => n29071, C1 => n39188, C2 =>
                           n29135, A => n36563, ZN => n36556);
   U33824 : OAI222_X1 port map( A1 => n31459, A2 => n39182, B1 => n31523, B2 =>
                           n39176, C1 => n31395, C2 => n39170, ZN => n36563);
   U33825 : AOI221_X1 port map( B1 => n39075, B2 => n32533, C1 => n39069, C2 =>
                           n27971, A => n36552, ZN => n36545);
   U33826 : OAI222_X1 port map( A1 => n30572, A2 => n39063, B1 => n30636, B2 =>
                           n39057, C1 => n30508, C2 => n39051, ZN => n36552);
   U33827 : AOI221_X1 port map( B1 => n39195, B2 => n29070, C1 => n39189, C2 =>
                           n29134, A => n36544, ZN => n36537);
   U33828 : OAI222_X1 port map( A1 => n31458, A2 => n39183, B1 => n31522, B2 =>
                           n39177, C1 => n31394, C2 => n39171, ZN => n36544);
   U33829 : AOI221_X1 port map( B1 => n39075, B2 => n32532, C1 => n39069, C2 =>
                           n27970, A => n36533, ZN => n36526);
   U33830 : OAI222_X1 port map( A1 => n30571, A2 => n39063, B1 => n30635, B2 =>
                           n39057, C1 => n30507, C2 => n39051, ZN => n36533);
   U33831 : AOI221_X1 port map( B1 => n39195, B2 => n29069, C1 => n39189, C2 =>
                           n29133, A => n36525, ZN => n36518);
   U33832 : OAI222_X1 port map( A1 => n31457, A2 => n39183, B1 => n31521, B2 =>
                           n39177, C1 => n31393, C2 => n39171, ZN => n36525);
   U33833 : AOI221_X1 port map( B1 => n39075, B2 => n32531, C1 => n39069, C2 =>
                           n27969, A => n36514, ZN => n36507);
   U33834 : OAI222_X1 port map( A1 => n30570, A2 => n39063, B1 => n30634, B2 =>
                           n39057, C1 => n30506, C2 => n39051, ZN => n36514);
   U33835 : AOI221_X1 port map( B1 => n39195, B2 => n29068, C1 => n39189, C2 =>
                           n29132, A => n36506, ZN => n36499);
   U33836 : OAI222_X1 port map( A1 => n31456, A2 => n39183, B1 => n31520, B2 =>
                           n39177, C1 => n31392, C2 => n39171, ZN => n36506);
   U33837 : AOI221_X1 port map( B1 => n39075, B2 => n32530, C1 => n39069, C2 =>
                           n27968, A => n36495, ZN => n36488);
   U33838 : OAI222_X1 port map( A1 => n30569, A2 => n39063, B1 => n30633, B2 =>
                           n39057, C1 => n30505, C2 => n39051, ZN => n36495);
   U33839 : AOI221_X1 port map( B1 => n39195, B2 => n29067, C1 => n39189, C2 =>
                           n29131, A => n36487, ZN => n36480);
   U33840 : OAI222_X1 port map( A1 => n31455, A2 => n39183, B1 => n31519, B2 =>
                           n39177, C1 => n31391, C2 => n39171, ZN => n36487);
   U33841 : AOI221_X1 port map( B1 => n39075, B2 => n32529, C1 => n39069, C2 =>
                           n27967, A => n36476, ZN => n36469);
   U33842 : OAI222_X1 port map( A1 => n30568, A2 => n39063, B1 => n30632, B2 =>
                           n39057, C1 => n30504, C2 => n39051, ZN => n36476);
   U33843 : AOI221_X1 port map( B1 => n39195, B2 => n29066, C1 => n39189, C2 =>
                           n29130, A => n36468, ZN => n36461);
   U33844 : OAI222_X1 port map( A1 => n31454, A2 => n39183, B1 => n31518, B2 =>
                           n39177, C1 => n31390, C2 => n39171, ZN => n36468);
   U33845 : AOI221_X1 port map( B1 => n39075, B2 => n32528, C1 => n39069, C2 =>
                           n27966, A => n36457, ZN => n36450);
   U33846 : OAI222_X1 port map( A1 => n30567, A2 => n39063, B1 => n30631, B2 =>
                           n39057, C1 => n30503, C2 => n39051, ZN => n36457);
   U33847 : AOI221_X1 port map( B1 => n39195, B2 => n29065, C1 => n39189, C2 =>
                           n29129, A => n36449, ZN => n36442);
   U33848 : OAI222_X1 port map( A1 => n31453, A2 => n39183, B1 => n31517, B2 =>
                           n39177, C1 => n31389, C2 => n39171, ZN => n36449);
   U33849 : AOI221_X1 port map( B1 => n39075, B2 => n32527, C1 => n39069, C2 =>
                           n27965, A => n36438, ZN => n36431);
   U33850 : OAI222_X1 port map( A1 => n30566, A2 => n39063, B1 => n30630, B2 =>
                           n39057, C1 => n30502, C2 => n39051, ZN => n36438);
   U33851 : AOI221_X1 port map( B1 => n39195, B2 => n29064, C1 => n39189, C2 =>
                           n29128, A => n36430, ZN => n36423);
   U33852 : OAI222_X1 port map( A1 => n31452, A2 => n39183, B1 => n31516, B2 =>
                           n39177, C1 => n31388, C2 => n39171, ZN => n36430);
   U33853 : AOI221_X1 port map( B1 => n39075, B2 => n32526, C1 => n39069, C2 =>
                           n27964, A => n36419, ZN => n36412);
   U33854 : OAI222_X1 port map( A1 => n30565, A2 => n39063, B1 => n30629, B2 =>
                           n39057, C1 => n30501, C2 => n39051, ZN => n36419);
   U33855 : AOI221_X1 port map( B1 => n39195, B2 => n29063, C1 => n39189, C2 =>
                           n29127, A => n36411, ZN => n36404);
   U33856 : OAI222_X1 port map( A1 => n31451, A2 => n39183, B1 => n31515, B2 =>
                           n39177, C1 => n31387, C2 => n39171, ZN => n36411);
   U33857 : AOI221_X1 port map( B1 => n39075, B2 => n32525, C1 => n39069, C2 =>
                           n27963, A => n36400, ZN => n36393);
   U33858 : OAI222_X1 port map( A1 => n30564, A2 => n39063, B1 => n30628, B2 =>
                           n39057, C1 => n30500, C2 => n39051, ZN => n36400);
   U33859 : AOI221_X1 port map( B1 => n39195, B2 => n29062, C1 => n39189, C2 =>
                           n29126, A => n36392, ZN => n36385);
   U33860 : OAI222_X1 port map( A1 => n31450, A2 => n39183, B1 => n31514, B2 =>
                           n39177, C1 => n31386, C2 => n39171, ZN => n36392);
   U33861 : AOI221_X1 port map( B1 => n39075, B2 => n32524, C1 => n39069, C2 =>
                           n27962, A => n36381, ZN => n36374);
   U33862 : OAI222_X1 port map( A1 => n30563, A2 => n39063, B1 => n30627, B2 =>
                           n39057, C1 => n30499, C2 => n39051, ZN => n36381);
   U33863 : AOI221_X1 port map( B1 => n39195, B2 => n29061, C1 => n39189, C2 =>
                           n29125, A => n36373, ZN => n36366);
   U33864 : OAI222_X1 port map( A1 => n31449, A2 => n39183, B1 => n31513, B2 =>
                           n39177, C1 => n31385, C2 => n39171, ZN => n36373);
   U33865 : AOI221_X1 port map( B1 => n39075, B2 => n32523, C1 => n39069, C2 =>
                           n27961, A => n36362, ZN => n36355);
   U33866 : OAI222_X1 port map( A1 => n30562, A2 => n39063, B1 => n30626, B2 =>
                           n39057, C1 => n30498, C2 => n39051, ZN => n36362);
   U33867 : AOI221_X1 port map( B1 => n39195, B2 => n29060, C1 => n39189, C2 =>
                           n29124, A => n36354, ZN => n36347);
   U33868 : OAI222_X1 port map( A1 => n31448, A2 => n39183, B1 => n31512, B2 =>
                           n39177, C1 => n31384, C2 => n39171, ZN => n36354);
   U33869 : AOI221_X1 port map( B1 => n39075, B2 => n32522, C1 => n39069, C2 =>
                           n27960, A => n36343, ZN => n36336);
   U33870 : OAI222_X1 port map( A1 => n30561, A2 => n39063, B1 => n30625, B2 =>
                           n39057, C1 => n30497, C2 => n39051, ZN => n36343);
   U33871 : AOI221_X1 port map( B1 => n39195, B2 => n29059, C1 => n39189, C2 =>
                           n29123, A => n36335, ZN => n36328);
   U33872 : OAI222_X1 port map( A1 => n31447, A2 => n39183, B1 => n31511, B2 =>
                           n39177, C1 => n31383, C2 => n39171, ZN => n36335);
   U33873 : AOI221_X1 port map( B1 => n39076, B2 => n32521, C1 => n39070, C2 =>
                           n27959, A => n36324, ZN => n36317);
   U33874 : OAI222_X1 port map( A1 => n30560, A2 => n39064, B1 => n30624, B2 =>
                           n39058, C1 => n30496, C2 => n39052, ZN => n36324);
   U33875 : AOI221_X1 port map( B1 => n39196, B2 => n29058, C1 => n39190, C2 =>
                           n29122, A => n36316, ZN => n36309);
   U33876 : OAI222_X1 port map( A1 => n31446, A2 => n39184, B1 => n31510, B2 =>
                           n39178, C1 => n31382, C2 => n39172, ZN => n36316);
   U33877 : AOI221_X1 port map( B1 => n39076, B2 => n32520, C1 => n39070, C2 =>
                           n27958, A => n36305, ZN => n36298);
   U33878 : OAI222_X1 port map( A1 => n30559, A2 => n39064, B1 => n30623, B2 =>
                           n39058, C1 => n30495, C2 => n39052, ZN => n36305);
   U33879 : AOI221_X1 port map( B1 => n39196, B2 => n29057, C1 => n39190, C2 =>
                           n29121, A => n36297, ZN => n36290);
   U33880 : OAI222_X1 port map( A1 => n31445, A2 => n39184, B1 => n31509, B2 =>
                           n39178, C1 => n31381, C2 => n39172, ZN => n36297);
   U33881 : AOI221_X1 port map( B1 => n39076, B2 => n32519, C1 => n39070, C2 =>
                           n27957, A => n36286, ZN => n36279);
   U33882 : OAI222_X1 port map( A1 => n30558, A2 => n39064, B1 => n30622, B2 =>
                           n39058, C1 => n30494, C2 => n39052, ZN => n36286);
   U33883 : AOI221_X1 port map( B1 => n39196, B2 => n29056, C1 => n39190, C2 =>
                           n29120, A => n36278, ZN => n36271);
   U33884 : OAI222_X1 port map( A1 => n31444, A2 => n39184, B1 => n31508, B2 =>
                           n39178, C1 => n31380, C2 => n39172, ZN => n36278);
   U33885 : AOI221_X1 port map( B1 => n39076, B2 => n32518, C1 => n39070, C2 =>
                           n27956, A => n36267, ZN => n36260);
   U33886 : OAI222_X1 port map( A1 => n30557, A2 => n39064, B1 => n30621, B2 =>
                           n39058, C1 => n30493, C2 => n39052, ZN => n36267);
   U33887 : AOI221_X1 port map( B1 => n39196, B2 => n29055, C1 => n39190, C2 =>
                           n29119, A => n36259, ZN => n36252);
   U33888 : OAI222_X1 port map( A1 => n31443, A2 => n39184, B1 => n31507, B2 =>
                           n39178, C1 => n31379, C2 => n39172, ZN => n36259);
   U33889 : AOI221_X1 port map( B1 => n39076, B2 => n32517, C1 => n39070, C2 =>
                           n27955, A => n36248, ZN => n36241);
   U33890 : OAI222_X1 port map( A1 => n30556, A2 => n39064, B1 => n30620, B2 =>
                           n39058, C1 => n30492, C2 => n39052, ZN => n36248);
   U33891 : AOI221_X1 port map( B1 => n39196, B2 => n29054, C1 => n39190, C2 =>
                           n29118, A => n36240, ZN => n36233);
   U33892 : OAI222_X1 port map( A1 => n31442, A2 => n39184, B1 => n31506, B2 =>
                           n39178, C1 => n31378, C2 => n39172, ZN => n36240);
   U33893 : AOI221_X1 port map( B1 => n39076, B2 => n32516, C1 => n39070, C2 =>
                           n27954, A => n36229, ZN => n36222);
   U33894 : OAI222_X1 port map( A1 => n30555, A2 => n39064, B1 => n30619, B2 =>
                           n39058, C1 => n30491, C2 => n39052, ZN => n36229);
   U33895 : AOI221_X1 port map( B1 => n39196, B2 => n29053, C1 => n39190, C2 =>
                           n29117, A => n36221, ZN => n36214);
   U33896 : OAI222_X1 port map( A1 => n31441, A2 => n39184, B1 => n31505, B2 =>
                           n39178, C1 => n31377, C2 => n39172, ZN => n36221);
   U33897 : AOI221_X1 port map( B1 => n39072, B2 => n30479, C1 => n39066, C2 =>
                           n28006, A => n37217, ZN => n37210);
   U33898 : OAI222_X1 port map( A1 => n30607, A2 => n39060, B1 => n30671, B2 =>
                           n39054, C1 => n30543, C2 => n39048, ZN => n37217);
   U33899 : AOI221_X1 port map( B1 => n39192, B2 => n29105, C1 => n39186, C2 =>
                           n29169, A => n37209, ZN => n37202);
   U33900 : OAI222_X1 port map( A1 => n31493, A2 => n39180, B1 => n31557, B2 =>
                           n39174, C1 => n31429, C2 => n39168, ZN => n37209);
   U33901 : AOI221_X1 port map( B1 => n39072, B2 => n30478, C1 => n39066, C2 =>
                           n28005, A => n37198, ZN => n37191);
   U33902 : OAI222_X1 port map( A1 => n30606, A2 => n39060, B1 => n30670, B2 =>
                           n39054, C1 => n30542, C2 => n39048, ZN => n37198);
   U33903 : AOI221_X1 port map( B1 => n39192, B2 => n29104, C1 => n39186, C2 =>
                           n29168, A => n37190, ZN => n37183);
   U33904 : OAI222_X1 port map( A1 => n31492, A2 => n39180, B1 => n31556, B2 =>
                           n39174, C1 => n31428, C2 => n39168, ZN => n37190);
   U33905 : AOI221_X1 port map( B1 => n39072, B2 => n30477, C1 => n39066, C2 =>
                           n28004, A => n37179, ZN => n37172);
   U33906 : OAI222_X1 port map( A1 => n30605, A2 => n39060, B1 => n30669, B2 =>
                           n39054, C1 => n30541, C2 => n39048, ZN => n37179);
   U33907 : AOI221_X1 port map( B1 => n39192, B2 => n29103, C1 => n39186, C2 =>
                           n29167, A => n37171, ZN => n37164);
   U33908 : OAI222_X1 port map( A1 => n31491, A2 => n39180, B1 => n31555, B2 =>
                           n39174, C1 => n31427, C2 => n39168, ZN => n37171);
   U33909 : AOI221_X1 port map( B1 => n39072, B2 => n30476, C1 => n39066, C2 =>
                           n28003, A => n37160, ZN => n37153);
   U33910 : OAI222_X1 port map( A1 => n30604, A2 => n39060, B1 => n30668, B2 =>
                           n39054, C1 => n30540, C2 => n39048, ZN => n37160);
   U33911 : AOI221_X1 port map( B1 => n39192, B2 => n29102, C1 => n39186, C2 =>
                           n29166, A => n37152, ZN => n37145);
   U33912 : OAI222_X1 port map( A1 => n31490, A2 => n39180, B1 => n31554, B2 =>
                           n39174, C1 => n31426, C2 => n39168, ZN => n37152);
   U33913 : AOI221_X1 port map( B1 => n39072, B2 => n30475, C1 => n39066, C2 =>
                           n28002, A => n37141, ZN => n37134);
   U33914 : OAI222_X1 port map( A1 => n30603, A2 => n39060, B1 => n30667, B2 =>
                           n39054, C1 => n30539, C2 => n39048, ZN => n37141);
   U33915 : AOI221_X1 port map( B1 => n39192, B2 => n29101, C1 => n39186, C2 =>
                           n29165, A => n37133, ZN => n37126);
   U33916 : OAI222_X1 port map( A1 => n31489, A2 => n39180, B1 => n31553, B2 =>
                           n39174, C1 => n31425, C2 => n39168, ZN => n37133);
   U33917 : AOI221_X1 port map( B1 => n39077, B2 => n32507, C1 => n39071, C2 =>
                           n27947, A => n36096, ZN => n36089);
   U33918 : OAI222_X1 port map( A1 => n30548, A2 => n39065, B1 => n30612, B2 =>
                           n39059, C1 => n30484, C2 => n39053, ZN => n36096);
   U33919 : AOI221_X1 port map( B1 => n39197, B2 => n29046, C1 => n39191, C2 =>
                           n29110, A => n36088, ZN => n36081);
   U33920 : OAI222_X1 port map( A1 => n31434, A2 => n39185, B1 => n31498, B2 =>
                           n39179, C1 => n31370, C2 => n39173, ZN => n36088);
   U33921 : AOI221_X1 port map( B1 => n39077, B2 => n32506, C1 => n39071, C2 =>
                           n27946, A => n36077, ZN => n36070);
   U33922 : OAI222_X1 port map( A1 => n30547, A2 => n39065, B1 => n30611, B2 =>
                           n39059, C1 => n30483, C2 => n39053, ZN => n36077);
   U33923 : AOI221_X1 port map( B1 => n39197, B2 => n29045, C1 => n39191, C2 =>
                           n29109, A => n36069, ZN => n36062);
   U33924 : OAI222_X1 port map( A1 => n31433, A2 => n39185, B1 => n31497, B2 =>
                           n39179, C1 => n31369, C2 => n39173, ZN => n36069);
   U33925 : AOI221_X1 port map( B1 => n39077, B2 => n32509, C1 => n39071, C2 =>
                           n27945, A => n36058, ZN => n36051);
   U33926 : OAI222_X1 port map( A1 => n30546, A2 => n39065, B1 => n30610, B2 =>
                           n39059, C1 => n30482, C2 => n39053, ZN => n36058);
   U33927 : AOI221_X1 port map( B1 => n39197, B2 => n29044, C1 => n39191, C2 =>
                           n29108, A => n36050, ZN => n36043);
   U33928 : OAI222_X1 port map( A1 => n31432, A2 => n39185, B1 => n31496, B2 =>
                           n39179, C1 => n31368, C2 => n39173, ZN => n36050);
   U33929 : AOI221_X1 port map( B1 => n39077, B2 => n32508, C1 => n39071, C2 =>
                           n27944, A => n36036, ZN => n36012);
   U33930 : OAI222_X1 port map( A1 => n30545, A2 => n39065, B1 => n30609, B2 =>
                           n39059, C1 => n30481, C2 => n39053, ZN => n36036);
   U33931 : AOI221_X1 port map( B1 => n39197, B2 => n29043, C1 => n39191, C2 =>
                           n29107, A => n36008, ZN => n35984);
   U33932 : OAI222_X1 port map( A1 => n31431, A2 => n39185, B1 => n31495, B2 =>
                           n39179, C1 => n31367, C2 => n39173, ZN => n36008);
   U33933 : AOI221_X1 port map( B1 => n39072, B2 => n30480, C1 => n39066, C2 =>
                           n28007, A => n37250, ZN => n37241);
   U33934 : OAI222_X1 port map( A1 => n30608, A2 => n39060, B1 => n30672, B2 =>
                           n39054, C1 => n30544, C2 => n39048, ZN => n37250);
   U33935 : AOI221_X1 port map( B1 => n39192, B2 => n29106, C1 => n39186, C2 =>
                           n29170, A => n37238, ZN => n37221);
   U33936 : OAI222_X1 port map( A1 => n31494, A2 => n39180, B1 => n31558, B2 =>
                           n39174, C1 => n31430, C2 => n39168, ZN => n37238);
   U33937 : AOI221_X1 port map( B1 => n39072, B2 => n30474, C1 => n39066, C2 =>
                           n28001, A => n37122, ZN => n37115);
   U33938 : OAI222_X1 port map( A1 => n30602, A2 => n39060, B1 => n30666, B2 =>
                           n39054, C1 => n30538, C2 => n39048, ZN => n37122);
   U33939 : AOI221_X1 port map( B1 => n39192, B2 => n29100, C1 => n39186, C2 =>
                           n29164, A => n37114, ZN => n37107);
   U33940 : OAI222_X1 port map( A1 => n31488, A2 => n39180, B1 => n31552, B2 =>
                           n39174, C1 => n31424, C2 => n39168, ZN => n37114);
   U33941 : AOI221_X1 port map( B1 => n39072, B2 => n30473, C1 => n39066, C2 =>
                           n28000, A => n37103, ZN => n37096);
   U33942 : OAI222_X1 port map( A1 => n30601, A2 => n39060, B1 => n30665, B2 =>
                           n39054, C1 => n30537, C2 => n39048, ZN => n37103);
   U33943 : AOI221_X1 port map( B1 => n39192, B2 => n29099, C1 => n39186, C2 =>
                           n29163, A => n37095, ZN => n37088);
   U33944 : OAI222_X1 port map( A1 => n31487, A2 => n39180, B1 => n31551, B2 =>
                           n39174, C1 => n31423, C2 => n39168, ZN => n37095);
   U33945 : AOI221_X1 port map( B1 => n39072, B2 => n30472, C1 => n39066, C2 =>
                           n27999, A => n37084, ZN => n37077);
   U33946 : OAI222_X1 port map( A1 => n30600, A2 => n39060, B1 => n30664, B2 =>
                           n39054, C1 => n30536, C2 => n39048, ZN => n37084);
   U33947 : AOI221_X1 port map( B1 => n39192, B2 => n29098, C1 => n39186, C2 =>
                           n29162, A => n37076, ZN => n37069);
   U33948 : OAI222_X1 port map( A1 => n31486, A2 => n39180, B1 => n31550, B2 =>
                           n39174, C1 => n31422, C2 => n39168, ZN => n37076);
   U33949 : AOI221_X1 port map( B1 => n39072, B2 => n30471, C1 => n39066, C2 =>
                           n27998, A => n37065, ZN => n37058);
   U33950 : OAI222_X1 port map( A1 => n30599, A2 => n39060, B1 => n30663, B2 =>
                           n39054, C1 => n30535, C2 => n39048, ZN => n37065);
   U33951 : AOI221_X1 port map( B1 => n39192, B2 => n29097, C1 => n39186, C2 =>
                           n29161, A => n37057, ZN => n37050);
   U33952 : OAI222_X1 port map( A1 => n31485, A2 => n39180, B1 => n31549, B2 =>
                           n39174, C1 => n31421, C2 => n39168, ZN => n37057);
   U33953 : AOI221_X1 port map( B1 => n39072, B2 => n30470, C1 => n39066, C2 =>
                           n27997, A => n37046, ZN => n37039);
   U33954 : OAI222_X1 port map( A1 => n30598, A2 => n39060, B1 => n30662, B2 =>
                           n39054, C1 => n30534, C2 => n39048, ZN => n37046);
   U33955 : AOI221_X1 port map( B1 => n39192, B2 => n29096, C1 => n39186, C2 =>
                           n29160, A => n37038, ZN => n37031);
   U33956 : OAI222_X1 port map( A1 => n31484, A2 => n39180, B1 => n31548, B2 =>
                           n39174, C1 => n31420, C2 => n39168, ZN => n37038);
   U33957 : AOI221_X1 port map( B1 => n39076, B2 => n32515, C1 => n39070, C2 =>
                           n27953, A => n36210, ZN => n36203);
   U33958 : OAI222_X1 port map( A1 => n30554, A2 => n39064, B1 => n30618, B2 =>
                           n39058, C1 => n30490, C2 => n39052, ZN => n36210);
   U33959 : AOI221_X1 port map( B1 => n39196, B2 => n29052, C1 => n39190, C2 =>
                           n29116, A => n36202, ZN => n36195);
   U33960 : OAI222_X1 port map( A1 => n31440, A2 => n39184, B1 => n31504, B2 =>
                           n39178, C1 => n31376, C2 => n39172, ZN => n36202);
   U33961 : AOI221_X1 port map( B1 => n39076, B2 => n32514, C1 => n39070, C2 =>
                           n27952, A => n36191, ZN => n36184);
   U33962 : OAI222_X1 port map( A1 => n30553, A2 => n39064, B1 => n30617, B2 =>
                           n39058, C1 => n30489, C2 => n39052, ZN => n36191);
   U33963 : AOI221_X1 port map( B1 => n39196, B2 => n29051, C1 => n39190, C2 =>
                           n29115, A => n36183, ZN => n36176);
   U33964 : OAI222_X1 port map( A1 => n31439, A2 => n39184, B1 => n31503, B2 =>
                           n39178, C1 => n31375, C2 => n39172, ZN => n36183);
   U33965 : AOI221_X1 port map( B1 => n39076, B2 => n32513, C1 => n39070, C2 =>
                           n27951, A => n36172, ZN => n36165);
   U33966 : OAI222_X1 port map( A1 => n30552, A2 => n39064, B1 => n30616, B2 =>
                           n39058, C1 => n30488, C2 => n39052, ZN => n36172);
   U33967 : AOI221_X1 port map( B1 => n39196, B2 => n29050, C1 => n39190, C2 =>
                           n29114, A => n36164, ZN => n36157);
   U33968 : OAI222_X1 port map( A1 => n31438, A2 => n39184, B1 => n31502, B2 =>
                           n39178, C1 => n31374, C2 => n39172, ZN => n36164);
   U33969 : AOI221_X1 port map( B1 => n39076, B2 => n32512, C1 => n39070, C2 =>
                           n27950, A => n36153, ZN => n36146);
   U33970 : OAI222_X1 port map( A1 => n30551, A2 => n39064, B1 => n30615, B2 =>
                           n39058, C1 => n30487, C2 => n39052, ZN => n36153);
   U33971 : AOI221_X1 port map( B1 => n39196, B2 => n29049, C1 => n39190, C2 =>
                           n29113, A => n36145, ZN => n36138);
   U33972 : OAI222_X1 port map( A1 => n31437, A2 => n39184, B1 => n31501, B2 =>
                           n39178, C1 => n31373, C2 => n39172, ZN => n36145);
   U33973 : AOI221_X1 port map( B1 => n39076, B2 => n32511, C1 => n39070, C2 =>
                           n27949, A => n36134, ZN => n36127);
   U33974 : OAI222_X1 port map( A1 => n30550, A2 => n39064, B1 => n30614, B2 =>
                           n39058, C1 => n30486, C2 => n39052, ZN => n36134);
   U33975 : AOI221_X1 port map( B1 => n39196, B2 => n29048, C1 => n39190, C2 =>
                           n29112, A => n36126, ZN => n36119);
   U33976 : OAI222_X1 port map( A1 => n31436, A2 => n39184, B1 => n31500, B2 =>
                           n39178, C1 => n31372, C2 => n39172, ZN => n36126);
   U33977 : AOI221_X1 port map( B1 => n39076, B2 => n32510, C1 => n39070, C2 =>
                           n27948, A => n36115, ZN => n36108);
   U33978 : OAI222_X1 port map( A1 => n30549, A2 => n39064, B1 => n30613, B2 =>
                           n39058, C1 => n30485, C2 => n39052, ZN => n36115);
   U33979 : AOI221_X1 port map( B1 => n39196, B2 => n29047, C1 => n39190, C2 =>
                           n29111, A => n36107, ZN => n36100);
   U33980 : OAI222_X1 port map( A1 => n31435, A2 => n39184, B1 => n31499, B2 =>
                           n39178, C1 => n31371, C2 => n39172, ZN => n36107);
   U33981 : AOI221_X1 port map( B1 => n39579, B2 => n30480, C1 => n39573, C2 =>
                           n28007, A => n33481, ZN => n33457);
   U33982 : OAI222_X1 port map( A1 => n30608, A2 => n39567, B1 => n30672, B2 =>
                           n39561, C1 => n30544, C2 => n39555, ZN => n33481);
   U33983 : AOI221_X1 port map( B1 => n39699, B2 => n29106, C1 => n39693, C2 =>
                           n29170, A => n33453, ZN => n33429);
   U33984 : OAI222_X1 port map( A1 => n31494, A2 => n39687, B1 => n31558, B2 =>
                           n39681, C1 => n31430, C2 => n39675, ZN => n33453);
   U33985 : AOI221_X1 port map( B1 => n39327, B2 => n30480, C1 => n39321, C2 =>
                           n28007, A => n34755, ZN => n34731);
   U33986 : OAI222_X1 port map( A1 => n30608, A2 => n39315, B1 => n30672, B2 =>
                           n39309, C1 => n30544, C2 => n39303, ZN => n34755);
   U33987 : AOI221_X1 port map( B1 => n39447, B2 => n29106, C1 => n39441, C2 =>
                           n29170, A => n34727, ZN => n34703);
   U33988 : OAI222_X1 port map( A1 => n31494, A2 => n39435, B1 => n31558, B2 =>
                           n39429, C1 => n31430, C2 => n39423, ZN => n34727);
   U33989 : AOI221_X1 port map( B1 => n39579, B2 => n30479, C1 => n39573, C2 =>
                           n28006, A => n33503, ZN => n33496);
   U33990 : OAI222_X1 port map( A1 => n30607, A2 => n39567, B1 => n30671, B2 =>
                           n39561, C1 => n30543, C2 => n39555, ZN => n33503);
   U33991 : AOI221_X1 port map( B1 => n39699, B2 => n29105, C1 => n39693, C2 =>
                           n29169, A => n33495, ZN => n33488);
   U33992 : OAI222_X1 port map( A1 => n31493, A2 => n39687, B1 => n31557, B2 =>
                           n39681, C1 => n31429, C2 => n39675, ZN => n33495);
   U33993 : AOI221_X1 port map( B1 => n39327, B2 => n30479, C1 => n39321, C2 =>
                           n28006, A => n34777, ZN => n34770);
   U33994 : OAI222_X1 port map( A1 => n30607, A2 => n39315, B1 => n30671, B2 =>
                           n39309, C1 => n30543, C2 => n39303, ZN => n34777);
   U33995 : AOI221_X1 port map( B1 => n39447, B2 => n29105, C1 => n39441, C2 =>
                           n29169, A => n34769, ZN => n34762);
   U33996 : OAI222_X1 port map( A1 => n31493, A2 => n39435, B1 => n31557, B2 =>
                           n39429, C1 => n31429, C2 => n39423, ZN => n34769);
   U33997 : AOI221_X1 port map( B1 => n39579, B2 => n30478, C1 => n39573, C2 =>
                           n28005, A => n33522, ZN => n33515);
   U33998 : OAI222_X1 port map( A1 => n30606, A2 => n39567, B1 => n30670, B2 =>
                           n39561, C1 => n30542, C2 => n39555, ZN => n33522);
   U33999 : AOI221_X1 port map( B1 => n39699, B2 => n29104, C1 => n39693, C2 =>
                           n29168, A => n33514, ZN => n33507);
   U34000 : OAI222_X1 port map( A1 => n31492, A2 => n39687, B1 => n31556, B2 =>
                           n39681, C1 => n31428, C2 => n39675, ZN => n33514);
   U34001 : AOI221_X1 port map( B1 => n39327, B2 => n30478, C1 => n39321, C2 =>
                           n28005, A => n34796, ZN => n34789);
   U34002 : OAI222_X1 port map( A1 => n30606, A2 => n39315, B1 => n30670, B2 =>
                           n39309, C1 => n30542, C2 => n39303, ZN => n34796);
   U34003 : AOI221_X1 port map( B1 => n39447, B2 => n29104, C1 => n39441, C2 =>
                           n29168, A => n34788, ZN => n34781);
   U34004 : OAI222_X1 port map( A1 => n31492, A2 => n39435, B1 => n31556, B2 =>
                           n39429, C1 => n31428, C2 => n39423, ZN => n34788);
   U34005 : AOI221_X1 port map( B1 => n39579, B2 => n30477, C1 => n39573, C2 =>
                           n28004, A => n33541, ZN => n33534);
   U34006 : OAI222_X1 port map( A1 => n30605, A2 => n39567, B1 => n30669, B2 =>
                           n39561, C1 => n30541, C2 => n39555, ZN => n33541);
   U34007 : AOI221_X1 port map( B1 => n39699, B2 => n29103, C1 => n39693, C2 =>
                           n29167, A => n33533, ZN => n33526);
   U34008 : OAI222_X1 port map( A1 => n31491, A2 => n39687, B1 => n31555, B2 =>
                           n39681, C1 => n31427, C2 => n39675, ZN => n33533);
   U34009 : AOI221_X1 port map( B1 => n39327, B2 => n30477, C1 => n39321, C2 =>
                           n28004, A => n34815, ZN => n34808);
   U34010 : OAI222_X1 port map( A1 => n30605, A2 => n39315, B1 => n30669, B2 =>
                           n39309, C1 => n30541, C2 => n39303, ZN => n34815);
   U34011 : AOI221_X1 port map( B1 => n39447, B2 => n29103, C1 => n39441, C2 =>
                           n29167, A => n34807, ZN => n34800);
   U34012 : OAI222_X1 port map( A1 => n31491, A2 => n39435, B1 => n31555, B2 =>
                           n39429, C1 => n31427, C2 => n39423, ZN => n34807);
   U34013 : AOI221_X1 port map( B1 => n39578, B2 => n30476, C1 => n39572, C2 =>
                           n28003, A => n33560, ZN => n33553);
   U34014 : OAI222_X1 port map( A1 => n30604, A2 => n39566, B1 => n30668, B2 =>
                           n39560, C1 => n30540, C2 => n39554, ZN => n33560);
   U34015 : AOI221_X1 port map( B1 => n39698, B2 => n29102, C1 => n39692, C2 =>
                           n29166, A => n33552, ZN => n33545);
   U34016 : OAI222_X1 port map( A1 => n31490, A2 => n39686, B1 => n31554, B2 =>
                           n39680, C1 => n31426, C2 => n39674, ZN => n33552);
   U34017 : AOI221_X1 port map( B1 => n39326, B2 => n30476, C1 => n39320, C2 =>
                           n28003, A => n34834, ZN => n34827);
   U34018 : OAI222_X1 port map( A1 => n30604, A2 => n39314, B1 => n30668, B2 =>
                           n39308, C1 => n30540, C2 => n39302, ZN => n34834);
   U34019 : AOI221_X1 port map( B1 => n39446, B2 => n29102, C1 => n39440, C2 =>
                           n29166, A => n34826, ZN => n34819);
   U34020 : OAI222_X1 port map( A1 => n31490, A2 => n39434, B1 => n31554, B2 =>
                           n39428, C1 => n31426, C2 => n39422, ZN => n34826);
   U34021 : AOI221_X1 port map( B1 => n39578, B2 => n30475, C1 => n39572, C2 =>
                           n28002, A => n33579, ZN => n33572);
   U34022 : OAI222_X1 port map( A1 => n30603, A2 => n39566, B1 => n30667, B2 =>
                           n39560, C1 => n30539, C2 => n39554, ZN => n33579);
   U34023 : AOI221_X1 port map( B1 => n39698, B2 => n29101, C1 => n39692, C2 =>
                           n29165, A => n33571, ZN => n33564);
   U34024 : OAI222_X1 port map( A1 => n31489, A2 => n39686, B1 => n31553, B2 =>
                           n39680, C1 => n31425, C2 => n39674, ZN => n33571);
   U34025 : AOI221_X1 port map( B1 => n39326, B2 => n30475, C1 => n39320, C2 =>
                           n28002, A => n34853, ZN => n34846);
   U34026 : OAI222_X1 port map( A1 => n30603, A2 => n39314, B1 => n30667, B2 =>
                           n39308, C1 => n30539, C2 => n39302, ZN => n34853);
   U34027 : AOI221_X1 port map( B1 => n39446, B2 => n29101, C1 => n39440, C2 =>
                           n29165, A => n34845, ZN => n34838);
   U34028 : OAI222_X1 port map( A1 => n31489, A2 => n39434, B1 => n31553, B2 =>
                           n39428, C1 => n31425, C2 => n39422, ZN => n34845);
   U34029 : AOI221_X1 port map( B1 => n39578, B2 => n30474, C1 => n39572, C2 =>
                           n28001, A => n33598, ZN => n33591);
   U34030 : OAI222_X1 port map( A1 => n30602, A2 => n39566, B1 => n30666, B2 =>
                           n39560, C1 => n30538, C2 => n39554, ZN => n33598);
   U34031 : AOI221_X1 port map( B1 => n39698, B2 => n29100, C1 => n39692, C2 =>
                           n29164, A => n33590, ZN => n33583);
   U34032 : OAI222_X1 port map( A1 => n31488, A2 => n39686, B1 => n31552, B2 =>
                           n39680, C1 => n31424, C2 => n39674, ZN => n33590);
   U34033 : AOI221_X1 port map( B1 => n39326, B2 => n30474, C1 => n39320, C2 =>
                           n28001, A => n34872, ZN => n34865);
   U34034 : OAI222_X1 port map( A1 => n30602, A2 => n39314, B1 => n30666, B2 =>
                           n39308, C1 => n30538, C2 => n39302, ZN => n34872);
   U34035 : AOI221_X1 port map( B1 => n39446, B2 => n29100, C1 => n39440, C2 =>
                           n29164, A => n34864, ZN => n34857);
   U34036 : OAI222_X1 port map( A1 => n31488, A2 => n39434, B1 => n31552, B2 =>
                           n39428, C1 => n31424, C2 => n39422, ZN => n34864);
   U34037 : AOI221_X1 port map( B1 => n39578, B2 => n30473, C1 => n39572, C2 =>
                           n28000, A => n33617, ZN => n33610);
   U34038 : OAI222_X1 port map( A1 => n30601, A2 => n39566, B1 => n30665, B2 =>
                           n39560, C1 => n30537, C2 => n39554, ZN => n33617);
   U34039 : AOI221_X1 port map( B1 => n39698, B2 => n29099, C1 => n39692, C2 =>
                           n29163, A => n33609, ZN => n33602);
   U34040 : OAI222_X1 port map( A1 => n31487, A2 => n39686, B1 => n31551, B2 =>
                           n39680, C1 => n31423, C2 => n39674, ZN => n33609);
   U34041 : AOI221_X1 port map( B1 => n39326, B2 => n30473, C1 => n39320, C2 =>
                           n28000, A => n34891, ZN => n34884);
   U34042 : OAI222_X1 port map( A1 => n30601, A2 => n39314, B1 => n30665, B2 =>
                           n39308, C1 => n30537, C2 => n39302, ZN => n34891);
   U34043 : AOI221_X1 port map( B1 => n39446, B2 => n29099, C1 => n39440, C2 =>
                           n29163, A => n34883, ZN => n34876);
   U34044 : OAI222_X1 port map( A1 => n31487, A2 => n39434, B1 => n31551, B2 =>
                           n39428, C1 => n31423, C2 => n39422, ZN => n34883);
   U34045 : AOI221_X1 port map( B1 => n39578, B2 => n30472, C1 => n39572, C2 =>
                           n27999, A => n33636, ZN => n33629);
   U34046 : OAI222_X1 port map( A1 => n30600, A2 => n39566, B1 => n30664, B2 =>
                           n39560, C1 => n30536, C2 => n39554, ZN => n33636);
   U34047 : AOI221_X1 port map( B1 => n39698, B2 => n29098, C1 => n39692, C2 =>
                           n29162, A => n33628, ZN => n33621);
   U34048 : OAI222_X1 port map( A1 => n31486, A2 => n39686, B1 => n31550, B2 =>
                           n39680, C1 => n31422, C2 => n39674, ZN => n33628);
   U34049 : AOI221_X1 port map( B1 => n39326, B2 => n30472, C1 => n39320, C2 =>
                           n27999, A => n34910, ZN => n34903);
   U34050 : OAI222_X1 port map( A1 => n30600, A2 => n39314, B1 => n30664, B2 =>
                           n39308, C1 => n30536, C2 => n39302, ZN => n34910);
   U34051 : AOI221_X1 port map( B1 => n39446, B2 => n29098, C1 => n39440, C2 =>
                           n29162, A => n34902, ZN => n34895);
   U34052 : OAI222_X1 port map( A1 => n31486, A2 => n39434, B1 => n31550, B2 =>
                           n39428, C1 => n31422, C2 => n39422, ZN => n34902);
   U34053 : AOI221_X1 port map( B1 => n39578, B2 => n30471, C1 => n39572, C2 =>
                           n27998, A => n33655, ZN => n33648);
   U34054 : OAI222_X1 port map( A1 => n30599, A2 => n39566, B1 => n30663, B2 =>
                           n39560, C1 => n30535, C2 => n39554, ZN => n33655);
   U34055 : AOI221_X1 port map( B1 => n39698, B2 => n29097, C1 => n39692, C2 =>
                           n29161, A => n33647, ZN => n33640);
   U34056 : OAI222_X1 port map( A1 => n31485, A2 => n39686, B1 => n31549, B2 =>
                           n39680, C1 => n31421, C2 => n39674, ZN => n33647);
   U34057 : AOI221_X1 port map( B1 => n39326, B2 => n30471, C1 => n39320, C2 =>
                           n27998, A => n34929, ZN => n34922);
   U34058 : OAI222_X1 port map( A1 => n30599, A2 => n39314, B1 => n30663, B2 =>
                           n39308, C1 => n30535, C2 => n39302, ZN => n34929);
   U34059 : AOI221_X1 port map( B1 => n39446, B2 => n29097, C1 => n39440, C2 =>
                           n29161, A => n34921, ZN => n34914);
   U34060 : OAI222_X1 port map( A1 => n31485, A2 => n39434, B1 => n31549, B2 =>
                           n39428, C1 => n31421, C2 => n39422, ZN => n34921);
   U34061 : AOI221_X1 port map( B1 => n39578, B2 => n30470, C1 => n39572, C2 =>
                           n27997, A => n33674, ZN => n33667);
   U34062 : OAI222_X1 port map( A1 => n30598, A2 => n39566, B1 => n30662, B2 =>
                           n39560, C1 => n30534, C2 => n39554, ZN => n33674);
   U34063 : AOI221_X1 port map( B1 => n39698, B2 => n29096, C1 => n39692, C2 =>
                           n29160, A => n33666, ZN => n33659);
   U34064 : OAI222_X1 port map( A1 => n31484, A2 => n39686, B1 => n31548, B2 =>
                           n39680, C1 => n31420, C2 => n39674, ZN => n33666);
   U34065 : AOI221_X1 port map( B1 => n39326, B2 => n30470, C1 => n39320, C2 =>
                           n27997, A => n34948, ZN => n34941);
   U34066 : OAI222_X1 port map( A1 => n30598, A2 => n39314, B1 => n30662, B2 =>
                           n39308, C1 => n30534, C2 => n39302, ZN => n34948);
   U34067 : AOI221_X1 port map( B1 => n39446, B2 => n29096, C1 => n39440, C2 =>
                           n29160, A => n34940, ZN => n34933);
   U34068 : OAI222_X1 port map( A1 => n31484, A2 => n39434, B1 => n31548, B2 =>
                           n39428, C1 => n31420, C2 => n39422, ZN => n34940);
   U34069 : AOI221_X1 port map( B1 => n39578, B2 => n30469, C1 => n39572, C2 =>
                           n27996, A => n33693, ZN => n33686);
   U34070 : OAI222_X1 port map( A1 => n30597, A2 => n39566, B1 => n30661, B2 =>
                           n39560, C1 => n30533, C2 => n39554, ZN => n33693);
   U34071 : AOI221_X1 port map( B1 => n39698, B2 => n29095, C1 => n39692, C2 =>
                           n29159, A => n33685, ZN => n33678);
   U34072 : OAI222_X1 port map( A1 => n31483, A2 => n39686, B1 => n31547, B2 =>
                           n39680, C1 => n31419, C2 => n39674, ZN => n33685);
   U34073 : AOI221_X1 port map( B1 => n39326, B2 => n30469, C1 => n39320, C2 =>
                           n27996, A => n34967, ZN => n34960);
   U34074 : OAI222_X1 port map( A1 => n30597, A2 => n39314, B1 => n30661, B2 =>
                           n39308, C1 => n30533, C2 => n39302, ZN => n34967);
   U34075 : AOI221_X1 port map( B1 => n39446, B2 => n29095, C1 => n39440, C2 =>
                           n29159, A => n34959, ZN => n34952);
   U34076 : OAI222_X1 port map( A1 => n31483, A2 => n39434, B1 => n31547, B2 =>
                           n39428, C1 => n31419, C2 => n39422, ZN => n34959);
   U34077 : AOI221_X1 port map( B1 => n39578, B2 => n30468, C1 => n39572, C2 =>
                           n27995, A => n33712, ZN => n33705);
   U34078 : OAI222_X1 port map( A1 => n30596, A2 => n39566, B1 => n30660, B2 =>
                           n39560, C1 => n30532, C2 => n39554, ZN => n33712);
   U34079 : AOI221_X1 port map( B1 => n39698, B2 => n29094, C1 => n39692, C2 =>
                           n29158, A => n33704, ZN => n33697);
   U34080 : OAI222_X1 port map( A1 => n31482, A2 => n39686, B1 => n31546, B2 =>
                           n39680, C1 => n31418, C2 => n39674, ZN => n33704);
   U34081 : AOI221_X1 port map( B1 => n39326, B2 => n30468, C1 => n39320, C2 =>
                           n27995, A => n34986, ZN => n34979);
   U34082 : OAI222_X1 port map( A1 => n30596, A2 => n39314, B1 => n30660, B2 =>
                           n39308, C1 => n30532, C2 => n39302, ZN => n34986);
   U34083 : AOI221_X1 port map( B1 => n39446, B2 => n29094, C1 => n39440, C2 =>
                           n29158, A => n34978, ZN => n34971);
   U34084 : OAI222_X1 port map( A1 => n31482, A2 => n39434, B1 => n31546, B2 =>
                           n39428, C1 => n31418, C2 => n39422, ZN => n34978);
   U34085 : AOI221_X1 port map( B1 => n39578, B2 => n30467, C1 => n39572, C2 =>
                           n27994, A => n33731, ZN => n33724);
   U34086 : OAI222_X1 port map( A1 => n30595, A2 => n39566, B1 => n30659, B2 =>
                           n39560, C1 => n30531, C2 => n39554, ZN => n33731);
   U34087 : AOI221_X1 port map( B1 => n39698, B2 => n29093, C1 => n39692, C2 =>
                           n29157, A => n33723, ZN => n33716);
   U34088 : OAI222_X1 port map( A1 => n31481, A2 => n39686, B1 => n31545, B2 =>
                           n39680, C1 => n31417, C2 => n39674, ZN => n33723);
   U34089 : AOI221_X1 port map( B1 => n39326, B2 => n30467, C1 => n39320, C2 =>
                           n27994, A => n35005, ZN => n34998);
   U34090 : OAI222_X1 port map( A1 => n30595, A2 => n39314, B1 => n30659, B2 =>
                           n39308, C1 => n30531, C2 => n39302, ZN => n35005);
   U34091 : AOI221_X1 port map( B1 => n39446, B2 => n29093, C1 => n39440, C2 =>
                           n29157, A => n34997, ZN => n34990);
   U34092 : OAI222_X1 port map( A1 => n31481, A2 => n39434, B1 => n31545, B2 =>
                           n39428, C1 => n31417, C2 => n39422, ZN => n34997);
   U34093 : AOI221_X1 port map( B1 => n39578, B2 => n30466, C1 => n39572, C2 =>
                           n27993, A => n33750, ZN => n33743);
   U34094 : OAI222_X1 port map( A1 => n30594, A2 => n39566, B1 => n30658, B2 =>
                           n39560, C1 => n30530, C2 => n39554, ZN => n33750);
   U34095 : AOI221_X1 port map( B1 => n39698, B2 => n29092, C1 => n39692, C2 =>
                           n29156, A => n33742, ZN => n33735);
   U34096 : OAI222_X1 port map( A1 => n31480, A2 => n39686, B1 => n31544, B2 =>
                           n39680, C1 => n31416, C2 => n39674, ZN => n33742);
   U34097 : AOI221_X1 port map( B1 => n39326, B2 => n30466, C1 => n39320, C2 =>
                           n27993, A => n35024, ZN => n35017);
   U34098 : OAI222_X1 port map( A1 => n30594, A2 => n39314, B1 => n30658, B2 =>
                           n39308, C1 => n30530, C2 => n39302, ZN => n35024);
   U34099 : AOI221_X1 port map( B1 => n39446, B2 => n29092, C1 => n39440, C2 =>
                           n29156, A => n35016, ZN => n35009);
   U34100 : OAI222_X1 port map( A1 => n31480, A2 => n39434, B1 => n31544, B2 =>
                           n39428, C1 => n31416, C2 => n39422, ZN => n35016);
   U34101 : AOI221_X1 port map( B1 => n39578, B2 => n30465, C1 => n39572, C2 =>
                           n27992, A => n33769, ZN => n33762);
   U34102 : OAI222_X1 port map( A1 => n30593, A2 => n39566, B1 => n30657, B2 =>
                           n39560, C1 => n30529, C2 => n39554, ZN => n33769);
   U34103 : AOI221_X1 port map( B1 => n39698, B2 => n29091, C1 => n39692, C2 =>
                           n29155, A => n33761, ZN => n33754);
   U34104 : OAI222_X1 port map( A1 => n31479, A2 => n39686, B1 => n31543, B2 =>
                           n39680, C1 => n31415, C2 => n39674, ZN => n33761);
   U34105 : AOI221_X1 port map( B1 => n39326, B2 => n30465, C1 => n39320, C2 =>
                           n27992, A => n35043, ZN => n35036);
   U34106 : OAI222_X1 port map( A1 => n30593, A2 => n39314, B1 => n30657, B2 =>
                           n39308, C1 => n30529, C2 => n39302, ZN => n35043);
   U34107 : AOI221_X1 port map( B1 => n39446, B2 => n29091, C1 => n39440, C2 =>
                           n29155, A => n35035, ZN => n35028);
   U34108 : OAI222_X1 port map( A1 => n31479, A2 => n39434, B1 => n31543, B2 =>
                           n39428, C1 => n31415, C2 => n39422, ZN => n35035);
   U34109 : AOI221_X1 port map( B1 => n39577, B2 => n30464, C1 => n39571, C2 =>
                           n27991, A => n33788, ZN => n33781);
   U34110 : OAI222_X1 port map( A1 => n30592, A2 => n39565, B1 => n30656, B2 =>
                           n39559, C1 => n30528, C2 => n39553, ZN => n33788);
   U34111 : AOI221_X1 port map( B1 => n39697, B2 => n29090, C1 => n39691, C2 =>
                           n29154, A => n33780, ZN => n33773);
   U34112 : OAI222_X1 port map( A1 => n31478, A2 => n39685, B1 => n31542, B2 =>
                           n39679, C1 => n31414, C2 => n39673, ZN => n33780);
   U34113 : AOI221_X1 port map( B1 => n39325, B2 => n30464, C1 => n39319, C2 =>
                           n27991, A => n35062, ZN => n35055);
   U34114 : OAI222_X1 port map( A1 => n30592, A2 => n39313, B1 => n30656, B2 =>
                           n39307, C1 => n30528, C2 => n39301, ZN => n35062);
   U34115 : AOI221_X1 port map( B1 => n39445, B2 => n29090, C1 => n39439, C2 =>
                           n29154, A => n35054, ZN => n35047);
   U34116 : OAI222_X1 port map( A1 => n31478, A2 => n39433, B1 => n31542, B2 =>
                           n39427, C1 => n31414, C2 => n39421, ZN => n35054);
   U34117 : AOI221_X1 port map( B1 => n39577, B2 => n30463, C1 => n39571, C2 =>
                           n27990, A => n33807, ZN => n33800);
   U34118 : OAI222_X1 port map( A1 => n30591, A2 => n39565, B1 => n30655, B2 =>
                           n39559, C1 => n30527, C2 => n39553, ZN => n33807);
   U34119 : AOI221_X1 port map( B1 => n39697, B2 => n29089, C1 => n39691, C2 =>
                           n29153, A => n33799, ZN => n33792);
   U34120 : OAI222_X1 port map( A1 => n31477, A2 => n39685, B1 => n31541, B2 =>
                           n39679, C1 => n31413, C2 => n39673, ZN => n33799);
   U34121 : AOI221_X1 port map( B1 => n39325, B2 => n30463, C1 => n39319, C2 =>
                           n27990, A => n35081, ZN => n35074);
   U34122 : OAI222_X1 port map( A1 => n30591, A2 => n39313, B1 => n30655, B2 =>
                           n39307, C1 => n30527, C2 => n39301, ZN => n35081);
   U34123 : AOI221_X1 port map( B1 => n39445, B2 => n29089, C1 => n39439, C2 =>
                           n29153, A => n35073, ZN => n35066);
   U34124 : OAI222_X1 port map( A1 => n31477, A2 => n39433, B1 => n31541, B2 =>
                           n39427, C1 => n31413, C2 => n39421, ZN => n35073);
   U34125 : AOI221_X1 port map( B1 => n39577, B2 => n30462, C1 => n39571, C2 =>
                           n27989, A => n33826, ZN => n33819);
   U34126 : OAI222_X1 port map( A1 => n30590, A2 => n39565, B1 => n30654, B2 =>
                           n39559, C1 => n30526, C2 => n39553, ZN => n33826);
   U34127 : AOI221_X1 port map( B1 => n39697, B2 => n29088, C1 => n39691, C2 =>
                           n29152, A => n33818, ZN => n33811);
   U34128 : OAI222_X1 port map( A1 => n31476, A2 => n39685, B1 => n31540, B2 =>
                           n39679, C1 => n31412, C2 => n39673, ZN => n33818);
   U34129 : AOI221_X1 port map( B1 => n39325, B2 => n30462, C1 => n39319, C2 =>
                           n27989, A => n35100, ZN => n35093);
   U34130 : OAI222_X1 port map( A1 => n30590, A2 => n39313, B1 => n30654, B2 =>
                           n39307, C1 => n30526, C2 => n39301, ZN => n35100);
   U34131 : AOI221_X1 port map( B1 => n39445, B2 => n29088, C1 => n39439, C2 =>
                           n29152, A => n35092, ZN => n35085);
   U34132 : OAI222_X1 port map( A1 => n31476, A2 => n39433, B1 => n31540, B2 =>
                           n39427, C1 => n31412, C2 => n39421, ZN => n35092);
   U34133 : AOI221_X1 port map( B1 => n39577, B2 => n30461, C1 => n39571, C2 =>
                           n27988, A => n33845, ZN => n33838);
   U34134 : OAI222_X1 port map( A1 => n30589, A2 => n39565, B1 => n30653, B2 =>
                           n39559, C1 => n30525, C2 => n39553, ZN => n33845);
   U34135 : AOI221_X1 port map( B1 => n39697, B2 => n29087, C1 => n39691, C2 =>
                           n29151, A => n33837, ZN => n33830);
   U34136 : OAI222_X1 port map( A1 => n31475, A2 => n39685, B1 => n31539, B2 =>
                           n39679, C1 => n31411, C2 => n39673, ZN => n33837);
   U34137 : AOI221_X1 port map( B1 => n39325, B2 => n30461, C1 => n39319, C2 =>
                           n27988, A => n35119, ZN => n35112);
   U34138 : OAI222_X1 port map( A1 => n30589, A2 => n39313, B1 => n30653, B2 =>
                           n39307, C1 => n30525, C2 => n39301, ZN => n35119);
   U34139 : AOI221_X1 port map( B1 => n39445, B2 => n29087, C1 => n39439, C2 =>
                           n29151, A => n35111, ZN => n35104);
   U34140 : OAI222_X1 port map( A1 => n31475, A2 => n39433, B1 => n31539, B2 =>
                           n39427, C1 => n31411, C2 => n39421, ZN => n35111);
   U34141 : AOI221_X1 port map( B1 => n39577, B2 => n30460, C1 => n39571, C2 =>
                           n27987, A => n33864, ZN => n33857);
   U34142 : OAI222_X1 port map( A1 => n30588, A2 => n39565, B1 => n30652, B2 =>
                           n39559, C1 => n30524, C2 => n39553, ZN => n33864);
   U34143 : AOI221_X1 port map( B1 => n39697, B2 => n29086, C1 => n39691, C2 =>
                           n29150, A => n33856, ZN => n33849);
   U34144 : OAI222_X1 port map( A1 => n31474, A2 => n39685, B1 => n31538, B2 =>
                           n39679, C1 => n31410, C2 => n39673, ZN => n33856);
   U34145 : AOI221_X1 port map( B1 => n39325, B2 => n30460, C1 => n39319, C2 =>
                           n27987, A => n35138, ZN => n35131);
   U34146 : OAI222_X1 port map( A1 => n30588, A2 => n39313, B1 => n30652, B2 =>
                           n39307, C1 => n30524, C2 => n39301, ZN => n35138);
   U34147 : AOI221_X1 port map( B1 => n39445, B2 => n29086, C1 => n39439, C2 =>
                           n29150, A => n35130, ZN => n35123);
   U34148 : OAI222_X1 port map( A1 => n31474, A2 => n39433, B1 => n31538, B2 =>
                           n39427, C1 => n31410, C2 => n39421, ZN => n35130);
   U34149 : AOI221_X1 port map( B1 => n39577, B2 => n30459, C1 => n39571, C2 =>
                           n27986, A => n33883, ZN => n33876);
   U34150 : OAI222_X1 port map( A1 => n30587, A2 => n39565, B1 => n30651, B2 =>
                           n39559, C1 => n30523, C2 => n39553, ZN => n33883);
   U34151 : AOI221_X1 port map( B1 => n39697, B2 => n29085, C1 => n39691, C2 =>
                           n29149, A => n33875, ZN => n33868);
   U34152 : OAI222_X1 port map( A1 => n31473, A2 => n39685, B1 => n31537, B2 =>
                           n39679, C1 => n31409, C2 => n39673, ZN => n33875);
   U34153 : AOI221_X1 port map( B1 => n39325, B2 => n30459, C1 => n39319, C2 =>
                           n27986, A => n35157, ZN => n35150);
   U34154 : OAI222_X1 port map( A1 => n30587, A2 => n39313, B1 => n30651, B2 =>
                           n39307, C1 => n30523, C2 => n39301, ZN => n35157);
   U34155 : AOI221_X1 port map( B1 => n39445, B2 => n29085, C1 => n39439, C2 =>
                           n29149, A => n35149, ZN => n35142);
   U34156 : OAI222_X1 port map( A1 => n31473, A2 => n39433, B1 => n31537, B2 =>
                           n39427, C1 => n31409, C2 => n39421, ZN => n35149);
   U34157 : AOI221_X1 port map( B1 => n39577, B2 => n30458, C1 => n39571, C2 =>
                           n27985, A => n33902, ZN => n33895);
   U34158 : OAI222_X1 port map( A1 => n30586, A2 => n39565, B1 => n30650, B2 =>
                           n39559, C1 => n30522, C2 => n39553, ZN => n33902);
   U34159 : AOI221_X1 port map( B1 => n39697, B2 => n29084, C1 => n39691, C2 =>
                           n29148, A => n33894, ZN => n33887);
   U34160 : OAI222_X1 port map( A1 => n31472, A2 => n39685, B1 => n31536, B2 =>
                           n39679, C1 => n31408, C2 => n39673, ZN => n33894);
   U34161 : AOI221_X1 port map( B1 => n39325, B2 => n30458, C1 => n39319, C2 =>
                           n27985, A => n35176, ZN => n35169);
   U34162 : OAI222_X1 port map( A1 => n30586, A2 => n39313, B1 => n30650, B2 =>
                           n39307, C1 => n30522, C2 => n39301, ZN => n35176);
   U34163 : AOI221_X1 port map( B1 => n39445, B2 => n29084, C1 => n39439, C2 =>
                           n29148, A => n35168, ZN => n35161);
   U34164 : OAI222_X1 port map( A1 => n31472, A2 => n39433, B1 => n31536, B2 =>
                           n39427, C1 => n31408, C2 => n39421, ZN => n35168);
   U34165 : AOI221_X1 port map( B1 => n39577, B2 => n32546, C1 => n39571, C2 =>
                           n27984, A => n33921, ZN => n33914);
   U34166 : OAI222_X1 port map( A1 => n30585, A2 => n39565, B1 => n30649, B2 =>
                           n39559, C1 => n30521, C2 => n39553, ZN => n33921);
   U34167 : AOI221_X1 port map( B1 => n39697, B2 => n29083, C1 => n39691, C2 =>
                           n29147, A => n33913, ZN => n33906);
   U34168 : OAI222_X1 port map( A1 => n31471, A2 => n39685, B1 => n31535, B2 =>
                           n39679, C1 => n31407, C2 => n39673, ZN => n33913);
   U34169 : AOI221_X1 port map( B1 => n39325, B2 => n32546, C1 => n39319, C2 =>
                           n27984, A => n35195, ZN => n35188);
   U34170 : OAI222_X1 port map( A1 => n30585, A2 => n39313, B1 => n30649, B2 =>
                           n39307, C1 => n30521, C2 => n39301, ZN => n35195);
   U34171 : AOI221_X1 port map( B1 => n39445, B2 => n29083, C1 => n39439, C2 =>
                           n29147, A => n35187, ZN => n35180);
   U34172 : OAI222_X1 port map( A1 => n31471, A2 => n39433, B1 => n31535, B2 =>
                           n39427, C1 => n31407, C2 => n39421, ZN => n35187);
   U34173 : AOI221_X1 port map( B1 => n39577, B2 => n32545, C1 => n39571, C2 =>
                           n27983, A => n33940, ZN => n33933);
   U34174 : OAI222_X1 port map( A1 => n30584, A2 => n39565, B1 => n30648, B2 =>
                           n39559, C1 => n30520, C2 => n39553, ZN => n33940);
   U34175 : AOI221_X1 port map( B1 => n39697, B2 => n29082, C1 => n39691, C2 =>
                           n29146, A => n33932, ZN => n33925);
   U34176 : OAI222_X1 port map( A1 => n31470, A2 => n39685, B1 => n31534, B2 =>
                           n39679, C1 => n31406, C2 => n39673, ZN => n33932);
   U34177 : AOI221_X1 port map( B1 => n39325, B2 => n32545, C1 => n39319, C2 =>
                           n27983, A => n35214, ZN => n35207);
   U34178 : OAI222_X1 port map( A1 => n30584, A2 => n39313, B1 => n30648, B2 =>
                           n39307, C1 => n30520, C2 => n39301, ZN => n35214);
   U34179 : AOI221_X1 port map( B1 => n39445, B2 => n29082, C1 => n39439, C2 =>
                           n29146, A => n35206, ZN => n35199);
   U34180 : OAI222_X1 port map( A1 => n31470, A2 => n39433, B1 => n31534, B2 =>
                           n39427, C1 => n31406, C2 => n39421, ZN => n35206);
   U34181 : AOI221_X1 port map( B1 => n39577, B2 => n32544, C1 => n39571, C2 =>
                           n27982, A => n33959, ZN => n33952);
   U34182 : OAI222_X1 port map( A1 => n30583, A2 => n39565, B1 => n30647, B2 =>
                           n39559, C1 => n30519, C2 => n39553, ZN => n33959);
   U34183 : AOI221_X1 port map( B1 => n39697, B2 => n29081, C1 => n39691, C2 =>
                           n29145, A => n33951, ZN => n33944);
   U34184 : OAI222_X1 port map( A1 => n31469, A2 => n39685, B1 => n31533, B2 =>
                           n39679, C1 => n31405, C2 => n39673, ZN => n33951);
   U34185 : AOI221_X1 port map( B1 => n39325, B2 => n32544, C1 => n39319, C2 =>
                           n27982, A => n35233, ZN => n35226);
   U34186 : OAI222_X1 port map( A1 => n30583, A2 => n39313, B1 => n30647, B2 =>
                           n39307, C1 => n30519, C2 => n39301, ZN => n35233);
   U34187 : AOI221_X1 port map( B1 => n39445, B2 => n29081, C1 => n39439, C2 =>
                           n29145, A => n35225, ZN => n35218);
   U34188 : OAI222_X1 port map( A1 => n31469, A2 => n39433, B1 => n31533, B2 =>
                           n39427, C1 => n31405, C2 => n39421, ZN => n35225);
   U34189 : AOI221_X1 port map( B1 => n39577, B2 => n32543, C1 => n39571, C2 =>
                           n27981, A => n33978, ZN => n33971);
   U34190 : OAI222_X1 port map( A1 => n30582, A2 => n39565, B1 => n30646, B2 =>
                           n39559, C1 => n30518, C2 => n39553, ZN => n33978);
   U34191 : AOI221_X1 port map( B1 => n39697, B2 => n29080, C1 => n39691, C2 =>
                           n29144, A => n33970, ZN => n33963);
   U34192 : OAI222_X1 port map( A1 => n31468, A2 => n39685, B1 => n31532, B2 =>
                           n39679, C1 => n31404, C2 => n39673, ZN => n33970);
   U34193 : AOI221_X1 port map( B1 => n39325, B2 => n32543, C1 => n39319, C2 =>
                           n27981, A => n35252, ZN => n35245);
   U34194 : OAI222_X1 port map( A1 => n30582, A2 => n39313, B1 => n30646, B2 =>
                           n39307, C1 => n30518, C2 => n39301, ZN => n35252);
   U34195 : AOI221_X1 port map( B1 => n39445, B2 => n29080, C1 => n39439, C2 =>
                           n29144, A => n35244, ZN => n35237);
   U34196 : OAI222_X1 port map( A1 => n31468, A2 => n39433, B1 => n31532, B2 =>
                           n39427, C1 => n31404, C2 => n39421, ZN => n35244);
   U34197 : AOI221_X1 port map( B1 => n39577, B2 => n32542, C1 => n39571, C2 =>
                           n27980, A => n33997, ZN => n33990);
   U34198 : OAI222_X1 port map( A1 => n30581, A2 => n39565, B1 => n30645, B2 =>
                           n39559, C1 => n30517, C2 => n39553, ZN => n33997);
   U34199 : AOI221_X1 port map( B1 => n39697, B2 => n29079, C1 => n39691, C2 =>
                           n29143, A => n33989, ZN => n33982);
   U34200 : OAI222_X1 port map( A1 => n31467, A2 => n39685, B1 => n31531, B2 =>
                           n39679, C1 => n31403, C2 => n39673, ZN => n33989);
   U34201 : AOI221_X1 port map( B1 => n39325, B2 => n32542, C1 => n39319, C2 =>
                           n27980, A => n35271, ZN => n35264);
   U34202 : OAI222_X1 port map( A1 => n30581, A2 => n39313, B1 => n30645, B2 =>
                           n39307, C1 => n30517, C2 => n39301, ZN => n35271);
   U34203 : AOI221_X1 port map( B1 => n39445, B2 => n29079, C1 => n39439, C2 =>
                           n29143, A => n35263, ZN => n35256);
   U34204 : OAI222_X1 port map( A1 => n31467, A2 => n39433, B1 => n31531, B2 =>
                           n39427, C1 => n31403, C2 => n39421, ZN => n35263);
   U34205 : AOI221_X1 port map( B1 => n39576, B2 => n32541, C1 => n39570, C2 =>
                           n27979, A => n34016, ZN => n34009);
   U34206 : OAI222_X1 port map( A1 => n30580, A2 => n39564, B1 => n30644, B2 =>
                           n39558, C1 => n30516, C2 => n39552, ZN => n34016);
   U34207 : AOI221_X1 port map( B1 => n39696, B2 => n29078, C1 => n39690, C2 =>
                           n29142, A => n34008, ZN => n34001);
   U34208 : OAI222_X1 port map( A1 => n31466, A2 => n39684, B1 => n31530, B2 =>
                           n39678, C1 => n31402, C2 => n39672, ZN => n34008);
   U34209 : AOI221_X1 port map( B1 => n39324, B2 => n32541, C1 => n39318, C2 =>
                           n27979, A => n35290, ZN => n35283);
   U34210 : OAI222_X1 port map( A1 => n30580, A2 => n39312, B1 => n30644, B2 =>
                           n39306, C1 => n30516, C2 => n39300, ZN => n35290);
   U34211 : AOI221_X1 port map( B1 => n39444, B2 => n29078, C1 => n39438, C2 =>
                           n29142, A => n35282, ZN => n35275);
   U34212 : OAI222_X1 port map( A1 => n31466, A2 => n39432, B1 => n31530, B2 =>
                           n39426, C1 => n31402, C2 => n39420, ZN => n35282);
   U34213 : AOI221_X1 port map( B1 => n39576, B2 => n32540, C1 => n39570, C2 =>
                           n27978, A => n34035, ZN => n34028);
   U34214 : OAI222_X1 port map( A1 => n30579, A2 => n39564, B1 => n30643, B2 =>
                           n39558, C1 => n30515, C2 => n39552, ZN => n34035);
   U34215 : AOI221_X1 port map( B1 => n39696, B2 => n29077, C1 => n39690, C2 =>
                           n29141, A => n34027, ZN => n34020);
   U34216 : OAI222_X1 port map( A1 => n31465, A2 => n39684, B1 => n31529, B2 =>
                           n39678, C1 => n31401, C2 => n39672, ZN => n34027);
   U34217 : AOI221_X1 port map( B1 => n39324, B2 => n32540, C1 => n39318, C2 =>
                           n27978, A => n35309, ZN => n35302);
   U34218 : OAI222_X1 port map( A1 => n30579, A2 => n39312, B1 => n30643, B2 =>
                           n39306, C1 => n30515, C2 => n39300, ZN => n35309);
   U34219 : AOI221_X1 port map( B1 => n39444, B2 => n29077, C1 => n39438, C2 =>
                           n29141, A => n35301, ZN => n35294);
   U34220 : OAI222_X1 port map( A1 => n31465, A2 => n39432, B1 => n31529, B2 =>
                           n39426, C1 => n31401, C2 => n39420, ZN => n35301);
   U34221 : AOI221_X1 port map( B1 => n39576, B2 => n32539, C1 => n39570, C2 =>
                           n27977, A => n34054, ZN => n34047);
   U34222 : OAI222_X1 port map( A1 => n30578, A2 => n39564, B1 => n30642, B2 =>
                           n39558, C1 => n30514, C2 => n39552, ZN => n34054);
   U34223 : AOI221_X1 port map( B1 => n39696, B2 => n29076, C1 => n39690, C2 =>
                           n29140, A => n34046, ZN => n34039);
   U34224 : OAI222_X1 port map( A1 => n31464, A2 => n39684, B1 => n31528, B2 =>
                           n39678, C1 => n31400, C2 => n39672, ZN => n34046);
   U34225 : AOI221_X1 port map( B1 => n39324, B2 => n32539, C1 => n39318, C2 =>
                           n27977, A => n35328, ZN => n35321);
   U34226 : OAI222_X1 port map( A1 => n30578, A2 => n39312, B1 => n30642, B2 =>
                           n39306, C1 => n30514, C2 => n39300, ZN => n35328);
   U34227 : AOI221_X1 port map( B1 => n39444, B2 => n29076, C1 => n39438, C2 =>
                           n29140, A => n35320, ZN => n35313);
   U34228 : OAI222_X1 port map( A1 => n31464, A2 => n39432, B1 => n31528, B2 =>
                           n39426, C1 => n31400, C2 => n39420, ZN => n35320);
   U34229 : AOI221_X1 port map( B1 => n39576, B2 => n32538, C1 => n39570, C2 =>
                           n27976, A => n34073, ZN => n34066);
   U34230 : OAI222_X1 port map( A1 => n30577, A2 => n39564, B1 => n30641, B2 =>
                           n39558, C1 => n30513, C2 => n39552, ZN => n34073);
   U34231 : AOI221_X1 port map( B1 => n39696, B2 => n29075, C1 => n39690, C2 =>
                           n29139, A => n34065, ZN => n34058);
   U34232 : OAI222_X1 port map( A1 => n31463, A2 => n39684, B1 => n31527, B2 =>
                           n39678, C1 => n31399, C2 => n39672, ZN => n34065);
   U34233 : AOI221_X1 port map( B1 => n39324, B2 => n32538, C1 => n39318, C2 =>
                           n27976, A => n35347, ZN => n35340);
   U34234 : OAI222_X1 port map( A1 => n30577, A2 => n39312, B1 => n30641, B2 =>
                           n39306, C1 => n30513, C2 => n39300, ZN => n35347);
   U34235 : AOI221_X1 port map( B1 => n39444, B2 => n29075, C1 => n39438, C2 =>
                           n29139, A => n35339, ZN => n35332);
   U34236 : OAI222_X1 port map( A1 => n31463, A2 => n39432, B1 => n31527, B2 =>
                           n39426, C1 => n31399, C2 => n39420, ZN => n35339);
   U34237 : AOI221_X1 port map( B1 => n39576, B2 => n32537, C1 => n39570, C2 =>
                           n27975, A => n34092, ZN => n34085);
   U34238 : OAI222_X1 port map( A1 => n30576, A2 => n39564, B1 => n30640, B2 =>
                           n39558, C1 => n30512, C2 => n39552, ZN => n34092);
   U34239 : AOI221_X1 port map( B1 => n39696, B2 => n29074, C1 => n39690, C2 =>
                           n29138, A => n34084, ZN => n34077);
   U34240 : OAI222_X1 port map( A1 => n31462, A2 => n39684, B1 => n31526, B2 =>
                           n39678, C1 => n31398, C2 => n39672, ZN => n34084);
   U34241 : AOI221_X1 port map( B1 => n39324, B2 => n32537, C1 => n39318, C2 =>
                           n27975, A => n35366, ZN => n35359);
   U34242 : OAI222_X1 port map( A1 => n30576, A2 => n39312, B1 => n30640, B2 =>
                           n39306, C1 => n30512, C2 => n39300, ZN => n35366);
   U34243 : AOI221_X1 port map( B1 => n39444, B2 => n29074, C1 => n39438, C2 =>
                           n29138, A => n35358, ZN => n35351);
   U34244 : OAI222_X1 port map( A1 => n31462, A2 => n39432, B1 => n31526, B2 =>
                           n39426, C1 => n31398, C2 => n39420, ZN => n35358);
   U34245 : AOI221_X1 port map( B1 => n39576, B2 => n32536, C1 => n39570, C2 =>
                           n27974, A => n34111, ZN => n34104);
   U34246 : OAI222_X1 port map( A1 => n30575, A2 => n39564, B1 => n30639, B2 =>
                           n39558, C1 => n30511, C2 => n39552, ZN => n34111);
   U34247 : AOI221_X1 port map( B1 => n39696, B2 => n29073, C1 => n39690, C2 =>
                           n29137, A => n34103, ZN => n34096);
   U34248 : OAI222_X1 port map( A1 => n31461, A2 => n39684, B1 => n31525, B2 =>
                           n39678, C1 => n31397, C2 => n39672, ZN => n34103);
   U34249 : AOI221_X1 port map( B1 => n39324, B2 => n32536, C1 => n39318, C2 =>
                           n27974, A => n35385, ZN => n35378);
   U34250 : OAI222_X1 port map( A1 => n30575, A2 => n39312, B1 => n30639, B2 =>
                           n39306, C1 => n30511, C2 => n39300, ZN => n35385);
   U34251 : AOI221_X1 port map( B1 => n39444, B2 => n29073, C1 => n39438, C2 =>
                           n29137, A => n35377, ZN => n35370);
   U34252 : OAI222_X1 port map( A1 => n31461, A2 => n39432, B1 => n31525, B2 =>
                           n39426, C1 => n31397, C2 => n39420, ZN => n35377);
   U34253 : AOI221_X1 port map( B1 => n39576, B2 => n32535, C1 => n39570, C2 =>
                           n27973, A => n34130, ZN => n34123);
   U34254 : OAI222_X1 port map( A1 => n30574, A2 => n39564, B1 => n30638, B2 =>
                           n39558, C1 => n30510, C2 => n39552, ZN => n34130);
   U34255 : AOI221_X1 port map( B1 => n39696, B2 => n29072, C1 => n39690, C2 =>
                           n29136, A => n34122, ZN => n34115);
   U34256 : OAI222_X1 port map( A1 => n31460, A2 => n39684, B1 => n31524, B2 =>
                           n39678, C1 => n31396, C2 => n39672, ZN => n34122);
   U34257 : AOI221_X1 port map( B1 => n39324, B2 => n32535, C1 => n39318, C2 =>
                           n27973, A => n35404, ZN => n35397);
   U34258 : OAI222_X1 port map( A1 => n30574, A2 => n39312, B1 => n30638, B2 =>
                           n39306, C1 => n30510, C2 => n39300, ZN => n35404);
   U34259 : AOI221_X1 port map( B1 => n39444, B2 => n29072, C1 => n39438, C2 =>
                           n29136, A => n35396, ZN => n35389);
   U34260 : OAI222_X1 port map( A1 => n31460, A2 => n39432, B1 => n31524, B2 =>
                           n39426, C1 => n31396, C2 => n39420, ZN => n35396);
   U34261 : AOI221_X1 port map( B1 => n39576, B2 => n32534, C1 => n39570, C2 =>
                           n27972, A => n34149, ZN => n34142);
   U34262 : OAI222_X1 port map( A1 => n30573, A2 => n39564, B1 => n30637, B2 =>
                           n39558, C1 => n30509, C2 => n39552, ZN => n34149);
   U34263 : AOI221_X1 port map( B1 => n39696, B2 => n29071, C1 => n39690, C2 =>
                           n29135, A => n34141, ZN => n34134);
   U34264 : OAI222_X1 port map( A1 => n31459, A2 => n39684, B1 => n31523, B2 =>
                           n39678, C1 => n31395, C2 => n39672, ZN => n34141);
   U34265 : AOI221_X1 port map( B1 => n39324, B2 => n32534, C1 => n39318, C2 =>
                           n27972, A => n35423, ZN => n35416);
   U34266 : OAI222_X1 port map( A1 => n30573, A2 => n39312, B1 => n30637, B2 =>
                           n39306, C1 => n30509, C2 => n39300, ZN => n35423);
   U34267 : AOI221_X1 port map( B1 => n39444, B2 => n29071, C1 => n39438, C2 =>
                           n29135, A => n35415, ZN => n35408);
   U34268 : OAI222_X1 port map( A1 => n31459, A2 => n39432, B1 => n31523, B2 =>
                           n39426, C1 => n31395, C2 => n39420, ZN => n35415);
   U34269 : AOI221_X1 port map( B1 => n39576, B2 => n32533, C1 => n39570, C2 =>
                           n27971, A => n34168, ZN => n34161);
   U34270 : OAI222_X1 port map( A1 => n30572, A2 => n39564, B1 => n30636, B2 =>
                           n39558, C1 => n30508, C2 => n39552, ZN => n34168);
   U34271 : AOI221_X1 port map( B1 => n39696, B2 => n29070, C1 => n39690, C2 =>
                           n29134, A => n34160, ZN => n34153);
   U34272 : OAI222_X1 port map( A1 => n31458, A2 => n39684, B1 => n31522, B2 =>
                           n39678, C1 => n31394, C2 => n39672, ZN => n34160);
   U34273 : AOI221_X1 port map( B1 => n39324, B2 => n32533, C1 => n39318, C2 =>
                           n27971, A => n35442, ZN => n35435);
   U34274 : OAI222_X1 port map( A1 => n30572, A2 => n39312, B1 => n30636, B2 =>
                           n39306, C1 => n30508, C2 => n39300, ZN => n35442);
   U34275 : AOI221_X1 port map( B1 => n39444, B2 => n29070, C1 => n39438, C2 =>
                           n29134, A => n35434, ZN => n35427);
   U34276 : OAI222_X1 port map( A1 => n31458, A2 => n39432, B1 => n31522, B2 =>
                           n39426, C1 => n31394, C2 => n39420, ZN => n35434);
   U34277 : AOI221_X1 port map( B1 => n39576, B2 => n32532, C1 => n39570, C2 =>
                           n27970, A => n34187, ZN => n34180);
   U34278 : OAI222_X1 port map( A1 => n30571, A2 => n39564, B1 => n30635, B2 =>
                           n39558, C1 => n30507, C2 => n39552, ZN => n34187);
   U34279 : AOI221_X1 port map( B1 => n39696, B2 => n29069, C1 => n39690, C2 =>
                           n29133, A => n34179, ZN => n34172);
   U34280 : OAI222_X1 port map( A1 => n31457, A2 => n39684, B1 => n31521, B2 =>
                           n39678, C1 => n31393, C2 => n39672, ZN => n34179);
   U34281 : AOI221_X1 port map( B1 => n39324, B2 => n32532, C1 => n39318, C2 =>
                           n27970, A => n35461, ZN => n35454);
   U34282 : OAI222_X1 port map( A1 => n30571, A2 => n39312, B1 => n30635, B2 =>
                           n39306, C1 => n30507, C2 => n39300, ZN => n35461);
   U34283 : AOI221_X1 port map( B1 => n39444, B2 => n29069, C1 => n39438, C2 =>
                           n29133, A => n35453, ZN => n35446);
   U34284 : OAI222_X1 port map( A1 => n31457, A2 => n39432, B1 => n31521, B2 =>
                           n39426, C1 => n31393, C2 => n39420, ZN => n35453);
   U34285 : AOI221_X1 port map( B1 => n39576, B2 => n32531, C1 => n39570, C2 =>
                           n27969, A => n34206, ZN => n34199);
   U34286 : OAI222_X1 port map( A1 => n30570, A2 => n39564, B1 => n30634, B2 =>
                           n39558, C1 => n30506, C2 => n39552, ZN => n34206);
   U34287 : AOI221_X1 port map( B1 => n39696, B2 => n29068, C1 => n39690, C2 =>
                           n29132, A => n34198, ZN => n34191);
   U34288 : OAI222_X1 port map( A1 => n31456, A2 => n39684, B1 => n31520, B2 =>
                           n39678, C1 => n31392, C2 => n39672, ZN => n34198);
   U34289 : AOI221_X1 port map( B1 => n39324, B2 => n32531, C1 => n39318, C2 =>
                           n27969, A => n35480, ZN => n35473);
   U34290 : OAI222_X1 port map( A1 => n30570, A2 => n39312, B1 => n30634, B2 =>
                           n39306, C1 => n30506, C2 => n39300, ZN => n35480);
   U34291 : AOI221_X1 port map( B1 => n39444, B2 => n29068, C1 => n39438, C2 =>
                           n29132, A => n35472, ZN => n35465);
   U34292 : OAI222_X1 port map( A1 => n31456, A2 => n39432, B1 => n31520, B2 =>
                           n39426, C1 => n31392, C2 => n39420, ZN => n35472);
   U34293 : AOI221_X1 port map( B1 => n39576, B2 => n32530, C1 => n39570, C2 =>
                           n27968, A => n34225, ZN => n34218);
   U34294 : OAI222_X1 port map( A1 => n30569, A2 => n39564, B1 => n30633, B2 =>
                           n39558, C1 => n30505, C2 => n39552, ZN => n34225);
   U34295 : AOI221_X1 port map( B1 => n39696, B2 => n29067, C1 => n39690, C2 =>
                           n29131, A => n34217, ZN => n34210);
   U34296 : OAI222_X1 port map( A1 => n31455, A2 => n39684, B1 => n31519, B2 =>
                           n39678, C1 => n31391, C2 => n39672, ZN => n34217);
   U34297 : AOI221_X1 port map( B1 => n39324, B2 => n32530, C1 => n39318, C2 =>
                           n27968, A => n35499, ZN => n35492);
   U34298 : OAI222_X1 port map( A1 => n30569, A2 => n39312, B1 => n30633, B2 =>
                           n39306, C1 => n30505, C2 => n39300, ZN => n35499);
   U34299 : AOI221_X1 port map( B1 => n39444, B2 => n29067, C1 => n39438, C2 =>
                           n29131, A => n35491, ZN => n35484);
   U34300 : OAI222_X1 port map( A1 => n31455, A2 => n39432, B1 => n31519, B2 =>
                           n39426, C1 => n31391, C2 => n39420, ZN => n35491);
   U34301 : AOI221_X1 port map( B1 => n39575, B2 => n32529, C1 => n39569, C2 =>
                           n27967, A => n34244, ZN => n34237);
   U34302 : OAI222_X1 port map( A1 => n30568, A2 => n39563, B1 => n30632, B2 =>
                           n39557, C1 => n30504, C2 => n39551, ZN => n34244);
   U34303 : AOI221_X1 port map( B1 => n39695, B2 => n29066, C1 => n39689, C2 =>
                           n29130, A => n34236, ZN => n34229);
   U34304 : OAI222_X1 port map( A1 => n31454, A2 => n39683, B1 => n31518, B2 =>
                           n39677, C1 => n31390, C2 => n39671, ZN => n34236);
   U34305 : AOI221_X1 port map( B1 => n39323, B2 => n32529, C1 => n39317, C2 =>
                           n27967, A => n35518, ZN => n35511);
   U34306 : OAI222_X1 port map( A1 => n30568, A2 => n39311, B1 => n30632, B2 =>
                           n39305, C1 => n30504, C2 => n39299, ZN => n35518);
   U34307 : AOI221_X1 port map( B1 => n39443, B2 => n29066, C1 => n39437, C2 =>
                           n29130, A => n35510, ZN => n35503);
   U34308 : OAI222_X1 port map( A1 => n31454, A2 => n39431, B1 => n31518, B2 =>
                           n39425, C1 => n31390, C2 => n39419, ZN => n35510);
   U34309 : AOI221_X1 port map( B1 => n39575, B2 => n32528, C1 => n39569, C2 =>
                           n27966, A => n34263, ZN => n34256);
   U34310 : OAI222_X1 port map( A1 => n30567, A2 => n39563, B1 => n30631, B2 =>
                           n39557, C1 => n30503, C2 => n39551, ZN => n34263);
   U34311 : AOI221_X1 port map( B1 => n39695, B2 => n29065, C1 => n39689, C2 =>
                           n29129, A => n34255, ZN => n34248);
   U34312 : OAI222_X1 port map( A1 => n31453, A2 => n39683, B1 => n31517, B2 =>
                           n39677, C1 => n31389, C2 => n39671, ZN => n34255);
   U34313 : AOI221_X1 port map( B1 => n39323, B2 => n32528, C1 => n39317, C2 =>
                           n27966, A => n35537, ZN => n35530);
   U34314 : OAI222_X1 port map( A1 => n30567, A2 => n39311, B1 => n30631, B2 =>
                           n39305, C1 => n30503, C2 => n39299, ZN => n35537);
   U34315 : AOI221_X1 port map( B1 => n39443, B2 => n29065, C1 => n39437, C2 =>
                           n29129, A => n35529, ZN => n35522);
   U34316 : OAI222_X1 port map( A1 => n31453, A2 => n39431, B1 => n31517, B2 =>
                           n39425, C1 => n31389, C2 => n39419, ZN => n35529);
   U34317 : AOI221_X1 port map( B1 => n39575, B2 => n32527, C1 => n39569, C2 =>
                           n27965, A => n34282, ZN => n34275);
   U34318 : OAI222_X1 port map( A1 => n30566, A2 => n39563, B1 => n30630, B2 =>
                           n39557, C1 => n30502, C2 => n39551, ZN => n34282);
   U34319 : AOI221_X1 port map( B1 => n39695, B2 => n29064, C1 => n39689, C2 =>
                           n29128, A => n34274, ZN => n34267);
   U34320 : OAI222_X1 port map( A1 => n31452, A2 => n39683, B1 => n31516, B2 =>
                           n39677, C1 => n31388, C2 => n39671, ZN => n34274);
   U34321 : AOI221_X1 port map( B1 => n39323, B2 => n32527, C1 => n39317, C2 =>
                           n27965, A => n35556, ZN => n35549);
   U34322 : OAI222_X1 port map( A1 => n30566, A2 => n39311, B1 => n30630, B2 =>
                           n39305, C1 => n30502, C2 => n39299, ZN => n35556);
   U34323 : AOI221_X1 port map( B1 => n39443, B2 => n29064, C1 => n39437, C2 =>
                           n29128, A => n35548, ZN => n35541);
   U34324 : OAI222_X1 port map( A1 => n31452, A2 => n39431, B1 => n31516, B2 =>
                           n39425, C1 => n31388, C2 => n39419, ZN => n35548);
   U34325 : AOI221_X1 port map( B1 => n39575, B2 => n32526, C1 => n39569, C2 =>
                           n27964, A => n34301, ZN => n34294);
   U34326 : OAI222_X1 port map( A1 => n30565, A2 => n39563, B1 => n30629, B2 =>
                           n39557, C1 => n30501, C2 => n39551, ZN => n34301);
   U34327 : AOI221_X1 port map( B1 => n39695, B2 => n29063, C1 => n39689, C2 =>
                           n29127, A => n34293, ZN => n34286);
   U34328 : OAI222_X1 port map( A1 => n31451, A2 => n39683, B1 => n31515, B2 =>
                           n39677, C1 => n31387, C2 => n39671, ZN => n34293);
   U34329 : AOI221_X1 port map( B1 => n39323, B2 => n32526, C1 => n39317, C2 =>
                           n27964, A => n35575, ZN => n35568);
   U34330 : OAI222_X1 port map( A1 => n30565, A2 => n39311, B1 => n30629, B2 =>
                           n39305, C1 => n30501, C2 => n39299, ZN => n35575);
   U34331 : AOI221_X1 port map( B1 => n39443, B2 => n29063, C1 => n39437, C2 =>
                           n29127, A => n35567, ZN => n35560);
   U34332 : OAI222_X1 port map( A1 => n31451, A2 => n39431, B1 => n31515, B2 =>
                           n39425, C1 => n31387, C2 => n39419, ZN => n35567);
   U34333 : AOI221_X1 port map( B1 => n39575, B2 => n32525, C1 => n39569, C2 =>
                           n27963, A => n34320, ZN => n34313);
   U34334 : OAI222_X1 port map( A1 => n30564, A2 => n39563, B1 => n30628, B2 =>
                           n39557, C1 => n30500, C2 => n39551, ZN => n34320);
   U34335 : AOI221_X1 port map( B1 => n39695, B2 => n29062, C1 => n39689, C2 =>
                           n29126, A => n34312, ZN => n34305);
   U34336 : OAI222_X1 port map( A1 => n31450, A2 => n39683, B1 => n31514, B2 =>
                           n39677, C1 => n31386, C2 => n39671, ZN => n34312);
   U34337 : AOI221_X1 port map( B1 => n39323, B2 => n32525, C1 => n39317, C2 =>
                           n27963, A => n35594, ZN => n35587);
   U34338 : OAI222_X1 port map( A1 => n30564, A2 => n39311, B1 => n30628, B2 =>
                           n39305, C1 => n30500, C2 => n39299, ZN => n35594);
   U34339 : AOI221_X1 port map( B1 => n39443, B2 => n29062, C1 => n39437, C2 =>
                           n29126, A => n35586, ZN => n35579);
   U34340 : OAI222_X1 port map( A1 => n31450, A2 => n39431, B1 => n31514, B2 =>
                           n39425, C1 => n31386, C2 => n39419, ZN => n35586);
   U34341 : AOI221_X1 port map( B1 => n39575, B2 => n32524, C1 => n39569, C2 =>
                           n27962, A => n34339, ZN => n34332);
   U34342 : OAI222_X1 port map( A1 => n30563, A2 => n39563, B1 => n30627, B2 =>
                           n39557, C1 => n30499, C2 => n39551, ZN => n34339);
   U34343 : AOI221_X1 port map( B1 => n39695, B2 => n29061, C1 => n39689, C2 =>
                           n29125, A => n34331, ZN => n34324);
   U34344 : OAI222_X1 port map( A1 => n31449, A2 => n39683, B1 => n31513, B2 =>
                           n39677, C1 => n31385, C2 => n39671, ZN => n34331);
   U34345 : AOI221_X1 port map( B1 => n39323, B2 => n32524, C1 => n39317, C2 =>
                           n27962, A => n35613, ZN => n35606);
   U34346 : OAI222_X1 port map( A1 => n30563, A2 => n39311, B1 => n30627, B2 =>
                           n39305, C1 => n30499, C2 => n39299, ZN => n35613);
   U34347 : AOI221_X1 port map( B1 => n39443, B2 => n29061, C1 => n39437, C2 =>
                           n29125, A => n35605, ZN => n35598);
   U34348 : OAI222_X1 port map( A1 => n31449, A2 => n39431, B1 => n31513, B2 =>
                           n39425, C1 => n31385, C2 => n39419, ZN => n35605);
   U34349 : AOI221_X1 port map( B1 => n39575, B2 => n32523, C1 => n39569, C2 =>
                           n27961, A => n34358, ZN => n34351);
   U34350 : OAI222_X1 port map( A1 => n30562, A2 => n39563, B1 => n30626, B2 =>
                           n39557, C1 => n30498, C2 => n39551, ZN => n34358);
   U34351 : AOI221_X1 port map( B1 => n39695, B2 => n29060, C1 => n39689, C2 =>
                           n29124, A => n34350, ZN => n34343);
   U34352 : OAI222_X1 port map( A1 => n31448, A2 => n39683, B1 => n31512, B2 =>
                           n39677, C1 => n31384, C2 => n39671, ZN => n34350);
   U34353 : AOI221_X1 port map( B1 => n39323, B2 => n32523, C1 => n39317, C2 =>
                           n27961, A => n35632, ZN => n35625);
   U34354 : OAI222_X1 port map( A1 => n30562, A2 => n39311, B1 => n30626, B2 =>
                           n39305, C1 => n30498, C2 => n39299, ZN => n35632);
   U34355 : AOI221_X1 port map( B1 => n39443, B2 => n29060, C1 => n39437, C2 =>
                           n29124, A => n35624, ZN => n35617);
   U34356 : OAI222_X1 port map( A1 => n31448, A2 => n39431, B1 => n31512, B2 =>
                           n39425, C1 => n31384, C2 => n39419, ZN => n35624);
   U34357 : AOI221_X1 port map( B1 => n39575, B2 => n32522, C1 => n39569, C2 =>
                           n27960, A => n34377, ZN => n34370);
   U34358 : OAI222_X1 port map( A1 => n30561, A2 => n39563, B1 => n30625, B2 =>
                           n39557, C1 => n30497, C2 => n39551, ZN => n34377);
   U34359 : AOI221_X1 port map( B1 => n39695, B2 => n29059, C1 => n39689, C2 =>
                           n29123, A => n34369, ZN => n34362);
   U34360 : OAI222_X1 port map( A1 => n31447, A2 => n39683, B1 => n31511, B2 =>
                           n39677, C1 => n31383, C2 => n39671, ZN => n34369);
   U34361 : AOI221_X1 port map( B1 => n39323, B2 => n32522, C1 => n39317, C2 =>
                           n27960, A => n35651, ZN => n35644);
   U34362 : OAI222_X1 port map( A1 => n30561, A2 => n39311, B1 => n30625, B2 =>
                           n39305, C1 => n30497, C2 => n39299, ZN => n35651);
   U34363 : AOI221_X1 port map( B1 => n39443, B2 => n29059, C1 => n39437, C2 =>
                           n29123, A => n35643, ZN => n35636);
   U34364 : OAI222_X1 port map( A1 => n31447, A2 => n39431, B1 => n31511, B2 =>
                           n39425, C1 => n31383, C2 => n39419, ZN => n35643);
   U34365 : AOI221_X1 port map( B1 => n39575, B2 => n32521, C1 => n39569, C2 =>
                           n27959, A => n34396, ZN => n34389);
   U34366 : OAI222_X1 port map( A1 => n30560, A2 => n39563, B1 => n30624, B2 =>
                           n39557, C1 => n30496, C2 => n39551, ZN => n34396);
   U34367 : AOI221_X1 port map( B1 => n39695, B2 => n29058, C1 => n39689, C2 =>
                           n29122, A => n34388, ZN => n34381);
   U34368 : OAI222_X1 port map( A1 => n31446, A2 => n39683, B1 => n31510, B2 =>
                           n39677, C1 => n31382, C2 => n39671, ZN => n34388);
   U34369 : AOI221_X1 port map( B1 => n39323, B2 => n32521, C1 => n39317, C2 =>
                           n27959, A => n35670, ZN => n35663);
   U34370 : OAI222_X1 port map( A1 => n30560, A2 => n39311, B1 => n30624, B2 =>
                           n39305, C1 => n30496, C2 => n39299, ZN => n35670);
   U34371 : AOI221_X1 port map( B1 => n39443, B2 => n29058, C1 => n39437, C2 =>
                           n29122, A => n35662, ZN => n35655);
   U34372 : OAI222_X1 port map( A1 => n31446, A2 => n39431, B1 => n31510, B2 =>
                           n39425, C1 => n31382, C2 => n39419, ZN => n35662);
   U34373 : AOI221_X1 port map( B1 => n39575, B2 => n32520, C1 => n39569, C2 =>
                           n27958, A => n34415, ZN => n34408);
   U34374 : OAI222_X1 port map( A1 => n30559, A2 => n39563, B1 => n30623, B2 =>
                           n39557, C1 => n30495, C2 => n39551, ZN => n34415);
   U34375 : AOI221_X1 port map( B1 => n39695, B2 => n29057, C1 => n39689, C2 =>
                           n29121, A => n34407, ZN => n34400);
   U34376 : OAI222_X1 port map( A1 => n31445, A2 => n39683, B1 => n31509, B2 =>
                           n39677, C1 => n31381, C2 => n39671, ZN => n34407);
   U34377 : AOI221_X1 port map( B1 => n39323, B2 => n32520, C1 => n39317, C2 =>
                           n27958, A => n35689, ZN => n35682);
   U34378 : OAI222_X1 port map( A1 => n30559, A2 => n39311, B1 => n30623, B2 =>
                           n39305, C1 => n30495, C2 => n39299, ZN => n35689);
   U34379 : AOI221_X1 port map( B1 => n39443, B2 => n29057, C1 => n39437, C2 =>
                           n29121, A => n35681, ZN => n35674);
   U34380 : OAI222_X1 port map( A1 => n31445, A2 => n39431, B1 => n31509, B2 =>
                           n39425, C1 => n31381, C2 => n39419, ZN => n35681);
   U34381 : AOI221_X1 port map( B1 => n39575, B2 => n32519, C1 => n39569, C2 =>
                           n27957, A => n34434, ZN => n34427);
   U34382 : OAI222_X1 port map( A1 => n30558, A2 => n39563, B1 => n30622, B2 =>
                           n39557, C1 => n30494, C2 => n39551, ZN => n34434);
   U34383 : AOI221_X1 port map( B1 => n39695, B2 => n29056, C1 => n39689, C2 =>
                           n29120, A => n34426, ZN => n34419);
   U34384 : OAI222_X1 port map( A1 => n31444, A2 => n39683, B1 => n31508, B2 =>
                           n39677, C1 => n31380, C2 => n39671, ZN => n34426);
   U34385 : AOI221_X1 port map( B1 => n39323, B2 => n32519, C1 => n39317, C2 =>
                           n27957, A => n35708, ZN => n35701);
   U34386 : OAI222_X1 port map( A1 => n30558, A2 => n39311, B1 => n30622, B2 =>
                           n39305, C1 => n30494, C2 => n39299, ZN => n35708);
   U34387 : AOI221_X1 port map( B1 => n39443, B2 => n29056, C1 => n39437, C2 =>
                           n29120, A => n35700, ZN => n35693);
   U34388 : OAI222_X1 port map( A1 => n31444, A2 => n39431, B1 => n31508, B2 =>
                           n39425, C1 => n31380, C2 => n39419, ZN => n35700);
   U34389 : AOI221_X1 port map( B1 => n39575, B2 => n32518, C1 => n39569, C2 =>
                           n27956, A => n34453, ZN => n34446);
   U34390 : OAI222_X1 port map( A1 => n30557, A2 => n39563, B1 => n30621, B2 =>
                           n39557, C1 => n30493, C2 => n39551, ZN => n34453);
   U34391 : AOI221_X1 port map( B1 => n39695, B2 => n29055, C1 => n39689, C2 =>
                           n29119, A => n34445, ZN => n34438);
   U34392 : OAI222_X1 port map( A1 => n31443, A2 => n39683, B1 => n31507, B2 =>
                           n39677, C1 => n31379, C2 => n39671, ZN => n34445);
   U34393 : AOI221_X1 port map( B1 => n39323, B2 => n32518, C1 => n39317, C2 =>
                           n27956, A => n35727, ZN => n35720);
   U34394 : OAI222_X1 port map( A1 => n30557, A2 => n39311, B1 => n30621, B2 =>
                           n39305, C1 => n30493, C2 => n39299, ZN => n35727);
   U34395 : AOI221_X1 port map( B1 => n39443, B2 => n29055, C1 => n39437, C2 =>
                           n29119, A => n35719, ZN => n35712);
   U34396 : OAI222_X1 port map( A1 => n31443, A2 => n39431, B1 => n31507, B2 =>
                           n39425, C1 => n31379, C2 => n39419, ZN => n35719);
   U34397 : AOI221_X1 port map( B1 => n39574, B2 => n32517, C1 => n39568, C2 =>
                           n27955, A => n34472, ZN => n34465);
   U34398 : OAI222_X1 port map( A1 => n30556, A2 => n39562, B1 => n30620, B2 =>
                           n39556, C1 => n30492, C2 => n39550, ZN => n34472);
   U34399 : AOI221_X1 port map( B1 => n39694, B2 => n29054, C1 => n39688, C2 =>
                           n29118, A => n34464, ZN => n34457);
   U34400 : OAI222_X1 port map( A1 => n31442, A2 => n39682, B1 => n31506, B2 =>
                           n39676, C1 => n31378, C2 => n39670, ZN => n34464);
   U34401 : AOI221_X1 port map( B1 => n39322, B2 => n32517, C1 => n39316, C2 =>
                           n27955, A => n35746, ZN => n35739);
   U34402 : OAI222_X1 port map( A1 => n30556, A2 => n39310, B1 => n30620, B2 =>
                           n39304, C1 => n30492, C2 => n39298, ZN => n35746);
   U34403 : AOI221_X1 port map( B1 => n39442, B2 => n29054, C1 => n39436, C2 =>
                           n29118, A => n35738, ZN => n35731);
   U34404 : OAI222_X1 port map( A1 => n31442, A2 => n39430, B1 => n31506, B2 =>
                           n39424, C1 => n31378, C2 => n39418, ZN => n35738);
   U34405 : AOI221_X1 port map( B1 => n39574, B2 => n32516, C1 => n39568, C2 =>
                           n27954, A => n34491, ZN => n34484);
   U34406 : OAI222_X1 port map( A1 => n30555, A2 => n39562, B1 => n30619, B2 =>
                           n39556, C1 => n30491, C2 => n39550, ZN => n34491);
   U34407 : AOI221_X1 port map( B1 => n39694, B2 => n29053, C1 => n39688, C2 =>
                           n29117, A => n34483, ZN => n34476);
   U34408 : OAI222_X1 port map( A1 => n31441, A2 => n39682, B1 => n31505, B2 =>
                           n39676, C1 => n31377, C2 => n39670, ZN => n34483);
   U34409 : AOI221_X1 port map( B1 => n39322, B2 => n32516, C1 => n39316, C2 =>
                           n27954, A => n35765, ZN => n35758);
   U34410 : OAI222_X1 port map( A1 => n30555, A2 => n39310, B1 => n30619, B2 =>
                           n39304, C1 => n30491, C2 => n39298, ZN => n35765);
   U34411 : AOI221_X1 port map( B1 => n39442, B2 => n29053, C1 => n39436, C2 =>
                           n29117, A => n35757, ZN => n35750);
   U34412 : OAI222_X1 port map( A1 => n31441, A2 => n39430, B1 => n31505, B2 =>
                           n39424, C1 => n31377, C2 => n39418, ZN => n35757);
   U34413 : AOI221_X1 port map( B1 => n39574, B2 => n32515, C1 => n39568, C2 =>
                           n27953, A => n34510, ZN => n34503);
   U34414 : OAI222_X1 port map( A1 => n30554, A2 => n39562, B1 => n30618, B2 =>
                           n39556, C1 => n30490, C2 => n39550, ZN => n34510);
   U34415 : AOI221_X1 port map( B1 => n39694, B2 => n29052, C1 => n39688, C2 =>
                           n29116, A => n34502, ZN => n34495);
   U34416 : OAI222_X1 port map( A1 => n31440, A2 => n39682, B1 => n31504, B2 =>
                           n39676, C1 => n31376, C2 => n39670, ZN => n34502);
   U34417 : AOI221_X1 port map( B1 => n39322, B2 => n32515, C1 => n39316, C2 =>
                           n27953, A => n35784, ZN => n35777);
   U34418 : OAI222_X1 port map( A1 => n30554, A2 => n39310, B1 => n30618, B2 =>
                           n39304, C1 => n30490, C2 => n39298, ZN => n35784);
   U34419 : AOI221_X1 port map( B1 => n39442, B2 => n29052, C1 => n39436, C2 =>
                           n29116, A => n35776, ZN => n35769);
   U34420 : OAI222_X1 port map( A1 => n31440, A2 => n39430, B1 => n31504, B2 =>
                           n39424, C1 => n31376, C2 => n39418, ZN => n35776);
   U34421 : AOI221_X1 port map( B1 => n39574, B2 => n32514, C1 => n39568, C2 =>
                           n27952, A => n34529, ZN => n34522);
   U34422 : OAI222_X1 port map( A1 => n30553, A2 => n39562, B1 => n30617, B2 =>
                           n39556, C1 => n30489, C2 => n39550, ZN => n34529);
   U34423 : AOI221_X1 port map( B1 => n39694, B2 => n29051, C1 => n39688, C2 =>
                           n29115, A => n34521, ZN => n34514);
   U34424 : OAI222_X1 port map( A1 => n31439, A2 => n39682, B1 => n31503, B2 =>
                           n39676, C1 => n31375, C2 => n39670, ZN => n34521);
   U34425 : AOI221_X1 port map( B1 => n39322, B2 => n32514, C1 => n39316, C2 =>
                           n27952, A => n35803, ZN => n35796);
   U34426 : OAI222_X1 port map( A1 => n30553, A2 => n39310, B1 => n30617, B2 =>
                           n39304, C1 => n30489, C2 => n39298, ZN => n35803);
   U34427 : AOI221_X1 port map( B1 => n39442, B2 => n29051, C1 => n39436, C2 =>
                           n29115, A => n35795, ZN => n35788);
   U34428 : OAI222_X1 port map( A1 => n31439, A2 => n39430, B1 => n31503, B2 =>
                           n39424, C1 => n31375, C2 => n39418, ZN => n35795);
   U34429 : AOI221_X1 port map( B1 => n39574, B2 => n32513, C1 => n39568, C2 =>
                           n27951, A => n34548, ZN => n34541);
   U34430 : OAI222_X1 port map( A1 => n30552, A2 => n39562, B1 => n30616, B2 =>
                           n39556, C1 => n30488, C2 => n39550, ZN => n34548);
   U34431 : AOI221_X1 port map( B1 => n39694, B2 => n29050, C1 => n39688, C2 =>
                           n29114, A => n34540, ZN => n34533);
   U34432 : OAI222_X1 port map( A1 => n31438, A2 => n39682, B1 => n31502, B2 =>
                           n39676, C1 => n31374, C2 => n39670, ZN => n34540);
   U34433 : AOI221_X1 port map( B1 => n39322, B2 => n32513, C1 => n39316, C2 =>
                           n27951, A => n35822, ZN => n35815);
   U34434 : OAI222_X1 port map( A1 => n30552, A2 => n39310, B1 => n30616, B2 =>
                           n39304, C1 => n30488, C2 => n39298, ZN => n35822);
   U34435 : AOI221_X1 port map( B1 => n39442, B2 => n29050, C1 => n39436, C2 =>
                           n29114, A => n35814, ZN => n35807);
   U34436 : OAI222_X1 port map( A1 => n31438, A2 => n39430, B1 => n31502, B2 =>
                           n39424, C1 => n31374, C2 => n39418, ZN => n35814);
   U34437 : AOI221_X1 port map( B1 => n39574, B2 => n32512, C1 => n39568, C2 =>
                           n27950, A => n34567, ZN => n34560);
   U34438 : OAI222_X1 port map( A1 => n30551, A2 => n39562, B1 => n30615, B2 =>
                           n39556, C1 => n30487, C2 => n39550, ZN => n34567);
   U34439 : AOI221_X1 port map( B1 => n39694, B2 => n29049, C1 => n39688, C2 =>
                           n29113, A => n34559, ZN => n34552);
   U34440 : OAI222_X1 port map( A1 => n31437, A2 => n39682, B1 => n31501, B2 =>
                           n39676, C1 => n31373, C2 => n39670, ZN => n34559);
   U34441 : AOI221_X1 port map( B1 => n39322, B2 => n32512, C1 => n39316, C2 =>
                           n27950, A => n35841, ZN => n35834);
   U34442 : OAI222_X1 port map( A1 => n30551, A2 => n39310, B1 => n30615, B2 =>
                           n39304, C1 => n30487, C2 => n39298, ZN => n35841);
   U34443 : AOI221_X1 port map( B1 => n39442, B2 => n29049, C1 => n39436, C2 =>
                           n29113, A => n35833, ZN => n35826);
   U34444 : OAI222_X1 port map( A1 => n31437, A2 => n39430, B1 => n31501, B2 =>
                           n39424, C1 => n31373, C2 => n39418, ZN => n35833);
   U34445 : AOI221_X1 port map( B1 => n39574, B2 => n32511, C1 => n39568, C2 =>
                           n27949, A => n34586, ZN => n34579);
   U34446 : OAI222_X1 port map( A1 => n30550, A2 => n39562, B1 => n30614, B2 =>
                           n39556, C1 => n30486, C2 => n39550, ZN => n34586);
   U34447 : AOI221_X1 port map( B1 => n39694, B2 => n29048, C1 => n39688, C2 =>
                           n29112, A => n34578, ZN => n34571);
   U34448 : OAI222_X1 port map( A1 => n31436, A2 => n39682, B1 => n31500, B2 =>
                           n39676, C1 => n31372, C2 => n39670, ZN => n34578);
   U34449 : AOI221_X1 port map( B1 => n39322, B2 => n32511, C1 => n39316, C2 =>
                           n27949, A => n35860, ZN => n35853);
   U34450 : OAI222_X1 port map( A1 => n30550, A2 => n39310, B1 => n30614, B2 =>
                           n39304, C1 => n30486, C2 => n39298, ZN => n35860);
   U34451 : AOI221_X1 port map( B1 => n39442, B2 => n29048, C1 => n39436, C2 =>
                           n29112, A => n35852, ZN => n35845);
   U34452 : OAI222_X1 port map( A1 => n31436, A2 => n39430, B1 => n31500, B2 =>
                           n39424, C1 => n31372, C2 => n39418, ZN => n35852);
   U34453 : AOI221_X1 port map( B1 => n39574, B2 => n32510, C1 => n39568, C2 =>
                           n27948, A => n34605, ZN => n34598);
   U34454 : OAI222_X1 port map( A1 => n30549, A2 => n39562, B1 => n30613, B2 =>
                           n39556, C1 => n30485, C2 => n39550, ZN => n34605);
   U34455 : AOI221_X1 port map( B1 => n39694, B2 => n29047, C1 => n39688, C2 =>
                           n29111, A => n34597, ZN => n34590);
   U34456 : OAI222_X1 port map( A1 => n31435, A2 => n39682, B1 => n31499, B2 =>
                           n39676, C1 => n31371, C2 => n39670, ZN => n34597);
   U34457 : AOI221_X1 port map( B1 => n39322, B2 => n32510, C1 => n39316, C2 =>
                           n27948, A => n35879, ZN => n35872);
   U34458 : OAI222_X1 port map( A1 => n30549, A2 => n39310, B1 => n30613, B2 =>
                           n39304, C1 => n30485, C2 => n39298, ZN => n35879);
   U34459 : AOI221_X1 port map( B1 => n39442, B2 => n29047, C1 => n39436, C2 =>
                           n29111, A => n35871, ZN => n35864);
   U34460 : OAI222_X1 port map( A1 => n31435, A2 => n39430, B1 => n31499, B2 =>
                           n39424, C1 => n31371, C2 => n39418, ZN => n35871);
   U34461 : AOI221_X1 port map( B1 => n39574, B2 => n32507, C1 => n39568, C2 =>
                           n27947, A => n34624, ZN => n34617);
   U34462 : OAI222_X1 port map( A1 => n30548, A2 => n39562, B1 => n30612, B2 =>
                           n39556, C1 => n30484, C2 => n39550, ZN => n34624);
   U34463 : AOI221_X1 port map( B1 => n39694, B2 => n29046, C1 => n39688, C2 =>
                           n29110, A => n34616, ZN => n34609);
   U34464 : OAI222_X1 port map( A1 => n31434, A2 => n39682, B1 => n31498, B2 =>
                           n39676, C1 => n31370, C2 => n39670, ZN => n34616);
   U34465 : AOI221_X1 port map( B1 => n39322, B2 => n32507, C1 => n39316, C2 =>
                           n27947, A => n35898, ZN => n35891);
   U34466 : OAI222_X1 port map( A1 => n30548, A2 => n39310, B1 => n30612, B2 =>
                           n39304, C1 => n30484, C2 => n39298, ZN => n35898);
   U34467 : AOI221_X1 port map( B1 => n39442, B2 => n29046, C1 => n39436, C2 =>
                           n29110, A => n35890, ZN => n35883);
   U34468 : OAI222_X1 port map( A1 => n31434, A2 => n39430, B1 => n31498, B2 =>
                           n39424, C1 => n31370, C2 => n39418, ZN => n35890);
   U34469 : AOI221_X1 port map( B1 => n39574, B2 => n32506, C1 => n39568, C2 =>
                           n27946, A => n34643, ZN => n34636);
   U34470 : OAI222_X1 port map( A1 => n30547, A2 => n39562, B1 => n30611, B2 =>
                           n39556, C1 => n30483, C2 => n39550, ZN => n34643);
   U34471 : AOI221_X1 port map( B1 => n39694, B2 => n29045, C1 => n39688, C2 =>
                           n29109, A => n34635, ZN => n34628);
   U34472 : OAI222_X1 port map( A1 => n31433, A2 => n39682, B1 => n31497, B2 =>
                           n39676, C1 => n31369, C2 => n39670, ZN => n34635);
   U34473 : AOI221_X1 port map( B1 => n39322, B2 => n32506, C1 => n39316, C2 =>
                           n27946, A => n35917, ZN => n35910);
   U34474 : OAI222_X1 port map( A1 => n30547, A2 => n39310, B1 => n30611, B2 =>
                           n39304, C1 => n30483, C2 => n39298, ZN => n35917);
   U34475 : AOI221_X1 port map( B1 => n39442, B2 => n29045, C1 => n39436, C2 =>
                           n29109, A => n35909, ZN => n35902);
   U34476 : OAI222_X1 port map( A1 => n31433, A2 => n39430, B1 => n31497, B2 =>
                           n39424, C1 => n31369, C2 => n39418, ZN => n35909);
   U34477 : AOI221_X1 port map( B1 => n39574, B2 => n32509, C1 => n39568, C2 =>
                           n27945, A => n34662, ZN => n34655);
   U34478 : OAI222_X1 port map( A1 => n30546, A2 => n39562, B1 => n30610, B2 =>
                           n39556, C1 => n30482, C2 => n39550, ZN => n34662);
   U34479 : AOI221_X1 port map( B1 => n39694, B2 => n29044, C1 => n39688, C2 =>
                           n29108, A => n34654, ZN => n34647);
   U34480 : OAI222_X1 port map( A1 => n31432, A2 => n39682, B1 => n31496, B2 =>
                           n39676, C1 => n31368, C2 => n39670, ZN => n34654);
   U34481 : AOI221_X1 port map( B1 => n39322, B2 => n32509, C1 => n39316, C2 =>
                           n27945, A => n35936, ZN => n35929);
   U34482 : OAI222_X1 port map( A1 => n30546, A2 => n39310, B1 => n30610, B2 =>
                           n39304, C1 => n30482, C2 => n39298, ZN => n35936);
   U34483 : AOI221_X1 port map( B1 => n39442, B2 => n29044, C1 => n39436, C2 =>
                           n29108, A => n35928, ZN => n35921);
   U34484 : OAI222_X1 port map( A1 => n31432, A2 => n39430, B1 => n31496, B2 =>
                           n39424, C1 => n31368, C2 => n39418, ZN => n35928);
   U34485 : AOI221_X1 port map( B1 => n39574, B2 => n32508, C1 => n39568, C2 =>
                           n27944, A => n34695, ZN => n34685);
   U34486 : OAI222_X1 port map( A1 => n30545, A2 => n39562, B1 => n30609, B2 =>
                           n39556, C1 => n30481, C2 => n39550, ZN => n34695);
   U34487 : AOI221_X1 port map( B1 => n39694, B2 => n29043, C1 => n39688, C2 =>
                           n29107, A => n34683, ZN => n34666);
   U34488 : OAI222_X1 port map( A1 => n31431, A2 => n39682, B1 => n31495, B2 =>
                           n39676, C1 => n31367, C2 => n39670, ZN => n34683);
   U34489 : AOI221_X1 port map( B1 => n39322, B2 => n32508, C1 => n39316, C2 =>
                           n27944, A => n35969, ZN => n35959);
   U34490 : OAI222_X1 port map( A1 => n30545, A2 => n39310, B1 => n30609, B2 =>
                           n39304, C1 => n30481, C2 => n39298, ZN => n35969);
   U34491 : AOI221_X1 port map( B1 => n39442, B2 => n29043, C1 => n39436, C2 =>
                           n29107, A => n35957, ZN => n35940);
   U34492 : OAI222_X1 port map( A1 => n31431, A2 => n39430, B1 => n31495, B2 =>
                           n39424, C1 => n31367, C2 => n39418, ZN => n35957);
   U34493 : OAI22_X1 port map( A1 => n16938, A2 => n39295, B1 => n36078, B2 => 
                           n39293, ZN => n7198);
   U34494 : NOR2_X1 port map( A1 => n36079, A2 => n36080, ZN => n36078);
   U34495 : NAND4_X1 port map( A1 => n36081, A2 => n36082, A3 => n36083, A4 => 
                           n36084, ZN => n36080);
   U34496 : NAND4_X1 port map( A1 => n36089, A2 => n36090, A3 => n36091, A4 => 
                           n36092, ZN => n36079);
   U34497 : OAI22_X1 port map( A1 => n16939, A2 => n39294, B1 => n36059, B2 => 
                           n39293, ZN => n7199);
   U34498 : NOR2_X1 port map( A1 => n36060, A2 => n36061, ZN => n36059);
   U34499 : NAND4_X1 port map( A1 => n36062, A2 => n36063, A3 => n36064, A4 => 
                           n36065, ZN => n36061);
   U34500 : NAND4_X1 port map( A1 => n36070, A2 => n36071, A3 => n36072, A4 => 
                           n36073, ZN => n36060);
   U34501 : OAI22_X1 port map( A1 => n16940, A2 => n39296, B1 => n36040, B2 => 
                           n39293, ZN => n7200);
   U34502 : NOR2_X1 port map( A1 => n36041, A2 => n36042, ZN => n36040);
   U34503 : NAND4_X1 port map( A1 => n36043, A2 => n36044, A3 => n36045, A4 => 
                           n36046, ZN => n36042);
   U34504 : NAND4_X1 port map( A1 => n36051, A2 => n36052, A3 => n36053, A4 => 
                           n36054, ZN => n36041);
   U34505 : OAI22_X1 port map( A1 => n16941, A2 => n39295, B1 => n35980, B2 => 
                           n39293, ZN => n7201);
   U34506 : NOR2_X1 port map( A1 => n35982, A2 => n35983, ZN => n35980);
   U34507 : NAND4_X1 port map( A1 => n35984, A2 => n35985, A3 => n35986, A4 => 
                           n35987, ZN => n35983);
   U34508 : NAND4_X1 port map( A1 => n36012, A2 => n36013, A3 => n36014, A4 => 
                           n36015, ZN => n35982);
   U34509 : OAI22_X1 port map( A1 => n17069, A2 => n39801, B1 => n33425, B2 => 
                           n39795, ZN => n7330);
   U34510 : NOR2_X1 port map( A1 => n33427, A2 => n33428, ZN => n33425);
   U34511 : NAND4_X1 port map( A1 => n33429, A2 => n33430, A3 => n33431, A4 => 
                           n33432, ZN => n33428);
   U34512 : NAND4_X1 port map( A1 => n33457, A2 => n33458, A3 => n33459, A4 => 
                           n33460, ZN => n33427);
   U34513 : OAI22_X1 port map( A1 => n17005, A2 => n39549, B1 => n34699, B2 => 
                           n39543, ZN => n7266);
   U34514 : NOR2_X1 port map( A1 => n34701, A2 => n34702, ZN => n34699);
   U34515 : NAND4_X1 port map( A1 => n34703, A2 => n34704, A3 => n34705, A4 => 
                           n34706, ZN => n34702);
   U34516 : NAND4_X1 port map( A1 => n34731, A2 => n34732, A3 => n34733, A4 => 
                           n34734, ZN => n34701);
   U34517 : OAI22_X1 port map( A1 => n17068, A2 => n39801, B1 => n33485, B2 => 
                           n39795, ZN => n7329);
   U34518 : NOR2_X1 port map( A1 => n33486, A2 => n33487, ZN => n33485);
   U34519 : NAND4_X1 port map( A1 => n33488, A2 => n33489, A3 => n33490, A4 => 
                           n33491, ZN => n33487);
   U34520 : NAND4_X1 port map( A1 => n33496, A2 => n33497, A3 => n33498, A4 => 
                           n33499, ZN => n33486);
   U34521 : OAI22_X1 port map( A1 => n17004, A2 => n39549, B1 => n34759, B2 => 
                           n39543, ZN => n7265);
   U34522 : NOR2_X1 port map( A1 => n34760, A2 => n34761, ZN => n34759);
   U34523 : NAND4_X1 port map( A1 => n34762, A2 => n34763, A3 => n34764, A4 => 
                           n34765, ZN => n34761);
   U34524 : NAND4_X1 port map( A1 => n34770, A2 => n34771, A3 => n34772, A4 => 
                           n34773, ZN => n34760);
   U34525 : OAI22_X1 port map( A1 => n17067, A2 => n39801, B1 => n33504, B2 => 
                           n39795, ZN => n7328);
   U34526 : NOR2_X1 port map( A1 => n33505, A2 => n33506, ZN => n33504);
   U34527 : NAND4_X1 port map( A1 => n33507, A2 => n33508, A3 => n33509, A4 => 
                           n33510, ZN => n33506);
   U34528 : NAND4_X1 port map( A1 => n33515, A2 => n33516, A3 => n33517, A4 => 
                           n33518, ZN => n33505);
   U34529 : OAI22_X1 port map( A1 => n17003, A2 => n39549, B1 => n34778, B2 => 
                           n39543, ZN => n7264);
   U34530 : NOR2_X1 port map( A1 => n34779, A2 => n34780, ZN => n34778);
   U34531 : NAND4_X1 port map( A1 => n34781, A2 => n34782, A3 => n34783, A4 => 
                           n34784, ZN => n34780);
   U34532 : NAND4_X1 port map( A1 => n34789, A2 => n34790, A3 => n34791, A4 => 
                           n34792, ZN => n34779);
   U34533 : OAI22_X1 port map( A1 => n17066, A2 => n39801, B1 => n33523, B2 => 
                           n39795, ZN => n7327);
   U34534 : NOR2_X1 port map( A1 => n33524, A2 => n33525, ZN => n33523);
   U34535 : NAND4_X1 port map( A1 => n33526, A2 => n33527, A3 => n33528, A4 => 
                           n33529, ZN => n33525);
   U34536 : NAND4_X1 port map( A1 => n33534, A2 => n33535, A3 => n33536, A4 => 
                           n33537, ZN => n33524);
   U34537 : OAI22_X1 port map( A1 => n17002, A2 => n39549, B1 => n34797, B2 => 
                           n39543, ZN => n7263);
   U34538 : NOR2_X1 port map( A1 => n34798, A2 => n34799, ZN => n34797);
   U34539 : NAND4_X1 port map( A1 => n34800, A2 => n34801, A3 => n34802, A4 => 
                           n34803, ZN => n34799);
   U34540 : NAND4_X1 port map( A1 => n34808, A2 => n34809, A3 => n34810, A4 => 
                           n34811, ZN => n34798);
   U34541 : XOR2_X1 port map( A => n2683, B => n39047, Z => n33297);
   U34542 : NAND2_X1 port map( A1 => n32242, A2 => add_146_carry_4_port, ZN => 
                           n39047);
   U34543 : OAI22_X1 port map( A1 => n16878, A2 => n39296, B1 => n37218, B2 => 
                           n39288, ZN => n7138);
   U34544 : NOR2_X1 port map( A1 => n37219, A2 => n37220, ZN => n37218);
   U34545 : NAND4_X1 port map( A1 => n37221, A2 => n37222, A3 => n37223, A4 => 
                           n37224, ZN => n37220);
   U34546 : NAND4_X1 port map( A1 => n37241, A2 => n37242, A3 => n37243, A4 => 
                           n37244, ZN => n37219);
   U34547 : OAI22_X1 port map( A1 => n16932, A2 => n39295, B1 => n36192, B2 => 
                           n39292, ZN => n7192);
   U34548 : NOR2_X1 port map( A1 => n36193, A2 => n36194, ZN => n36192);
   U34549 : NAND4_X1 port map( A1 => n36195, A2 => n36196, A3 => n36197, A4 => 
                           n36198, ZN => n36194);
   U34550 : NAND4_X1 port map( A1 => n36203, A2 => n36204, A3 => n36205, A4 => 
                           n36206, ZN => n36193);
   U34551 : OAI22_X1 port map( A1 => n16933, A2 => n39294, B1 => n36173, B2 => 
                           n39292, ZN => n7193);
   U34552 : NOR2_X1 port map( A1 => n36174, A2 => n36175, ZN => n36173);
   U34553 : NAND4_X1 port map( A1 => n36176, A2 => n36177, A3 => n36178, A4 => 
                           n36179, ZN => n36175);
   U34554 : NAND4_X1 port map( A1 => n36184, A2 => n36185, A3 => n36186, A4 => 
                           n36187, ZN => n36174);
   U34555 : OAI22_X1 port map( A1 => n16934, A2 => n39296, B1 => n36154, B2 => 
                           n39292, ZN => n7194);
   U34556 : NOR2_X1 port map( A1 => n36155, A2 => n36156, ZN => n36154);
   U34557 : NAND4_X1 port map( A1 => n36157, A2 => n36158, A3 => n36159, A4 => 
                           n36160, ZN => n36156);
   U34558 : NAND4_X1 port map( A1 => n36165, A2 => n36166, A3 => n36167, A4 => 
                           n36168, ZN => n36155);
   U34559 : OAI22_X1 port map( A1 => n16935, A2 => n39295, B1 => n36135, B2 => 
                           n39292, ZN => n7195);
   U34560 : NOR2_X1 port map( A1 => n36136, A2 => n36137, ZN => n36135);
   U34561 : NAND4_X1 port map( A1 => n36138, A2 => n36139, A3 => n36140, A4 => 
                           n36141, ZN => n36137);
   U34562 : NAND4_X1 port map( A1 => n36146, A2 => n36147, A3 => n36148, A4 => 
                           n36149, ZN => n36136);
   U34563 : OAI22_X1 port map( A1 => n16936, A2 => n39294, B1 => n36116, B2 => 
                           n39292, ZN => n7196);
   U34564 : NOR2_X1 port map( A1 => n36117, A2 => n36118, ZN => n36116);
   U34565 : NAND4_X1 port map( A1 => n36119, A2 => n36120, A3 => n36121, A4 => 
                           n36122, ZN => n36118);
   U34566 : NAND4_X1 port map( A1 => n36127, A2 => n36128, A3 => n36129, A4 => 
                           n36130, ZN => n36117);
   U34567 : OAI22_X1 port map( A1 => n16937, A2 => n39296, B1 => n36097, B2 => 
                           n39292, ZN => n7197);
   U34568 : NOR2_X1 port map( A1 => n36098, A2 => n36099, ZN => n36097);
   U34569 : NAND4_X1 port map( A1 => n36100, A2 => n36101, A3 => n36102, A4 => 
                           n36103, ZN => n36099);
   U34570 : NAND4_X1 port map( A1 => n36108, A2 => n36109, A3 => n36110, A4 => 
                           n36111, ZN => n36098);
   U34571 : OAI22_X1 port map( A1 => n16889, A2 => n39296, B1 => n37009, B2 => 
                           n39288, ZN => n7149);
   U34572 : NOR2_X1 port map( A1 => n37010, A2 => n37011, ZN => n37009);
   U34573 : NAND4_X1 port map( A1 => n37012, A2 => n37013, A3 => n37014, A4 => 
                           n37015, ZN => n37011);
   U34574 : NAND4_X1 port map( A1 => n37020, A2 => n37021, A3 => n37022, A4 => 
                           n37023, ZN => n37010);
   U34575 : OAI22_X1 port map( A1 => n16890, A2 => n39296, B1 => n36990, B2 => 
                           n39289, ZN => n7150);
   U34576 : NOR2_X1 port map( A1 => n36991, A2 => n36992, ZN => n36990);
   U34577 : NAND4_X1 port map( A1 => n36993, A2 => n36994, A3 => n36995, A4 => 
                           n36996, ZN => n36992);
   U34578 : NAND4_X1 port map( A1 => n37001, A2 => n37002, A3 => n37003, A4 => 
                           n37004, ZN => n36991);
   U34579 : OAI22_X1 port map( A1 => n16891, A2 => n39296, B1 => n36971, B2 => 
                           n39289, ZN => n7151);
   U34580 : NOR2_X1 port map( A1 => n36972, A2 => n36973, ZN => n36971);
   U34581 : NAND4_X1 port map( A1 => n36974, A2 => n36975, A3 => n36976, A4 => 
                           n36977, ZN => n36973);
   U34582 : NAND4_X1 port map( A1 => n36982, A2 => n36983, A3 => n36984, A4 => 
                           n36985, ZN => n36972);
   U34583 : OAI22_X1 port map( A1 => n16892, A2 => n39296, B1 => n36952, B2 => 
                           n39289, ZN => n7152);
   U34584 : NOR2_X1 port map( A1 => n36953, A2 => n36954, ZN => n36952);
   U34585 : NAND4_X1 port map( A1 => n36955, A2 => n36956, A3 => n36957, A4 => 
                           n36958, ZN => n36954);
   U34586 : NAND4_X1 port map( A1 => n36963, A2 => n36964, A3 => n36965, A4 => 
                           n36966, ZN => n36953);
   U34587 : OAI22_X1 port map( A1 => n16893, A2 => n39296, B1 => n36933, B2 => 
                           n39289, ZN => n7153);
   U34588 : NOR2_X1 port map( A1 => n36934, A2 => n36935, ZN => n36933);
   U34589 : NAND4_X1 port map( A1 => n36936, A2 => n36937, A3 => n36938, A4 => 
                           n36939, ZN => n36935);
   U34590 : NAND4_X1 port map( A1 => n36944, A2 => n36945, A3 => n36946, A4 => 
                           n36947, ZN => n36934);
   U34591 : OAI22_X1 port map( A1 => n16894, A2 => n39296, B1 => n36914, B2 => 
                           n39289, ZN => n7154);
   U34592 : NOR2_X1 port map( A1 => n36915, A2 => n36916, ZN => n36914);
   U34593 : NAND4_X1 port map( A1 => n36917, A2 => n36918, A3 => n36919, A4 => 
                           n36920, ZN => n36916);
   U34594 : NAND4_X1 port map( A1 => n36925, A2 => n36926, A3 => n36927, A4 => 
                           n36928, ZN => n36915);
   U34595 : OAI22_X1 port map( A1 => n16895, A2 => n39296, B1 => n36895, B2 => 
                           n39289, ZN => n7155);
   U34596 : NOR2_X1 port map( A1 => n36896, A2 => n36897, ZN => n36895);
   U34597 : NAND4_X1 port map( A1 => n36898, A2 => n36899, A3 => n36900, A4 => 
                           n36901, ZN => n36897);
   U34598 : NAND4_X1 port map( A1 => n36906, A2 => n36907, A3 => n36908, A4 => 
                           n36909, ZN => n36896);
   U34599 : OAI22_X1 port map( A1 => n16896, A2 => n39296, B1 => n36876, B2 => 
                           n39289, ZN => n7156);
   U34600 : NOR2_X1 port map( A1 => n36877, A2 => n36878, ZN => n36876);
   U34601 : NAND4_X1 port map( A1 => n36879, A2 => n36880, A3 => n36881, A4 => 
                           n36882, ZN => n36878);
   U34602 : NAND4_X1 port map( A1 => n36887, A2 => n36888, A3 => n36889, A4 => 
                           n36890, ZN => n36877);
   U34603 : OAI22_X1 port map( A1 => n16897, A2 => n39295, B1 => n36857, B2 => 
                           n39289, ZN => n7157);
   U34604 : NOR2_X1 port map( A1 => n36858, A2 => n36859, ZN => n36857);
   U34605 : NAND4_X1 port map( A1 => n36860, A2 => n36861, A3 => n36862, A4 => 
                           n36863, ZN => n36859);
   U34606 : NAND4_X1 port map( A1 => n36868, A2 => n36869, A3 => n36870, A4 => 
                           n36871, ZN => n36858);
   U34607 : OAI22_X1 port map( A1 => n16898, A2 => n39296, B1 => n36838, B2 => 
                           n39289, ZN => n7158);
   U34608 : NOR2_X1 port map( A1 => n36839, A2 => n36840, ZN => n36838);
   U34609 : NAND4_X1 port map( A1 => n36841, A2 => n36842, A3 => n36843, A4 => 
                           n36844, ZN => n36840);
   U34610 : NAND4_X1 port map( A1 => n36849, A2 => n36850, A3 => n36851, A4 => 
                           n36852, ZN => n36839);
   U34611 : OAI22_X1 port map( A1 => n16899, A2 => n39295, B1 => n36819, B2 => 
                           n39289, ZN => n7159);
   U34612 : NOR2_X1 port map( A1 => n36820, A2 => n36821, ZN => n36819);
   U34613 : NAND4_X1 port map( A1 => n36822, A2 => n36823, A3 => n36824, A4 => 
                           n36825, ZN => n36821);
   U34614 : NAND4_X1 port map( A1 => n36830, A2 => n36831, A3 => n36832, A4 => 
                           n36833, ZN => n36820);
   U34615 : OAI22_X1 port map( A1 => n16900, A2 => n39296, B1 => n36800, B2 => 
                           n39289, ZN => n7160);
   U34616 : NOR2_X1 port map( A1 => n36801, A2 => n36802, ZN => n36800);
   U34617 : NAND4_X1 port map( A1 => n36803, A2 => n36804, A3 => n36805, A4 => 
                           n36806, ZN => n36802);
   U34618 : NAND4_X1 port map( A1 => n36811, A2 => n36812, A3 => n36813, A4 => 
                           n36814, ZN => n36801);
   U34619 : OAI22_X1 port map( A1 => n16901, A2 => n39295, B1 => n36781, B2 => 
                           n39289, ZN => n7161);
   U34620 : NOR2_X1 port map( A1 => n36782, A2 => n36783, ZN => n36781);
   U34621 : NAND4_X1 port map( A1 => n36784, A2 => n36785, A3 => n36786, A4 => 
                           n36787, ZN => n36783);
   U34622 : NAND4_X1 port map( A1 => n36792, A2 => n36793, A3 => n36794, A4 => 
                           n36795, ZN => n36782);
   U34623 : OAI22_X1 port map( A1 => n16902, A2 => n39296, B1 => n36762, B2 => 
                           n39290, ZN => n7162);
   U34624 : NOR2_X1 port map( A1 => n36763, A2 => n36764, ZN => n36762);
   U34625 : NAND4_X1 port map( A1 => n36765, A2 => n36766, A3 => n36767, A4 => 
                           n36768, ZN => n36764);
   U34626 : NAND4_X1 port map( A1 => n36773, A2 => n36774, A3 => n36775, A4 => 
                           n36776, ZN => n36763);
   U34627 : OAI22_X1 port map( A1 => n16903, A2 => n39295, B1 => n36743, B2 => 
                           n39290, ZN => n7163);
   U34628 : NOR2_X1 port map( A1 => n36744, A2 => n36745, ZN => n36743);
   U34629 : NAND4_X1 port map( A1 => n36746, A2 => n36747, A3 => n36748, A4 => 
                           n36749, ZN => n36745);
   U34630 : NAND4_X1 port map( A1 => n36754, A2 => n36755, A3 => n36756, A4 => 
                           n36757, ZN => n36744);
   U34631 : OAI22_X1 port map( A1 => n16904, A2 => n39296, B1 => n36724, B2 => 
                           n39290, ZN => n7164);
   U34632 : NOR2_X1 port map( A1 => n36725, A2 => n36726, ZN => n36724);
   U34633 : NAND4_X1 port map( A1 => n36727, A2 => n36728, A3 => n36729, A4 => 
                           n36730, ZN => n36726);
   U34634 : NAND4_X1 port map( A1 => n36735, A2 => n36736, A3 => n36737, A4 => 
                           n36738, ZN => n36725);
   U34635 : OAI22_X1 port map( A1 => n16905, A2 => n39295, B1 => n36705, B2 => 
                           n39290, ZN => n7165);
   U34636 : NOR2_X1 port map( A1 => n36706, A2 => n36707, ZN => n36705);
   U34637 : NAND4_X1 port map( A1 => n36708, A2 => n36709, A3 => n36710, A4 => 
                           n36711, ZN => n36707);
   U34638 : NAND4_X1 port map( A1 => n36716, A2 => n36717, A3 => n36718, A4 => 
                           n36719, ZN => n36706);
   U34639 : OAI22_X1 port map( A1 => n16906, A2 => n39296, B1 => n36686, B2 => 
                           n39290, ZN => n7166);
   U34640 : NOR2_X1 port map( A1 => n36687, A2 => n36688, ZN => n36686);
   U34641 : NAND4_X1 port map( A1 => n36689, A2 => n36690, A3 => n36691, A4 => 
                           n36692, ZN => n36688);
   U34642 : NAND4_X1 port map( A1 => n36697, A2 => n36698, A3 => n36699, A4 => 
                           n36700, ZN => n36687);
   U34643 : OAI22_X1 port map( A1 => n16907, A2 => n39295, B1 => n36667, B2 => 
                           n39290, ZN => n7167);
   U34644 : NOR2_X1 port map( A1 => n36668, A2 => n36669, ZN => n36667);
   U34645 : NAND4_X1 port map( A1 => n36670, A2 => n36671, A3 => n36672, A4 => 
                           n36673, ZN => n36669);
   U34646 : NAND4_X1 port map( A1 => n36678, A2 => n36679, A3 => n36680, A4 => 
                           n36681, ZN => n36668);
   U34647 : OAI22_X1 port map( A1 => n16908, A2 => n39295, B1 => n36648, B2 => 
                           n39290, ZN => n7168);
   U34648 : NOR2_X1 port map( A1 => n36649, A2 => n36650, ZN => n36648);
   U34649 : NAND4_X1 port map( A1 => n36651, A2 => n36652, A3 => n36653, A4 => 
                           n36654, ZN => n36650);
   U34650 : NAND4_X1 port map( A1 => n36659, A2 => n36660, A3 => n36661, A4 => 
                           n36662, ZN => n36649);
   U34651 : OAI22_X1 port map( A1 => n16909, A2 => n39295, B1 => n36629, B2 => 
                           n39290, ZN => n7169);
   U34652 : NOR2_X1 port map( A1 => n36630, A2 => n36631, ZN => n36629);
   U34653 : NAND4_X1 port map( A1 => n36632, A2 => n36633, A3 => n36634, A4 => 
                           n36635, ZN => n36631);
   U34654 : NAND4_X1 port map( A1 => n36640, A2 => n36641, A3 => n36642, A4 => 
                           n36643, ZN => n36630);
   U34655 : OAI22_X1 port map( A1 => n16910, A2 => n39295, B1 => n36610, B2 => 
                           n39290, ZN => n7170);
   U34656 : NOR2_X1 port map( A1 => n36611, A2 => n36612, ZN => n36610);
   U34657 : NAND4_X1 port map( A1 => n36613, A2 => n36614, A3 => n36615, A4 => 
                           n36616, ZN => n36612);
   U34658 : NAND4_X1 port map( A1 => n36621, A2 => n36622, A3 => n36623, A4 => 
                           n36624, ZN => n36611);
   U34659 : OAI22_X1 port map( A1 => n16911, A2 => n39295, B1 => n36591, B2 => 
                           n39290, ZN => n7171);
   U34660 : NOR2_X1 port map( A1 => n36592, A2 => n36593, ZN => n36591);
   U34661 : NAND4_X1 port map( A1 => n36594, A2 => n36595, A3 => n36596, A4 => 
                           n36597, ZN => n36593);
   U34662 : NAND4_X1 port map( A1 => n36602, A2 => n36603, A3 => n36604, A4 => 
                           n36605, ZN => n36592);
   U34663 : OAI22_X1 port map( A1 => n16912, A2 => n39295, B1 => n36572, B2 => 
                           n39290, ZN => n7172);
   U34664 : NOR2_X1 port map( A1 => n36573, A2 => n36574, ZN => n36572);
   U34665 : NAND4_X1 port map( A1 => n36575, A2 => n36576, A3 => n36577, A4 => 
                           n36578, ZN => n36574);
   U34666 : NAND4_X1 port map( A1 => n36583, A2 => n36584, A3 => n36585, A4 => 
                           n36586, ZN => n36573);
   U34667 : OAI22_X1 port map( A1 => n16913, A2 => n39295, B1 => n36553, B2 => 
                           n39290, ZN => n7173);
   U34668 : NOR2_X1 port map( A1 => n36554, A2 => n36555, ZN => n36553);
   U34669 : NAND4_X1 port map( A1 => n36556, A2 => n36557, A3 => n36558, A4 => 
                           n36559, ZN => n36555);
   U34670 : NAND4_X1 port map( A1 => n36564, A2 => n36565, A3 => n36566, A4 => 
                           n36567, ZN => n36554);
   U34671 : OAI22_X1 port map( A1 => n16914, A2 => n39295, B1 => n36534, B2 => 
                           n39291, ZN => n7174);
   U34672 : NOR2_X1 port map( A1 => n36535, A2 => n36536, ZN => n36534);
   U34673 : NAND4_X1 port map( A1 => n36537, A2 => n36538, A3 => n36539, A4 => 
                           n36540, ZN => n36536);
   U34674 : NAND4_X1 port map( A1 => n36545, A2 => n36546, A3 => n36547, A4 => 
                           n36548, ZN => n36535);
   U34675 : OAI22_X1 port map( A1 => n16915, A2 => n39295, B1 => n36515, B2 => 
                           n39291, ZN => n7175);
   U34676 : NOR2_X1 port map( A1 => n36516, A2 => n36517, ZN => n36515);
   U34677 : NAND4_X1 port map( A1 => n36518, A2 => n36519, A3 => n36520, A4 => 
                           n36521, ZN => n36517);
   U34678 : NAND4_X1 port map( A1 => n36526, A2 => n36527, A3 => n36528, A4 => 
                           n36529, ZN => n36516);
   U34679 : OAI22_X1 port map( A1 => n16916, A2 => n39295, B1 => n36496, B2 => 
                           n39291, ZN => n7176);
   U34680 : NOR2_X1 port map( A1 => n36497, A2 => n36498, ZN => n36496);
   U34681 : NAND4_X1 port map( A1 => n36499, A2 => n36500, A3 => n36501, A4 => 
                           n36502, ZN => n36498);
   U34682 : NAND4_X1 port map( A1 => n36507, A2 => n36508, A3 => n36509, A4 => 
                           n36510, ZN => n36497);
   U34683 : OAI22_X1 port map( A1 => n16917, A2 => n39295, B1 => n36477, B2 => 
                           n39291, ZN => n7177);
   U34684 : NOR2_X1 port map( A1 => n36478, A2 => n36479, ZN => n36477);
   U34685 : NAND4_X1 port map( A1 => n36480, A2 => n36481, A3 => n36482, A4 => 
                           n36483, ZN => n36479);
   U34686 : NAND4_X1 port map( A1 => n36488, A2 => n36489, A3 => n36490, A4 => 
                           n36491, ZN => n36478);
   U34687 : OAI22_X1 port map( A1 => n16918, A2 => n39295, B1 => n36458, B2 => 
                           n39291, ZN => n7178);
   U34688 : NOR2_X1 port map( A1 => n36459, A2 => n36460, ZN => n36458);
   U34689 : NAND4_X1 port map( A1 => n36461, A2 => n36462, A3 => n36463, A4 => 
                           n36464, ZN => n36460);
   U34690 : NAND4_X1 port map( A1 => n36469, A2 => n36470, A3 => n36471, A4 => 
                           n36472, ZN => n36459);
   U34691 : OAI22_X1 port map( A1 => n16919, A2 => n39294, B1 => n36439, B2 => 
                           n39291, ZN => n7179);
   U34692 : NOR2_X1 port map( A1 => n36440, A2 => n36441, ZN => n36439);
   U34693 : NAND4_X1 port map( A1 => n36442, A2 => n36443, A3 => n36444, A4 => 
                           n36445, ZN => n36441);
   U34694 : NAND4_X1 port map( A1 => n36450, A2 => n36451, A3 => n36452, A4 => 
                           n36453, ZN => n36440);
   U34695 : OAI22_X1 port map( A1 => n16920, A2 => n39294, B1 => n36420, B2 => 
                           n39291, ZN => n7180);
   U34696 : NOR2_X1 port map( A1 => n36421, A2 => n36422, ZN => n36420);
   U34697 : NAND4_X1 port map( A1 => n36423, A2 => n36424, A3 => n36425, A4 => 
                           n36426, ZN => n36422);
   U34698 : NAND4_X1 port map( A1 => n36431, A2 => n36432, A3 => n36433, A4 => 
                           n36434, ZN => n36421);
   U34699 : OAI22_X1 port map( A1 => n16921, A2 => n39294, B1 => n36401, B2 => 
                           n39291, ZN => n7181);
   U34700 : NOR2_X1 port map( A1 => n36402, A2 => n36403, ZN => n36401);
   U34701 : NAND4_X1 port map( A1 => n36404, A2 => n36405, A3 => n36406, A4 => 
                           n36407, ZN => n36403);
   U34702 : NAND4_X1 port map( A1 => n36412, A2 => n36413, A3 => n36414, A4 => 
                           n36415, ZN => n36402);
   U34703 : OAI22_X1 port map( A1 => n16922, A2 => n39294, B1 => n36382, B2 => 
                           n39291, ZN => n7182);
   U34704 : NOR2_X1 port map( A1 => n36383, A2 => n36384, ZN => n36382);
   U34705 : NAND4_X1 port map( A1 => n36385, A2 => n36386, A3 => n36387, A4 => 
                           n36388, ZN => n36384);
   U34706 : NAND4_X1 port map( A1 => n36393, A2 => n36394, A3 => n36395, A4 => 
                           n36396, ZN => n36383);
   U34707 : OAI22_X1 port map( A1 => n16923, A2 => n39294, B1 => n36363, B2 => 
                           n39291, ZN => n7183);
   U34708 : NOR2_X1 port map( A1 => n36364, A2 => n36365, ZN => n36363);
   U34709 : NAND4_X1 port map( A1 => n36366, A2 => n36367, A3 => n36368, A4 => 
                           n36369, ZN => n36365);
   U34710 : NAND4_X1 port map( A1 => n36374, A2 => n36375, A3 => n36376, A4 => 
                           n36377, ZN => n36364);
   U34711 : OAI22_X1 port map( A1 => n16924, A2 => n39294, B1 => n36344, B2 => 
                           n39291, ZN => n7184);
   U34712 : NOR2_X1 port map( A1 => n36345, A2 => n36346, ZN => n36344);
   U34713 : NAND4_X1 port map( A1 => n36347, A2 => n36348, A3 => n36349, A4 => 
                           n36350, ZN => n36346);
   U34714 : NAND4_X1 port map( A1 => n36355, A2 => n36356, A3 => n36357, A4 => 
                           n36358, ZN => n36345);
   U34715 : OAI22_X1 port map( A1 => n16925, A2 => n39294, B1 => n36325, B2 => 
                           n39291, ZN => n7185);
   U34716 : NOR2_X1 port map( A1 => n36326, A2 => n36327, ZN => n36325);
   U34717 : NAND4_X1 port map( A1 => n36328, A2 => n36329, A3 => n36330, A4 => 
                           n36331, ZN => n36327);
   U34718 : NAND4_X1 port map( A1 => n36336, A2 => n36337, A3 => n36338, A4 => 
                           n36339, ZN => n36326);
   U34719 : OAI22_X1 port map( A1 => n16926, A2 => n39294, B1 => n36306, B2 => 
                           n39292, ZN => n7186);
   U34720 : NOR2_X1 port map( A1 => n36307, A2 => n36308, ZN => n36306);
   U34721 : NAND4_X1 port map( A1 => n36309, A2 => n36310, A3 => n36311, A4 => 
                           n36312, ZN => n36308);
   U34722 : NAND4_X1 port map( A1 => n36317, A2 => n36318, A3 => n36319, A4 => 
                           n36320, ZN => n36307);
   U34723 : OAI22_X1 port map( A1 => n16927, A2 => n39295, B1 => n36287, B2 => 
                           n39292, ZN => n7187);
   U34724 : NOR2_X1 port map( A1 => n36288, A2 => n36289, ZN => n36287);
   U34725 : NAND4_X1 port map( A1 => n36290, A2 => n36291, A3 => n36292, A4 => 
                           n36293, ZN => n36289);
   U34726 : NAND4_X1 port map( A1 => n36298, A2 => n36299, A3 => n36300, A4 => 
                           n36301, ZN => n36288);
   U34727 : OAI22_X1 port map( A1 => n16928, A2 => n39294, B1 => n36268, B2 => 
                           n39292, ZN => n7188);
   U34728 : NOR2_X1 port map( A1 => n36269, A2 => n36270, ZN => n36268);
   U34729 : NAND4_X1 port map( A1 => n36271, A2 => n36272, A3 => n36273, A4 => 
                           n36274, ZN => n36270);
   U34730 : NAND4_X1 port map( A1 => n36279, A2 => n36280, A3 => n36281, A4 => 
                           n36282, ZN => n36269);
   U34731 : OAI22_X1 port map( A1 => n16929, A2 => n39294, B1 => n36249, B2 => 
                           n39292, ZN => n7189);
   U34732 : NOR2_X1 port map( A1 => n36250, A2 => n36251, ZN => n36249);
   U34733 : NAND4_X1 port map( A1 => n36252, A2 => n36253, A3 => n36254, A4 => 
                           n36255, ZN => n36251);
   U34734 : NAND4_X1 port map( A1 => n36260, A2 => n36261, A3 => n36262, A4 => 
                           n36263, ZN => n36250);
   U34735 : OAI22_X1 port map( A1 => n16930, A2 => n39294, B1 => n36230, B2 => 
                           n39292, ZN => n7190);
   U34736 : NOR2_X1 port map( A1 => n36231, A2 => n36232, ZN => n36230);
   U34737 : NAND4_X1 port map( A1 => n36233, A2 => n36234, A3 => n36235, A4 => 
                           n36236, ZN => n36232);
   U34738 : NAND4_X1 port map( A1 => n36241, A2 => n36242, A3 => n36243, A4 => 
                           n36244, ZN => n36231);
   U34739 : OAI22_X1 port map( A1 => n16931, A2 => n39294, B1 => n36211, B2 => 
                           n39292, ZN => n7191);
   U34740 : NOR2_X1 port map( A1 => n36212, A2 => n36213, ZN => n36211);
   U34741 : NAND4_X1 port map( A1 => n36214, A2 => n36215, A3 => n36216, A4 => 
                           n36217, ZN => n36213);
   U34742 : NAND4_X1 port map( A1 => n36222, A2 => n36223, A3 => n36224, A4 => 
                           n36225, ZN => n36212);
   U34743 : OAI22_X1 port map( A1 => n16879, A2 => n39295, B1 => n37199, B2 => 
                           n39288, ZN => n7139);
   U34744 : NOR2_X1 port map( A1 => n37200, A2 => n37201, ZN => n37199);
   U34745 : NAND4_X1 port map( A1 => n37202, A2 => n37203, A3 => n37204, A4 => 
                           n37205, ZN => n37201);
   U34746 : NAND4_X1 port map( A1 => n37210, A2 => n37211, A3 => n37212, A4 => 
                           n37213, ZN => n37200);
   U34747 : OAI22_X1 port map( A1 => n16880, A2 => n39294, B1 => n37180, B2 => 
                           n39288, ZN => n7140);
   U34748 : NOR2_X1 port map( A1 => n37181, A2 => n37182, ZN => n37180);
   U34749 : NAND4_X1 port map( A1 => n37183, A2 => n37184, A3 => n37185, A4 => 
                           n37186, ZN => n37182);
   U34750 : NAND4_X1 port map( A1 => n37191, A2 => n37192, A3 => n37193, A4 => 
                           n37194, ZN => n37181);
   U34751 : OAI22_X1 port map( A1 => n16881, A2 => n39296, B1 => n37161, B2 => 
                           n39288, ZN => n7141);
   U34752 : NOR2_X1 port map( A1 => n37162, A2 => n37163, ZN => n37161);
   U34753 : NAND4_X1 port map( A1 => n37164, A2 => n37165, A3 => n37166, A4 => 
                           n37167, ZN => n37163);
   U34754 : NAND4_X1 port map( A1 => n37172, A2 => n37173, A3 => n37174, A4 => 
                           n37175, ZN => n37162);
   U34755 : OAI22_X1 port map( A1 => n16882, A2 => n39295, B1 => n37142, B2 => 
                           n39288, ZN => n7142);
   U34756 : NOR2_X1 port map( A1 => n37143, A2 => n37144, ZN => n37142);
   U34757 : NAND4_X1 port map( A1 => n37145, A2 => n37146, A3 => n37147, A4 => 
                           n37148, ZN => n37144);
   U34758 : NAND4_X1 port map( A1 => n37153, A2 => n37154, A3 => n37155, A4 => 
                           n37156, ZN => n37143);
   U34759 : OAI22_X1 port map( A1 => n16883, A2 => n39294, B1 => n37123, B2 => 
                           n39288, ZN => n7143);
   U34760 : NOR2_X1 port map( A1 => n37124, A2 => n37125, ZN => n37123);
   U34761 : NAND4_X1 port map( A1 => n37126, A2 => n37127, A3 => n37128, A4 => 
                           n37129, ZN => n37125);
   U34762 : NAND4_X1 port map( A1 => n37134, A2 => n37135, A3 => n37136, A4 => 
                           n37137, ZN => n37124);
   U34763 : OAI22_X1 port map( A1 => n16884, A2 => n39296, B1 => n37104, B2 => 
                           n39288, ZN => n7144);
   U34764 : NOR2_X1 port map( A1 => n37105, A2 => n37106, ZN => n37104);
   U34765 : NAND4_X1 port map( A1 => n37107, A2 => n37108, A3 => n37109, A4 => 
                           n37110, ZN => n37106);
   U34766 : NAND4_X1 port map( A1 => n37115, A2 => n37116, A3 => n37117, A4 => 
                           n37118, ZN => n37105);
   U34767 : OAI22_X1 port map( A1 => n16885, A2 => n39296, B1 => n37085, B2 => 
                           n39288, ZN => n7145);
   U34768 : NOR2_X1 port map( A1 => n37086, A2 => n37087, ZN => n37085);
   U34769 : NAND4_X1 port map( A1 => n37088, A2 => n37089, A3 => n37090, A4 => 
                           n37091, ZN => n37087);
   U34770 : NAND4_X1 port map( A1 => n37096, A2 => n37097, A3 => n37098, A4 => 
                           n37099, ZN => n37086);
   U34771 : OAI22_X1 port map( A1 => n16886, A2 => n39296, B1 => n37066, B2 => 
                           n39288, ZN => n7146);
   U34772 : NOR2_X1 port map( A1 => n37067, A2 => n37068, ZN => n37066);
   U34773 : NAND4_X1 port map( A1 => n37069, A2 => n37070, A3 => n37071, A4 => 
                           n37072, ZN => n37068);
   U34774 : NAND4_X1 port map( A1 => n37077, A2 => n37078, A3 => n37079, A4 => 
                           n37080, ZN => n37067);
   U34775 : OAI22_X1 port map( A1 => n16887, A2 => n39296, B1 => n37047, B2 => 
                           n39288, ZN => n7147);
   U34776 : NOR2_X1 port map( A1 => n37048, A2 => n37049, ZN => n37047);
   U34777 : NAND4_X1 port map( A1 => n37050, A2 => n37051, A3 => n37052, A4 => 
                           n37053, ZN => n37049);
   U34778 : NAND4_X1 port map( A1 => n37058, A2 => n37059, A3 => n37060, A4 => 
                           n37061, ZN => n37048);
   U34779 : OAI22_X1 port map( A1 => n16888, A2 => n39296, B1 => n37028, B2 => 
                           n39288, ZN => n7148);
   U34780 : NOR2_X1 port map( A1 => n37029, A2 => n37030, ZN => n37028);
   U34781 : NAND4_X1 port map( A1 => n37031, A2 => n37032, A3 => n37033, A4 => 
                           n37034, ZN => n37030);
   U34782 : NAND4_X1 port map( A1 => n37039, A2 => n37040, A3 => n37041, A4 => 
                           n37042, ZN => n37029);
   U34783 : OAI22_X1 port map( A1 => n17065, A2 => n39801, B1 => n33542, B2 => 
                           n39794, ZN => n7326);
   U34784 : NOR2_X1 port map( A1 => n33543, A2 => n33544, ZN => n33542);
   U34785 : NAND4_X1 port map( A1 => n33545, A2 => n33546, A3 => n33547, A4 => 
                           n33548, ZN => n33544);
   U34786 : NAND4_X1 port map( A1 => n33553, A2 => n33554, A3 => n33555, A4 => 
                           n33556, ZN => n33543);
   U34787 : OAI22_X1 port map( A1 => n17001, A2 => n39549, B1 => n34816, B2 => 
                           n39542, ZN => n7262);
   U34788 : NOR2_X1 port map( A1 => n34817, A2 => n34818, ZN => n34816);
   U34789 : NAND4_X1 port map( A1 => n34819, A2 => n34820, A3 => n34821, A4 => 
                           n34822, ZN => n34818);
   U34790 : NAND4_X1 port map( A1 => n34827, A2 => n34828, A3 => n34829, A4 => 
                           n34830, ZN => n34817);
   U34791 : OAI22_X1 port map( A1 => n17064, A2 => n39800, B1 => n33561, B2 => 
                           n39794, ZN => n7325);
   U34792 : NOR2_X1 port map( A1 => n33562, A2 => n33563, ZN => n33561);
   U34793 : NAND4_X1 port map( A1 => n33564, A2 => n33565, A3 => n33566, A4 => 
                           n33567, ZN => n33563);
   U34794 : NAND4_X1 port map( A1 => n33572, A2 => n33573, A3 => n33574, A4 => 
                           n33575, ZN => n33562);
   U34795 : OAI22_X1 port map( A1 => n17000, A2 => n39548, B1 => n34835, B2 => 
                           n39542, ZN => n7261);
   U34796 : NOR2_X1 port map( A1 => n34836, A2 => n34837, ZN => n34835);
   U34797 : NAND4_X1 port map( A1 => n34838, A2 => n34839, A3 => n34840, A4 => 
                           n34841, ZN => n34837);
   U34798 : NAND4_X1 port map( A1 => n34846, A2 => n34847, A3 => n34848, A4 => 
                           n34849, ZN => n34836);
   U34799 : OAI22_X1 port map( A1 => n17063, A2 => n39800, B1 => n33580, B2 => 
                           n39794, ZN => n7324);
   U34800 : NOR2_X1 port map( A1 => n33581, A2 => n33582, ZN => n33580);
   U34801 : NAND4_X1 port map( A1 => n33583, A2 => n33584, A3 => n33585, A4 => 
                           n33586, ZN => n33582);
   U34802 : NAND4_X1 port map( A1 => n33591, A2 => n33592, A3 => n33593, A4 => 
                           n33594, ZN => n33581);
   U34803 : OAI22_X1 port map( A1 => n16999, A2 => n39548, B1 => n34854, B2 => 
                           n39542, ZN => n7260);
   U34804 : NOR2_X1 port map( A1 => n34855, A2 => n34856, ZN => n34854);
   U34805 : NAND4_X1 port map( A1 => n34857, A2 => n34858, A3 => n34859, A4 => 
                           n34860, ZN => n34856);
   U34806 : NAND4_X1 port map( A1 => n34865, A2 => n34866, A3 => n34867, A4 => 
                           n34868, ZN => n34855);
   U34807 : OAI22_X1 port map( A1 => n17062, A2 => n39800, B1 => n33599, B2 => 
                           n39794, ZN => n7323);
   U34808 : NOR2_X1 port map( A1 => n33600, A2 => n33601, ZN => n33599);
   U34809 : NAND4_X1 port map( A1 => n33602, A2 => n33603, A3 => n33604, A4 => 
                           n33605, ZN => n33601);
   U34810 : NAND4_X1 port map( A1 => n33610, A2 => n33611, A3 => n33612, A4 => 
                           n33613, ZN => n33600);
   U34811 : OAI22_X1 port map( A1 => n16998, A2 => n39548, B1 => n34873, B2 => 
                           n39542, ZN => n7259);
   U34812 : NOR2_X1 port map( A1 => n34874, A2 => n34875, ZN => n34873);
   U34813 : NAND4_X1 port map( A1 => n34876, A2 => n34877, A3 => n34878, A4 => 
                           n34879, ZN => n34875);
   U34814 : NAND4_X1 port map( A1 => n34884, A2 => n34885, A3 => n34886, A4 => 
                           n34887, ZN => n34874);
   U34815 : OAI22_X1 port map( A1 => n17061, A2 => n39800, B1 => n33618, B2 => 
                           n39794, ZN => n7322);
   U34816 : NOR2_X1 port map( A1 => n33619, A2 => n33620, ZN => n33618);
   U34817 : NAND4_X1 port map( A1 => n33621, A2 => n33622, A3 => n33623, A4 => 
                           n33624, ZN => n33620);
   U34818 : NAND4_X1 port map( A1 => n33629, A2 => n33630, A3 => n33631, A4 => 
                           n33632, ZN => n33619);
   U34819 : OAI22_X1 port map( A1 => n16997, A2 => n39548, B1 => n34892, B2 => 
                           n39542, ZN => n7258);
   U34820 : NOR2_X1 port map( A1 => n34893, A2 => n34894, ZN => n34892);
   U34821 : NAND4_X1 port map( A1 => n34895, A2 => n34896, A3 => n34897, A4 => 
                           n34898, ZN => n34894);
   U34822 : NAND4_X1 port map( A1 => n34903, A2 => n34904, A3 => n34905, A4 => 
                           n34906, ZN => n34893);
   U34823 : OAI22_X1 port map( A1 => n17060, A2 => n39800, B1 => n33637, B2 => 
                           n39794, ZN => n7321);
   U34824 : NOR2_X1 port map( A1 => n33638, A2 => n33639, ZN => n33637);
   U34825 : NAND4_X1 port map( A1 => n33640, A2 => n33641, A3 => n33642, A4 => 
                           n33643, ZN => n33639);
   U34826 : NAND4_X1 port map( A1 => n33648, A2 => n33649, A3 => n33650, A4 => 
                           n33651, ZN => n33638);
   U34827 : OAI22_X1 port map( A1 => n16996, A2 => n39548, B1 => n34911, B2 => 
                           n39542, ZN => n7257);
   U34828 : NOR2_X1 port map( A1 => n34912, A2 => n34913, ZN => n34911);
   U34829 : NAND4_X1 port map( A1 => n34914, A2 => n34915, A3 => n34916, A4 => 
                           n34917, ZN => n34913);
   U34830 : NAND4_X1 port map( A1 => n34922, A2 => n34923, A3 => n34924, A4 => 
                           n34925, ZN => n34912);
   U34831 : OAI22_X1 port map( A1 => n17059, A2 => n39800, B1 => n33656, B2 => 
                           n39794, ZN => n7320);
   U34832 : NOR2_X1 port map( A1 => n33657, A2 => n33658, ZN => n33656);
   U34833 : NAND4_X1 port map( A1 => n33659, A2 => n33660, A3 => n33661, A4 => 
                           n33662, ZN => n33658);
   U34834 : NAND4_X1 port map( A1 => n33667, A2 => n33668, A3 => n33669, A4 => 
                           n33670, ZN => n33657);
   U34835 : OAI22_X1 port map( A1 => n16995, A2 => n39548, B1 => n34930, B2 => 
                           n39542, ZN => n7256);
   U34836 : NOR2_X1 port map( A1 => n34931, A2 => n34932, ZN => n34930);
   U34837 : NAND4_X1 port map( A1 => n34933, A2 => n34934, A3 => n34935, A4 => 
                           n34936, ZN => n34932);
   U34838 : NAND4_X1 port map( A1 => n34941, A2 => n34942, A3 => n34943, A4 => 
                           n34944, ZN => n34931);
   U34839 : OAI22_X1 port map( A1 => n17058, A2 => n39800, B1 => n33675, B2 => 
                           n39794, ZN => n7319);
   U34840 : NOR2_X1 port map( A1 => n33676, A2 => n33677, ZN => n33675);
   U34841 : NAND4_X1 port map( A1 => n33678, A2 => n33679, A3 => n33680, A4 => 
                           n33681, ZN => n33677);
   U34842 : NAND4_X1 port map( A1 => n33686, A2 => n33687, A3 => n33688, A4 => 
                           n33689, ZN => n33676);
   U34843 : OAI22_X1 port map( A1 => n16994, A2 => n39548, B1 => n34949, B2 => 
                           n39542, ZN => n7255);
   U34844 : NOR2_X1 port map( A1 => n34950, A2 => n34951, ZN => n34949);
   U34845 : NAND4_X1 port map( A1 => n34952, A2 => n34953, A3 => n34954, A4 => 
                           n34955, ZN => n34951);
   U34846 : NAND4_X1 port map( A1 => n34960, A2 => n34961, A3 => n34962, A4 => 
                           n34963, ZN => n34950);
   U34847 : OAI22_X1 port map( A1 => n17057, A2 => n39800, B1 => n33694, B2 => 
                           n39794, ZN => n7318);
   U34848 : NOR2_X1 port map( A1 => n33695, A2 => n33696, ZN => n33694);
   U34849 : NAND4_X1 port map( A1 => n33697, A2 => n33698, A3 => n33699, A4 => 
                           n33700, ZN => n33696);
   U34850 : NAND4_X1 port map( A1 => n33705, A2 => n33706, A3 => n33707, A4 => 
                           n33708, ZN => n33695);
   U34851 : OAI22_X1 port map( A1 => n16993, A2 => n39548, B1 => n34968, B2 => 
                           n39542, ZN => n7254);
   U34852 : NOR2_X1 port map( A1 => n34969, A2 => n34970, ZN => n34968);
   U34853 : NAND4_X1 port map( A1 => n34971, A2 => n34972, A3 => n34973, A4 => 
                           n34974, ZN => n34970);
   U34854 : NAND4_X1 port map( A1 => n34979, A2 => n34980, A3 => n34981, A4 => 
                           n34982, ZN => n34969);
   U34855 : OAI22_X1 port map( A1 => n17056, A2 => n39800, B1 => n33713, B2 => 
                           n39794, ZN => n7317);
   U34856 : NOR2_X1 port map( A1 => n33714, A2 => n33715, ZN => n33713);
   U34857 : NAND4_X1 port map( A1 => n33716, A2 => n33717, A3 => n33718, A4 => 
                           n33719, ZN => n33715);
   U34858 : NAND4_X1 port map( A1 => n33724, A2 => n33725, A3 => n33726, A4 => 
                           n33727, ZN => n33714);
   U34859 : OAI22_X1 port map( A1 => n16992, A2 => n39548, B1 => n34987, B2 => 
                           n39542, ZN => n7253);
   U34860 : NOR2_X1 port map( A1 => n34988, A2 => n34989, ZN => n34987);
   U34861 : NAND4_X1 port map( A1 => n34990, A2 => n34991, A3 => n34992, A4 => 
                           n34993, ZN => n34989);
   U34862 : NAND4_X1 port map( A1 => n34998, A2 => n34999, A3 => n35000, A4 => 
                           n35001, ZN => n34988);
   U34863 : OAI22_X1 port map( A1 => n17055, A2 => n39800, B1 => n33732, B2 => 
                           n39794, ZN => n7316);
   U34864 : NOR2_X1 port map( A1 => n33733, A2 => n33734, ZN => n33732);
   U34865 : NAND4_X1 port map( A1 => n33735, A2 => n33736, A3 => n33737, A4 => 
                           n33738, ZN => n33734);
   U34866 : NAND4_X1 port map( A1 => n33743, A2 => n33744, A3 => n33745, A4 => 
                           n33746, ZN => n33733);
   U34867 : OAI22_X1 port map( A1 => n16991, A2 => n39548, B1 => n35006, B2 => 
                           n39542, ZN => n7252);
   U34868 : NOR2_X1 port map( A1 => n35007, A2 => n35008, ZN => n35006);
   U34869 : NAND4_X1 port map( A1 => n35009, A2 => n35010, A3 => n35011, A4 => 
                           n35012, ZN => n35008);
   U34870 : NAND4_X1 port map( A1 => n35017, A2 => n35018, A3 => n35019, A4 => 
                           n35020, ZN => n35007);
   U34871 : OAI22_X1 port map( A1 => n17054, A2 => n39800, B1 => n33751, B2 => 
                           n39794, ZN => n7315);
   U34872 : NOR2_X1 port map( A1 => n33752, A2 => n33753, ZN => n33751);
   U34873 : NAND4_X1 port map( A1 => n33754, A2 => n33755, A3 => n33756, A4 => 
                           n33757, ZN => n33753);
   U34874 : NAND4_X1 port map( A1 => n33762, A2 => n33763, A3 => n33764, A4 => 
                           n33765, ZN => n33752);
   U34875 : OAI22_X1 port map( A1 => n16990, A2 => n39548, B1 => n35025, B2 => 
                           n39542, ZN => n7251);
   U34876 : NOR2_X1 port map( A1 => n35026, A2 => n35027, ZN => n35025);
   U34877 : NAND4_X1 port map( A1 => n35028, A2 => n35029, A3 => n35030, A4 => 
                           n35031, ZN => n35027);
   U34878 : NAND4_X1 port map( A1 => n35036, A2 => n35037, A3 => n35038, A4 => 
                           n35039, ZN => n35026);
   U34879 : OAI22_X1 port map( A1 => n17053, A2 => n39800, B1 => n33770, B2 => 
                           n39793, ZN => n7314);
   U34880 : NOR2_X1 port map( A1 => n33771, A2 => n33772, ZN => n33770);
   U34881 : NAND4_X1 port map( A1 => n33773, A2 => n33774, A3 => n33775, A4 => 
                           n33776, ZN => n33772);
   U34882 : NAND4_X1 port map( A1 => n33781, A2 => n33782, A3 => n33783, A4 => 
                           n33784, ZN => n33771);
   U34883 : OAI22_X1 port map( A1 => n16989, A2 => n39548, B1 => n35044, B2 => 
                           n39541, ZN => n7250);
   U34884 : NOR2_X1 port map( A1 => n35045, A2 => n35046, ZN => n35044);
   U34885 : NAND4_X1 port map( A1 => n35047, A2 => n35048, A3 => n35049, A4 => 
                           n35050, ZN => n35046);
   U34886 : NAND4_X1 port map( A1 => n35055, A2 => n35056, A3 => n35057, A4 => 
                           n35058, ZN => n35045);
   U34887 : OAI22_X1 port map( A1 => n17052, A2 => n39799, B1 => n33789, B2 => 
                           n39793, ZN => n7313);
   U34888 : NOR2_X1 port map( A1 => n33790, A2 => n33791, ZN => n33789);
   U34889 : NAND4_X1 port map( A1 => n33792, A2 => n33793, A3 => n33794, A4 => 
                           n33795, ZN => n33791);
   U34890 : NAND4_X1 port map( A1 => n33800, A2 => n33801, A3 => n33802, A4 => 
                           n33803, ZN => n33790);
   U34891 : OAI22_X1 port map( A1 => n16988, A2 => n39547, B1 => n35063, B2 => 
                           n39541, ZN => n7249);
   U34892 : NOR2_X1 port map( A1 => n35064, A2 => n35065, ZN => n35063);
   U34893 : NAND4_X1 port map( A1 => n35066, A2 => n35067, A3 => n35068, A4 => 
                           n35069, ZN => n35065);
   U34894 : NAND4_X1 port map( A1 => n35074, A2 => n35075, A3 => n35076, A4 => 
                           n35077, ZN => n35064);
   U34895 : OAI22_X1 port map( A1 => n17051, A2 => n39799, B1 => n33808, B2 => 
                           n39793, ZN => n7312);
   U34896 : NOR2_X1 port map( A1 => n33809, A2 => n33810, ZN => n33808);
   U34897 : NAND4_X1 port map( A1 => n33811, A2 => n33812, A3 => n33813, A4 => 
                           n33814, ZN => n33810);
   U34898 : NAND4_X1 port map( A1 => n33819, A2 => n33820, A3 => n33821, A4 => 
                           n33822, ZN => n33809);
   U34899 : OAI22_X1 port map( A1 => n16987, A2 => n39547, B1 => n35082, B2 => 
                           n39541, ZN => n7248);
   U34900 : NOR2_X1 port map( A1 => n35083, A2 => n35084, ZN => n35082);
   U34901 : NAND4_X1 port map( A1 => n35085, A2 => n35086, A3 => n35087, A4 => 
                           n35088, ZN => n35084);
   U34902 : NAND4_X1 port map( A1 => n35093, A2 => n35094, A3 => n35095, A4 => 
                           n35096, ZN => n35083);
   U34903 : OAI22_X1 port map( A1 => n17050, A2 => n39799, B1 => n33827, B2 => 
                           n39793, ZN => n7311);
   U34904 : NOR2_X1 port map( A1 => n33828, A2 => n33829, ZN => n33827);
   U34905 : NAND4_X1 port map( A1 => n33830, A2 => n33831, A3 => n33832, A4 => 
                           n33833, ZN => n33829);
   U34906 : NAND4_X1 port map( A1 => n33838, A2 => n33839, A3 => n33840, A4 => 
                           n33841, ZN => n33828);
   U34907 : OAI22_X1 port map( A1 => n16986, A2 => n39547, B1 => n35101, B2 => 
                           n39541, ZN => n7247);
   U34908 : NOR2_X1 port map( A1 => n35102, A2 => n35103, ZN => n35101);
   U34909 : NAND4_X1 port map( A1 => n35104, A2 => n35105, A3 => n35106, A4 => 
                           n35107, ZN => n35103);
   U34910 : NAND4_X1 port map( A1 => n35112, A2 => n35113, A3 => n35114, A4 => 
                           n35115, ZN => n35102);
   U34911 : OAI22_X1 port map( A1 => n17049, A2 => n39799, B1 => n33846, B2 => 
                           n39793, ZN => n7310);
   U34912 : NOR2_X1 port map( A1 => n33847, A2 => n33848, ZN => n33846);
   U34913 : NAND4_X1 port map( A1 => n33849, A2 => n33850, A3 => n33851, A4 => 
                           n33852, ZN => n33848);
   U34914 : NAND4_X1 port map( A1 => n33857, A2 => n33858, A3 => n33859, A4 => 
                           n33860, ZN => n33847);
   U34915 : OAI22_X1 port map( A1 => n16985, A2 => n39547, B1 => n35120, B2 => 
                           n39541, ZN => n7246);
   U34916 : NOR2_X1 port map( A1 => n35121, A2 => n35122, ZN => n35120);
   U34917 : NAND4_X1 port map( A1 => n35123, A2 => n35124, A3 => n35125, A4 => 
                           n35126, ZN => n35122);
   U34918 : NAND4_X1 port map( A1 => n35131, A2 => n35132, A3 => n35133, A4 => 
                           n35134, ZN => n35121);
   U34919 : OAI22_X1 port map( A1 => n17048, A2 => n39799, B1 => n33865, B2 => 
                           n39793, ZN => n7309);
   U34920 : NOR2_X1 port map( A1 => n33866, A2 => n33867, ZN => n33865);
   U34921 : NAND4_X1 port map( A1 => n33868, A2 => n33869, A3 => n33870, A4 => 
                           n33871, ZN => n33867);
   U34922 : NAND4_X1 port map( A1 => n33876, A2 => n33877, A3 => n33878, A4 => 
                           n33879, ZN => n33866);
   U34923 : OAI22_X1 port map( A1 => n16984, A2 => n39547, B1 => n35139, B2 => 
                           n39541, ZN => n7245);
   U34924 : NOR2_X1 port map( A1 => n35140, A2 => n35141, ZN => n35139);
   U34925 : NAND4_X1 port map( A1 => n35142, A2 => n35143, A3 => n35144, A4 => 
                           n35145, ZN => n35141);
   U34926 : NAND4_X1 port map( A1 => n35150, A2 => n35151, A3 => n35152, A4 => 
                           n35153, ZN => n35140);
   U34927 : OAI22_X1 port map( A1 => n17047, A2 => n39799, B1 => n33884, B2 => 
                           n39793, ZN => n7308);
   U34928 : NOR2_X1 port map( A1 => n33885, A2 => n33886, ZN => n33884);
   U34929 : NAND4_X1 port map( A1 => n33887, A2 => n33888, A3 => n33889, A4 => 
                           n33890, ZN => n33886);
   U34930 : NAND4_X1 port map( A1 => n33895, A2 => n33896, A3 => n33897, A4 => 
                           n33898, ZN => n33885);
   U34931 : OAI22_X1 port map( A1 => n16983, A2 => n39547, B1 => n35158, B2 => 
                           n39541, ZN => n7244);
   U34932 : NOR2_X1 port map( A1 => n35159, A2 => n35160, ZN => n35158);
   U34933 : NAND4_X1 port map( A1 => n35161, A2 => n35162, A3 => n35163, A4 => 
                           n35164, ZN => n35160);
   U34934 : NAND4_X1 port map( A1 => n35169, A2 => n35170, A3 => n35171, A4 => 
                           n35172, ZN => n35159);
   U34935 : OAI22_X1 port map( A1 => n17046, A2 => n39799, B1 => n33903, B2 => 
                           n39793, ZN => n7307);
   U34936 : NOR2_X1 port map( A1 => n33904, A2 => n33905, ZN => n33903);
   U34937 : NAND4_X1 port map( A1 => n33906, A2 => n33907, A3 => n33908, A4 => 
                           n33909, ZN => n33905);
   U34938 : NAND4_X1 port map( A1 => n33914, A2 => n33915, A3 => n33916, A4 => 
                           n33917, ZN => n33904);
   U34939 : OAI22_X1 port map( A1 => n16982, A2 => n39547, B1 => n35177, B2 => 
                           n39541, ZN => n7243);
   U34940 : NOR2_X1 port map( A1 => n35178, A2 => n35179, ZN => n35177);
   U34941 : NAND4_X1 port map( A1 => n35180, A2 => n35181, A3 => n35182, A4 => 
                           n35183, ZN => n35179);
   U34942 : NAND4_X1 port map( A1 => n35188, A2 => n35189, A3 => n35190, A4 => 
                           n35191, ZN => n35178);
   U34943 : OAI22_X1 port map( A1 => n17045, A2 => n39799, B1 => n33922, B2 => 
                           n39793, ZN => n7306);
   U34944 : NOR2_X1 port map( A1 => n33923, A2 => n33924, ZN => n33922);
   U34945 : NAND4_X1 port map( A1 => n33925, A2 => n33926, A3 => n33927, A4 => 
                           n33928, ZN => n33924);
   U34946 : NAND4_X1 port map( A1 => n33933, A2 => n33934, A3 => n33935, A4 => 
                           n33936, ZN => n33923);
   U34947 : OAI22_X1 port map( A1 => n16981, A2 => n39547, B1 => n35196, B2 => 
                           n39541, ZN => n7242);
   U34948 : NOR2_X1 port map( A1 => n35197, A2 => n35198, ZN => n35196);
   U34949 : NAND4_X1 port map( A1 => n35199, A2 => n35200, A3 => n35201, A4 => 
                           n35202, ZN => n35198);
   U34950 : NAND4_X1 port map( A1 => n35207, A2 => n35208, A3 => n35209, A4 => 
                           n35210, ZN => n35197);
   U34951 : OAI22_X1 port map( A1 => n17044, A2 => n39799, B1 => n33941, B2 => 
                           n39793, ZN => n7305);
   U34952 : NOR2_X1 port map( A1 => n33942, A2 => n33943, ZN => n33941);
   U34953 : NAND4_X1 port map( A1 => n33944, A2 => n33945, A3 => n33946, A4 => 
                           n33947, ZN => n33943);
   U34954 : NAND4_X1 port map( A1 => n33952, A2 => n33953, A3 => n33954, A4 => 
                           n33955, ZN => n33942);
   U34955 : OAI22_X1 port map( A1 => n16980, A2 => n39547, B1 => n35215, B2 => 
                           n39541, ZN => n7241);
   U34956 : NOR2_X1 port map( A1 => n35216, A2 => n35217, ZN => n35215);
   U34957 : NAND4_X1 port map( A1 => n35218, A2 => n35219, A3 => n35220, A4 => 
                           n35221, ZN => n35217);
   U34958 : NAND4_X1 port map( A1 => n35226, A2 => n35227, A3 => n35228, A4 => 
                           n35229, ZN => n35216);
   U34959 : OAI22_X1 port map( A1 => n17043, A2 => n39799, B1 => n33960, B2 => 
                           n39793, ZN => n7304);
   U34960 : NOR2_X1 port map( A1 => n33961, A2 => n33962, ZN => n33960);
   U34961 : NAND4_X1 port map( A1 => n33963, A2 => n33964, A3 => n33965, A4 => 
                           n33966, ZN => n33962);
   U34962 : NAND4_X1 port map( A1 => n33971, A2 => n33972, A3 => n33973, A4 => 
                           n33974, ZN => n33961);
   U34963 : OAI22_X1 port map( A1 => n16979, A2 => n39547, B1 => n35234, B2 => 
                           n39541, ZN => n7240);
   U34964 : NOR2_X1 port map( A1 => n35235, A2 => n35236, ZN => n35234);
   U34965 : NAND4_X1 port map( A1 => n35237, A2 => n35238, A3 => n35239, A4 => 
                           n35240, ZN => n35236);
   U34966 : NAND4_X1 port map( A1 => n35245, A2 => n35246, A3 => n35247, A4 => 
                           n35248, ZN => n35235);
   U34967 : OAI22_X1 port map( A1 => n17042, A2 => n39799, B1 => n33979, B2 => 
                           n39793, ZN => n7303);
   U34968 : NOR2_X1 port map( A1 => n33980, A2 => n33981, ZN => n33979);
   U34969 : NAND4_X1 port map( A1 => n33982, A2 => n33983, A3 => n33984, A4 => 
                           n33985, ZN => n33981);
   U34970 : NAND4_X1 port map( A1 => n33990, A2 => n33991, A3 => n33992, A4 => 
                           n33993, ZN => n33980);
   U34971 : OAI22_X1 port map( A1 => n16978, A2 => n39547, B1 => n35253, B2 => 
                           n39541, ZN => n7239);
   U34972 : NOR2_X1 port map( A1 => n35254, A2 => n35255, ZN => n35253);
   U34973 : NAND4_X1 port map( A1 => n35256, A2 => n35257, A3 => n35258, A4 => 
                           n35259, ZN => n35255);
   U34974 : NAND4_X1 port map( A1 => n35264, A2 => n35265, A3 => n35266, A4 => 
                           n35267, ZN => n35254);
   U34975 : OAI22_X1 port map( A1 => n17041, A2 => n39799, B1 => n33998, B2 => 
                           n39792, ZN => n7302);
   U34976 : NOR2_X1 port map( A1 => n33999, A2 => n34000, ZN => n33998);
   U34977 : NAND4_X1 port map( A1 => n34001, A2 => n34002, A3 => n34003, A4 => 
                           n34004, ZN => n34000);
   U34978 : NAND4_X1 port map( A1 => n34009, A2 => n34010, A3 => n34011, A4 => 
                           n34012, ZN => n33999);
   U34979 : OAI22_X1 port map( A1 => n16977, A2 => n39547, B1 => n35272, B2 => 
                           n39540, ZN => n7238);
   U34980 : NOR2_X1 port map( A1 => n35273, A2 => n35274, ZN => n35272);
   U34981 : NAND4_X1 port map( A1 => n35275, A2 => n35276, A3 => n35277, A4 => 
                           n35278, ZN => n35274);
   U34982 : NAND4_X1 port map( A1 => n35283, A2 => n35284, A3 => n35285, A4 => 
                           n35286, ZN => n35273);
   U34983 : OAI22_X1 port map( A1 => n17040, A2 => n39798, B1 => n34017, B2 => 
                           n39792, ZN => n7301);
   U34984 : NOR2_X1 port map( A1 => n34018, A2 => n34019, ZN => n34017);
   U34985 : NAND4_X1 port map( A1 => n34020, A2 => n34021, A3 => n34022, A4 => 
                           n34023, ZN => n34019);
   U34986 : NAND4_X1 port map( A1 => n34028, A2 => n34029, A3 => n34030, A4 => 
                           n34031, ZN => n34018);
   U34987 : OAI22_X1 port map( A1 => n16976, A2 => n39546, B1 => n35291, B2 => 
                           n39540, ZN => n7237);
   U34988 : NOR2_X1 port map( A1 => n35292, A2 => n35293, ZN => n35291);
   U34989 : NAND4_X1 port map( A1 => n35294, A2 => n35295, A3 => n35296, A4 => 
                           n35297, ZN => n35293);
   U34990 : NAND4_X1 port map( A1 => n35302, A2 => n35303, A3 => n35304, A4 => 
                           n35305, ZN => n35292);
   U34991 : OAI22_X1 port map( A1 => n17039, A2 => n39798, B1 => n34036, B2 => 
                           n39792, ZN => n7300);
   U34992 : NOR2_X1 port map( A1 => n34037, A2 => n34038, ZN => n34036);
   U34993 : NAND4_X1 port map( A1 => n34039, A2 => n34040, A3 => n34041, A4 => 
                           n34042, ZN => n34038);
   U34994 : NAND4_X1 port map( A1 => n34047, A2 => n34048, A3 => n34049, A4 => 
                           n34050, ZN => n34037);
   U34995 : OAI22_X1 port map( A1 => n16975, A2 => n39546, B1 => n35310, B2 => 
                           n39540, ZN => n7236);
   U34996 : NOR2_X1 port map( A1 => n35311, A2 => n35312, ZN => n35310);
   U34997 : NAND4_X1 port map( A1 => n35313, A2 => n35314, A3 => n35315, A4 => 
                           n35316, ZN => n35312);
   U34998 : NAND4_X1 port map( A1 => n35321, A2 => n35322, A3 => n35323, A4 => 
                           n35324, ZN => n35311);
   U34999 : OAI22_X1 port map( A1 => n17038, A2 => n39798, B1 => n34055, B2 => 
                           n39792, ZN => n7299);
   U35000 : NOR2_X1 port map( A1 => n34056, A2 => n34057, ZN => n34055);
   U35001 : NAND4_X1 port map( A1 => n34058, A2 => n34059, A3 => n34060, A4 => 
                           n34061, ZN => n34057);
   U35002 : NAND4_X1 port map( A1 => n34066, A2 => n34067, A3 => n34068, A4 => 
                           n34069, ZN => n34056);
   U35003 : OAI22_X1 port map( A1 => n16974, A2 => n39546, B1 => n35329, B2 => 
                           n39540, ZN => n7235);
   U35004 : NOR2_X1 port map( A1 => n35330, A2 => n35331, ZN => n35329);
   U35005 : NAND4_X1 port map( A1 => n35332, A2 => n35333, A3 => n35334, A4 => 
                           n35335, ZN => n35331);
   U35006 : NAND4_X1 port map( A1 => n35340, A2 => n35341, A3 => n35342, A4 => 
                           n35343, ZN => n35330);
   U35007 : OAI22_X1 port map( A1 => n17037, A2 => n39798, B1 => n34074, B2 => 
                           n39792, ZN => n7298);
   U35008 : NOR2_X1 port map( A1 => n34075, A2 => n34076, ZN => n34074);
   U35009 : NAND4_X1 port map( A1 => n34077, A2 => n34078, A3 => n34079, A4 => 
                           n34080, ZN => n34076);
   U35010 : NAND4_X1 port map( A1 => n34085, A2 => n34086, A3 => n34087, A4 => 
                           n34088, ZN => n34075);
   U35011 : OAI22_X1 port map( A1 => n16973, A2 => n39546, B1 => n35348, B2 => 
                           n39540, ZN => n7234);
   U35012 : NOR2_X1 port map( A1 => n35349, A2 => n35350, ZN => n35348);
   U35013 : NAND4_X1 port map( A1 => n35351, A2 => n35352, A3 => n35353, A4 => 
                           n35354, ZN => n35350);
   U35014 : NAND4_X1 port map( A1 => n35359, A2 => n35360, A3 => n35361, A4 => 
                           n35362, ZN => n35349);
   U35015 : OAI22_X1 port map( A1 => n17036, A2 => n39798, B1 => n34093, B2 => 
                           n39792, ZN => n7297);
   U35016 : NOR2_X1 port map( A1 => n34094, A2 => n34095, ZN => n34093);
   U35017 : NAND4_X1 port map( A1 => n34096, A2 => n34097, A3 => n34098, A4 => 
                           n34099, ZN => n34095);
   U35018 : NAND4_X1 port map( A1 => n34104, A2 => n34105, A3 => n34106, A4 => 
                           n34107, ZN => n34094);
   U35019 : OAI22_X1 port map( A1 => n16972, A2 => n39546, B1 => n35367, B2 => 
                           n39540, ZN => n7233);
   U35020 : NOR2_X1 port map( A1 => n35368, A2 => n35369, ZN => n35367);
   U35021 : NAND4_X1 port map( A1 => n35370, A2 => n35371, A3 => n35372, A4 => 
                           n35373, ZN => n35369);
   U35022 : NAND4_X1 port map( A1 => n35378, A2 => n35379, A3 => n35380, A4 => 
                           n35381, ZN => n35368);
   U35023 : OAI22_X1 port map( A1 => n17035, A2 => n39798, B1 => n34112, B2 => 
                           n39792, ZN => n7296);
   U35024 : NOR2_X1 port map( A1 => n34113, A2 => n34114, ZN => n34112);
   U35025 : NAND4_X1 port map( A1 => n34115, A2 => n34116, A3 => n34117, A4 => 
                           n34118, ZN => n34114);
   U35026 : NAND4_X1 port map( A1 => n34123, A2 => n34124, A3 => n34125, A4 => 
                           n34126, ZN => n34113);
   U35027 : OAI22_X1 port map( A1 => n16971, A2 => n39546, B1 => n35386, B2 => 
                           n39540, ZN => n7232);
   U35028 : NOR2_X1 port map( A1 => n35387, A2 => n35388, ZN => n35386);
   U35029 : NAND4_X1 port map( A1 => n35389, A2 => n35390, A3 => n35391, A4 => 
                           n35392, ZN => n35388);
   U35030 : NAND4_X1 port map( A1 => n35397, A2 => n35398, A3 => n35399, A4 => 
                           n35400, ZN => n35387);
   U35031 : OAI22_X1 port map( A1 => n17034, A2 => n39798, B1 => n34131, B2 => 
                           n39792, ZN => n7295);
   U35032 : NOR2_X1 port map( A1 => n34132, A2 => n34133, ZN => n34131);
   U35033 : NAND4_X1 port map( A1 => n34134, A2 => n34135, A3 => n34136, A4 => 
                           n34137, ZN => n34133);
   U35034 : NAND4_X1 port map( A1 => n34142, A2 => n34143, A3 => n34144, A4 => 
                           n34145, ZN => n34132);
   U35035 : OAI22_X1 port map( A1 => n16970, A2 => n39546, B1 => n35405, B2 => 
                           n39540, ZN => n7231);
   U35036 : NOR2_X1 port map( A1 => n35406, A2 => n35407, ZN => n35405);
   U35037 : NAND4_X1 port map( A1 => n35408, A2 => n35409, A3 => n35410, A4 => 
                           n35411, ZN => n35407);
   U35038 : NAND4_X1 port map( A1 => n35416, A2 => n35417, A3 => n35418, A4 => 
                           n35419, ZN => n35406);
   U35039 : OAI22_X1 port map( A1 => n17033, A2 => n39798, B1 => n34150, B2 => 
                           n39792, ZN => n7294);
   U35040 : NOR2_X1 port map( A1 => n34151, A2 => n34152, ZN => n34150);
   U35041 : NAND4_X1 port map( A1 => n34153, A2 => n34154, A3 => n34155, A4 => 
                           n34156, ZN => n34152);
   U35042 : NAND4_X1 port map( A1 => n34161, A2 => n34162, A3 => n34163, A4 => 
                           n34164, ZN => n34151);
   U35043 : OAI22_X1 port map( A1 => n16969, A2 => n39546, B1 => n35424, B2 => 
                           n39540, ZN => n7230);
   U35044 : NOR2_X1 port map( A1 => n35425, A2 => n35426, ZN => n35424);
   U35045 : NAND4_X1 port map( A1 => n35427, A2 => n35428, A3 => n35429, A4 => 
                           n35430, ZN => n35426);
   U35046 : NAND4_X1 port map( A1 => n35435, A2 => n35436, A3 => n35437, A4 => 
                           n35438, ZN => n35425);
   U35047 : OAI22_X1 port map( A1 => n17032, A2 => n39798, B1 => n34169, B2 => 
                           n39792, ZN => n7293);
   U35048 : NOR2_X1 port map( A1 => n34170, A2 => n34171, ZN => n34169);
   U35049 : NAND4_X1 port map( A1 => n34172, A2 => n34173, A3 => n34174, A4 => 
                           n34175, ZN => n34171);
   U35050 : NAND4_X1 port map( A1 => n34180, A2 => n34181, A3 => n34182, A4 => 
                           n34183, ZN => n34170);
   U35051 : OAI22_X1 port map( A1 => n16968, A2 => n39546, B1 => n35443, B2 => 
                           n39540, ZN => n7229);
   U35052 : NOR2_X1 port map( A1 => n35444, A2 => n35445, ZN => n35443);
   U35053 : NAND4_X1 port map( A1 => n35446, A2 => n35447, A3 => n35448, A4 => 
                           n35449, ZN => n35445);
   U35054 : NAND4_X1 port map( A1 => n35454, A2 => n35455, A3 => n35456, A4 => 
                           n35457, ZN => n35444);
   U35055 : OAI22_X1 port map( A1 => n17031, A2 => n39798, B1 => n34188, B2 => 
                           n39792, ZN => n7292);
   U35056 : NOR2_X1 port map( A1 => n34189, A2 => n34190, ZN => n34188);
   U35057 : NAND4_X1 port map( A1 => n34191, A2 => n34192, A3 => n34193, A4 => 
                           n34194, ZN => n34190);
   U35058 : NAND4_X1 port map( A1 => n34199, A2 => n34200, A3 => n34201, A4 => 
                           n34202, ZN => n34189);
   U35059 : OAI22_X1 port map( A1 => n16967, A2 => n39546, B1 => n35462, B2 => 
                           n39540, ZN => n7228);
   U35060 : NOR2_X1 port map( A1 => n35463, A2 => n35464, ZN => n35462);
   U35061 : NAND4_X1 port map( A1 => n35465, A2 => n35466, A3 => n35467, A4 => 
                           n35468, ZN => n35464);
   U35062 : NAND4_X1 port map( A1 => n35473, A2 => n35474, A3 => n35475, A4 => 
                           n35476, ZN => n35463);
   U35063 : OAI22_X1 port map( A1 => n17030, A2 => n39798, B1 => n34207, B2 => 
                           n39792, ZN => n7291);
   U35064 : NOR2_X1 port map( A1 => n34208, A2 => n34209, ZN => n34207);
   U35065 : NAND4_X1 port map( A1 => n34210, A2 => n34211, A3 => n34212, A4 => 
                           n34213, ZN => n34209);
   U35066 : NAND4_X1 port map( A1 => n34218, A2 => n34219, A3 => n34220, A4 => 
                           n34221, ZN => n34208);
   U35067 : OAI22_X1 port map( A1 => n16966, A2 => n39546, B1 => n35481, B2 => 
                           n39540, ZN => n7227);
   U35068 : NOR2_X1 port map( A1 => n35482, A2 => n35483, ZN => n35481);
   U35069 : NAND4_X1 port map( A1 => n35484, A2 => n35485, A3 => n35486, A4 => 
                           n35487, ZN => n35483);
   U35070 : NAND4_X1 port map( A1 => n35492, A2 => n35493, A3 => n35494, A4 => 
                           n35495, ZN => n35482);
   U35071 : OAI22_X1 port map( A1 => n17029, A2 => n39798, B1 => n34226, B2 => 
                           n39791, ZN => n7290);
   U35072 : NOR2_X1 port map( A1 => n34227, A2 => n34228, ZN => n34226);
   U35073 : NAND4_X1 port map( A1 => n34229, A2 => n34230, A3 => n34231, A4 => 
                           n34232, ZN => n34228);
   U35074 : NAND4_X1 port map( A1 => n34237, A2 => n34238, A3 => n34239, A4 => 
                           n34240, ZN => n34227);
   U35075 : OAI22_X1 port map( A1 => n16965, A2 => n39546, B1 => n35500, B2 => 
                           n39539, ZN => n7226);
   U35076 : NOR2_X1 port map( A1 => n35501, A2 => n35502, ZN => n35500);
   U35077 : NAND4_X1 port map( A1 => n35503, A2 => n35504, A3 => n35505, A4 => 
                           n35506, ZN => n35502);
   U35078 : NAND4_X1 port map( A1 => n35511, A2 => n35512, A3 => n35513, A4 => 
                           n35514, ZN => n35501);
   U35079 : OAI22_X1 port map( A1 => n17028, A2 => n39797, B1 => n34245, B2 => 
                           n39791, ZN => n7289);
   U35080 : NOR2_X1 port map( A1 => n34246, A2 => n34247, ZN => n34245);
   U35081 : NAND4_X1 port map( A1 => n34248, A2 => n34249, A3 => n34250, A4 => 
                           n34251, ZN => n34247);
   U35082 : NAND4_X1 port map( A1 => n34256, A2 => n34257, A3 => n34258, A4 => 
                           n34259, ZN => n34246);
   U35083 : OAI22_X1 port map( A1 => n16964, A2 => n39545, B1 => n35519, B2 => 
                           n39539, ZN => n7225);
   U35084 : NOR2_X1 port map( A1 => n35520, A2 => n35521, ZN => n35519);
   U35085 : NAND4_X1 port map( A1 => n35522, A2 => n35523, A3 => n35524, A4 => 
                           n35525, ZN => n35521);
   U35086 : NAND4_X1 port map( A1 => n35530, A2 => n35531, A3 => n35532, A4 => 
                           n35533, ZN => n35520);
   U35087 : OAI22_X1 port map( A1 => n17027, A2 => n39797, B1 => n34264, B2 => 
                           n39791, ZN => n7288);
   U35088 : NOR2_X1 port map( A1 => n34265, A2 => n34266, ZN => n34264);
   U35089 : NAND4_X1 port map( A1 => n34267, A2 => n34268, A3 => n34269, A4 => 
                           n34270, ZN => n34266);
   U35090 : NAND4_X1 port map( A1 => n34275, A2 => n34276, A3 => n34277, A4 => 
                           n34278, ZN => n34265);
   U35091 : OAI22_X1 port map( A1 => n16963, A2 => n39545, B1 => n35538, B2 => 
                           n39539, ZN => n7224);
   U35092 : NOR2_X1 port map( A1 => n35539, A2 => n35540, ZN => n35538);
   U35093 : NAND4_X1 port map( A1 => n35541, A2 => n35542, A3 => n35543, A4 => 
                           n35544, ZN => n35540);
   U35094 : NAND4_X1 port map( A1 => n35549, A2 => n35550, A3 => n35551, A4 => 
                           n35552, ZN => n35539);
   U35095 : OAI22_X1 port map( A1 => n17026, A2 => n39797, B1 => n34283, B2 => 
                           n39791, ZN => n7287);
   U35096 : NOR2_X1 port map( A1 => n34284, A2 => n34285, ZN => n34283);
   U35097 : NAND4_X1 port map( A1 => n34286, A2 => n34287, A3 => n34288, A4 => 
                           n34289, ZN => n34285);
   U35098 : NAND4_X1 port map( A1 => n34294, A2 => n34295, A3 => n34296, A4 => 
                           n34297, ZN => n34284);
   U35099 : OAI22_X1 port map( A1 => n16962, A2 => n39545, B1 => n35557, B2 => 
                           n39539, ZN => n7223);
   U35100 : NOR2_X1 port map( A1 => n35558, A2 => n35559, ZN => n35557);
   U35101 : NAND4_X1 port map( A1 => n35560, A2 => n35561, A3 => n35562, A4 => 
                           n35563, ZN => n35559);
   U35102 : NAND4_X1 port map( A1 => n35568, A2 => n35569, A3 => n35570, A4 => 
                           n35571, ZN => n35558);
   U35103 : OAI22_X1 port map( A1 => n17025, A2 => n39797, B1 => n34302, B2 => 
                           n39791, ZN => n7286);
   U35104 : NOR2_X1 port map( A1 => n34303, A2 => n34304, ZN => n34302);
   U35105 : NAND4_X1 port map( A1 => n34305, A2 => n34306, A3 => n34307, A4 => 
                           n34308, ZN => n34304);
   U35106 : NAND4_X1 port map( A1 => n34313, A2 => n34314, A3 => n34315, A4 => 
                           n34316, ZN => n34303);
   U35107 : OAI22_X1 port map( A1 => n16961, A2 => n39545, B1 => n35576, B2 => 
                           n39539, ZN => n7222);
   U35108 : NOR2_X1 port map( A1 => n35577, A2 => n35578, ZN => n35576);
   U35109 : NAND4_X1 port map( A1 => n35579, A2 => n35580, A3 => n35581, A4 => 
                           n35582, ZN => n35578);
   U35110 : NAND4_X1 port map( A1 => n35587, A2 => n35588, A3 => n35589, A4 => 
                           n35590, ZN => n35577);
   U35111 : OAI22_X1 port map( A1 => n17024, A2 => n39797, B1 => n34321, B2 => 
                           n39791, ZN => n7285);
   U35112 : NOR2_X1 port map( A1 => n34322, A2 => n34323, ZN => n34321);
   U35113 : NAND4_X1 port map( A1 => n34324, A2 => n34325, A3 => n34326, A4 => 
                           n34327, ZN => n34323);
   U35114 : NAND4_X1 port map( A1 => n34332, A2 => n34333, A3 => n34334, A4 => 
                           n34335, ZN => n34322);
   U35115 : OAI22_X1 port map( A1 => n16960, A2 => n39545, B1 => n35595, B2 => 
                           n39539, ZN => n7221);
   U35116 : NOR2_X1 port map( A1 => n35596, A2 => n35597, ZN => n35595);
   U35117 : NAND4_X1 port map( A1 => n35598, A2 => n35599, A3 => n35600, A4 => 
                           n35601, ZN => n35597);
   U35118 : NAND4_X1 port map( A1 => n35606, A2 => n35607, A3 => n35608, A4 => 
                           n35609, ZN => n35596);
   U35119 : OAI22_X1 port map( A1 => n17023, A2 => n39797, B1 => n34340, B2 => 
                           n39791, ZN => n7284);
   U35120 : NOR2_X1 port map( A1 => n34341, A2 => n34342, ZN => n34340);
   U35121 : NAND4_X1 port map( A1 => n34343, A2 => n34344, A3 => n34345, A4 => 
                           n34346, ZN => n34342);
   U35122 : NAND4_X1 port map( A1 => n34351, A2 => n34352, A3 => n34353, A4 => 
                           n34354, ZN => n34341);
   U35123 : OAI22_X1 port map( A1 => n16959, A2 => n39545, B1 => n35614, B2 => 
                           n39539, ZN => n7220);
   U35124 : NOR2_X1 port map( A1 => n35615, A2 => n35616, ZN => n35614);
   U35125 : NAND4_X1 port map( A1 => n35617, A2 => n35618, A3 => n35619, A4 => 
                           n35620, ZN => n35616);
   U35126 : NAND4_X1 port map( A1 => n35625, A2 => n35626, A3 => n35627, A4 => 
                           n35628, ZN => n35615);
   U35127 : OAI22_X1 port map( A1 => n17022, A2 => n39797, B1 => n34359, B2 => 
                           n39791, ZN => n7283);
   U35128 : NOR2_X1 port map( A1 => n34360, A2 => n34361, ZN => n34359);
   U35129 : NAND4_X1 port map( A1 => n34362, A2 => n34363, A3 => n34364, A4 => 
                           n34365, ZN => n34361);
   U35130 : NAND4_X1 port map( A1 => n34370, A2 => n34371, A3 => n34372, A4 => 
                           n34373, ZN => n34360);
   U35131 : OAI22_X1 port map( A1 => n16958, A2 => n39545, B1 => n35633, B2 => 
                           n39539, ZN => n7219);
   U35132 : NOR2_X1 port map( A1 => n35634, A2 => n35635, ZN => n35633);
   U35133 : NAND4_X1 port map( A1 => n35636, A2 => n35637, A3 => n35638, A4 => 
                           n35639, ZN => n35635);
   U35134 : NAND4_X1 port map( A1 => n35644, A2 => n35645, A3 => n35646, A4 => 
                           n35647, ZN => n35634);
   U35135 : OAI22_X1 port map( A1 => n17021, A2 => n39797, B1 => n34378, B2 => 
                           n39791, ZN => n7282);
   U35136 : NOR2_X1 port map( A1 => n34379, A2 => n34380, ZN => n34378);
   U35137 : NAND4_X1 port map( A1 => n34381, A2 => n34382, A3 => n34383, A4 => 
                           n34384, ZN => n34380);
   U35138 : NAND4_X1 port map( A1 => n34389, A2 => n34390, A3 => n34391, A4 => 
                           n34392, ZN => n34379);
   U35139 : OAI22_X1 port map( A1 => n16957, A2 => n39545, B1 => n35652, B2 => 
                           n39539, ZN => n7218);
   U35140 : NOR2_X1 port map( A1 => n35653, A2 => n35654, ZN => n35652);
   U35141 : NAND4_X1 port map( A1 => n35655, A2 => n35656, A3 => n35657, A4 => 
                           n35658, ZN => n35654);
   U35142 : NAND4_X1 port map( A1 => n35663, A2 => n35664, A3 => n35665, A4 => 
                           n35666, ZN => n35653);
   U35143 : OAI22_X1 port map( A1 => n17020, A2 => n39797, B1 => n34397, B2 => 
                           n39791, ZN => n7281);
   U35144 : NOR2_X1 port map( A1 => n34398, A2 => n34399, ZN => n34397);
   U35145 : NAND4_X1 port map( A1 => n34400, A2 => n34401, A3 => n34402, A4 => 
                           n34403, ZN => n34399);
   U35146 : NAND4_X1 port map( A1 => n34408, A2 => n34409, A3 => n34410, A4 => 
                           n34411, ZN => n34398);
   U35147 : OAI22_X1 port map( A1 => n16956, A2 => n39545, B1 => n35671, B2 => 
                           n39539, ZN => n7217);
   U35148 : NOR2_X1 port map( A1 => n35672, A2 => n35673, ZN => n35671);
   U35149 : NAND4_X1 port map( A1 => n35674, A2 => n35675, A3 => n35676, A4 => 
                           n35677, ZN => n35673);
   U35150 : NAND4_X1 port map( A1 => n35682, A2 => n35683, A3 => n35684, A4 => 
                           n35685, ZN => n35672);
   U35151 : OAI22_X1 port map( A1 => n17019, A2 => n39797, B1 => n34416, B2 => 
                           n39791, ZN => n7280);
   U35152 : NOR2_X1 port map( A1 => n34417, A2 => n34418, ZN => n34416);
   U35153 : NAND4_X1 port map( A1 => n34419, A2 => n34420, A3 => n34421, A4 => 
                           n34422, ZN => n34418);
   U35154 : NAND4_X1 port map( A1 => n34427, A2 => n34428, A3 => n34429, A4 => 
                           n34430, ZN => n34417);
   U35155 : OAI22_X1 port map( A1 => n16955, A2 => n39545, B1 => n35690, B2 => 
                           n39539, ZN => n7216);
   U35156 : NOR2_X1 port map( A1 => n35691, A2 => n35692, ZN => n35690);
   U35157 : NAND4_X1 port map( A1 => n35693, A2 => n35694, A3 => n35695, A4 => 
                           n35696, ZN => n35692);
   U35158 : NAND4_X1 port map( A1 => n35701, A2 => n35702, A3 => n35703, A4 => 
                           n35704, ZN => n35691);
   U35159 : OAI22_X1 port map( A1 => n17018, A2 => n39797, B1 => n34435, B2 => 
                           n39791, ZN => n7279);
   U35160 : NOR2_X1 port map( A1 => n34436, A2 => n34437, ZN => n34435);
   U35161 : NAND4_X1 port map( A1 => n34438, A2 => n34439, A3 => n34440, A4 => 
                           n34441, ZN => n34437);
   U35162 : NAND4_X1 port map( A1 => n34446, A2 => n34447, A3 => n34448, A4 => 
                           n34449, ZN => n34436);
   U35163 : OAI22_X1 port map( A1 => n16954, A2 => n39545, B1 => n35709, B2 => 
                           n39539, ZN => n7215);
   U35164 : NOR2_X1 port map( A1 => n35710, A2 => n35711, ZN => n35709);
   U35165 : NAND4_X1 port map( A1 => n35712, A2 => n35713, A3 => n35714, A4 => 
                           n35715, ZN => n35711);
   U35166 : NAND4_X1 port map( A1 => n35720, A2 => n35721, A3 => n35722, A4 => 
                           n35723, ZN => n35710);
   U35167 : OAI22_X1 port map( A1 => n17017, A2 => n39797, B1 => n34454, B2 => 
                           n39790, ZN => n7278);
   U35168 : NOR2_X1 port map( A1 => n34455, A2 => n34456, ZN => n34454);
   U35169 : NAND4_X1 port map( A1 => n34457, A2 => n34458, A3 => n34459, A4 => 
                           n34460, ZN => n34456);
   U35170 : NAND4_X1 port map( A1 => n34465, A2 => n34466, A3 => n34467, A4 => 
                           n34468, ZN => n34455);
   U35171 : OAI22_X1 port map( A1 => n16953, A2 => n39545, B1 => n35728, B2 => 
                           n39538, ZN => n7214);
   U35172 : NOR2_X1 port map( A1 => n35729, A2 => n35730, ZN => n35728);
   U35173 : NAND4_X1 port map( A1 => n35731, A2 => n35732, A3 => n35733, A4 => 
                           n35734, ZN => n35730);
   U35174 : NAND4_X1 port map( A1 => n35739, A2 => n35740, A3 => n35741, A4 => 
                           n35742, ZN => n35729);
   U35175 : OAI22_X1 port map( A1 => n17016, A2 => n39796, B1 => n34473, B2 => 
                           n39790, ZN => n7277);
   U35176 : NOR2_X1 port map( A1 => n34474, A2 => n34475, ZN => n34473);
   U35177 : NAND4_X1 port map( A1 => n34476, A2 => n34477, A3 => n34478, A4 => 
                           n34479, ZN => n34475);
   U35178 : NAND4_X1 port map( A1 => n34484, A2 => n34485, A3 => n34486, A4 => 
                           n34487, ZN => n34474);
   U35179 : OAI22_X1 port map( A1 => n16952, A2 => n39544, B1 => n35747, B2 => 
                           n39538, ZN => n7213);
   U35180 : NOR2_X1 port map( A1 => n35748, A2 => n35749, ZN => n35747);
   U35181 : NAND4_X1 port map( A1 => n35750, A2 => n35751, A3 => n35752, A4 => 
                           n35753, ZN => n35749);
   U35182 : NAND4_X1 port map( A1 => n35758, A2 => n35759, A3 => n35760, A4 => 
                           n35761, ZN => n35748);
   U35183 : OAI22_X1 port map( A1 => n17015, A2 => n39796, B1 => n34492, B2 => 
                           n39790, ZN => n7276);
   U35184 : NOR2_X1 port map( A1 => n34493, A2 => n34494, ZN => n34492);
   U35185 : NAND4_X1 port map( A1 => n34495, A2 => n34496, A3 => n34497, A4 => 
                           n34498, ZN => n34494);
   U35186 : NAND4_X1 port map( A1 => n34503, A2 => n34504, A3 => n34505, A4 => 
                           n34506, ZN => n34493);
   U35187 : OAI22_X1 port map( A1 => n16951, A2 => n39544, B1 => n35766, B2 => 
                           n39538, ZN => n7212);
   U35188 : NOR2_X1 port map( A1 => n35767, A2 => n35768, ZN => n35766);
   U35189 : NAND4_X1 port map( A1 => n35769, A2 => n35770, A3 => n35771, A4 => 
                           n35772, ZN => n35768);
   U35190 : NAND4_X1 port map( A1 => n35777, A2 => n35778, A3 => n35779, A4 => 
                           n35780, ZN => n35767);
   U35191 : OAI22_X1 port map( A1 => n17014, A2 => n39796, B1 => n34511, B2 => 
                           n39790, ZN => n7275);
   U35192 : NOR2_X1 port map( A1 => n34512, A2 => n34513, ZN => n34511);
   U35193 : NAND4_X1 port map( A1 => n34514, A2 => n34515, A3 => n34516, A4 => 
                           n34517, ZN => n34513);
   U35194 : NAND4_X1 port map( A1 => n34522, A2 => n34523, A3 => n34524, A4 => 
                           n34525, ZN => n34512);
   U35195 : OAI22_X1 port map( A1 => n16950, A2 => n39544, B1 => n35785, B2 => 
                           n39538, ZN => n7211);
   U35196 : NOR2_X1 port map( A1 => n35786, A2 => n35787, ZN => n35785);
   U35197 : NAND4_X1 port map( A1 => n35788, A2 => n35789, A3 => n35790, A4 => 
                           n35791, ZN => n35787);
   U35198 : NAND4_X1 port map( A1 => n35796, A2 => n35797, A3 => n35798, A4 => 
                           n35799, ZN => n35786);
   U35199 : OAI22_X1 port map( A1 => n17013, A2 => n39796, B1 => n34530, B2 => 
                           n39790, ZN => n7274);
   U35200 : NOR2_X1 port map( A1 => n34531, A2 => n34532, ZN => n34530);
   U35201 : NAND4_X1 port map( A1 => n34533, A2 => n34534, A3 => n34535, A4 => 
                           n34536, ZN => n34532);
   U35202 : NAND4_X1 port map( A1 => n34541, A2 => n34542, A3 => n34543, A4 => 
                           n34544, ZN => n34531);
   U35203 : OAI22_X1 port map( A1 => n16949, A2 => n39544, B1 => n35804, B2 => 
                           n39538, ZN => n7210);
   U35204 : NOR2_X1 port map( A1 => n35805, A2 => n35806, ZN => n35804);
   U35205 : NAND4_X1 port map( A1 => n35807, A2 => n35808, A3 => n35809, A4 => 
                           n35810, ZN => n35806);
   U35206 : NAND4_X1 port map( A1 => n35815, A2 => n35816, A3 => n35817, A4 => 
                           n35818, ZN => n35805);
   U35207 : OAI22_X1 port map( A1 => n17012, A2 => n39796, B1 => n34549, B2 => 
                           n39790, ZN => n7273);
   U35208 : NOR2_X1 port map( A1 => n34550, A2 => n34551, ZN => n34549);
   U35209 : NAND4_X1 port map( A1 => n34552, A2 => n34553, A3 => n34554, A4 => 
                           n34555, ZN => n34551);
   U35210 : NAND4_X1 port map( A1 => n34560, A2 => n34561, A3 => n34562, A4 => 
                           n34563, ZN => n34550);
   U35211 : OAI22_X1 port map( A1 => n16948, A2 => n39544, B1 => n35823, B2 => 
                           n39538, ZN => n7209);
   U35212 : NOR2_X1 port map( A1 => n35824, A2 => n35825, ZN => n35823);
   U35213 : NAND4_X1 port map( A1 => n35826, A2 => n35827, A3 => n35828, A4 => 
                           n35829, ZN => n35825);
   U35214 : NAND4_X1 port map( A1 => n35834, A2 => n35835, A3 => n35836, A4 => 
                           n35837, ZN => n35824);
   U35215 : OAI22_X1 port map( A1 => n17011, A2 => n39796, B1 => n34568, B2 => 
                           n39790, ZN => n7272);
   U35216 : NOR2_X1 port map( A1 => n34569, A2 => n34570, ZN => n34568);
   U35217 : NAND4_X1 port map( A1 => n34571, A2 => n34572, A3 => n34573, A4 => 
                           n34574, ZN => n34570);
   U35218 : NAND4_X1 port map( A1 => n34579, A2 => n34580, A3 => n34581, A4 => 
                           n34582, ZN => n34569);
   U35219 : OAI22_X1 port map( A1 => n16947, A2 => n39544, B1 => n35842, B2 => 
                           n39538, ZN => n7208);
   U35220 : NOR2_X1 port map( A1 => n35843, A2 => n35844, ZN => n35842);
   U35221 : NAND4_X1 port map( A1 => n35845, A2 => n35846, A3 => n35847, A4 => 
                           n35848, ZN => n35844);
   U35222 : NAND4_X1 port map( A1 => n35853, A2 => n35854, A3 => n35855, A4 => 
                           n35856, ZN => n35843);
   U35223 : OAI22_X1 port map( A1 => n17010, A2 => n39796, B1 => n34587, B2 => 
                           n39790, ZN => n7271);
   U35224 : NOR2_X1 port map( A1 => n34588, A2 => n34589, ZN => n34587);
   U35225 : NAND4_X1 port map( A1 => n34590, A2 => n34591, A3 => n34592, A4 => 
                           n34593, ZN => n34589);
   U35226 : NAND4_X1 port map( A1 => n34598, A2 => n34599, A3 => n34600, A4 => 
                           n34601, ZN => n34588);
   U35227 : OAI22_X1 port map( A1 => n16946, A2 => n39544, B1 => n35861, B2 => 
                           n39538, ZN => n7207);
   U35228 : NOR2_X1 port map( A1 => n35862, A2 => n35863, ZN => n35861);
   U35229 : NAND4_X1 port map( A1 => n35864, A2 => n35865, A3 => n35866, A4 => 
                           n35867, ZN => n35863);
   U35230 : NAND4_X1 port map( A1 => n35872, A2 => n35873, A3 => n35874, A4 => 
                           n35875, ZN => n35862);
   U35231 : OAI22_X1 port map( A1 => n17009, A2 => n39796, B1 => n34606, B2 => 
                           n39790, ZN => n7270);
   U35232 : NOR2_X1 port map( A1 => n34607, A2 => n34608, ZN => n34606);
   U35233 : NAND4_X1 port map( A1 => n34609, A2 => n34610, A3 => n34611, A4 => 
                           n34612, ZN => n34608);
   U35234 : NAND4_X1 port map( A1 => n34617, A2 => n34618, A3 => n34619, A4 => 
                           n34620, ZN => n34607);
   U35235 : OAI22_X1 port map( A1 => n16945, A2 => n39544, B1 => n35880, B2 => 
                           n39538, ZN => n7206);
   U35236 : NOR2_X1 port map( A1 => n35881, A2 => n35882, ZN => n35880);
   U35237 : NAND4_X1 port map( A1 => n35883, A2 => n35884, A3 => n35885, A4 => 
                           n35886, ZN => n35882);
   U35238 : NAND4_X1 port map( A1 => n35891, A2 => n35892, A3 => n35893, A4 => 
                           n35894, ZN => n35881);
   U35239 : OAI22_X1 port map( A1 => n17008, A2 => n39796, B1 => n34625, B2 => 
                           n39790, ZN => n7269);
   U35240 : NOR2_X1 port map( A1 => n34626, A2 => n34627, ZN => n34625);
   U35241 : NAND4_X1 port map( A1 => n34628, A2 => n34629, A3 => n34630, A4 => 
                           n34631, ZN => n34627);
   U35242 : NAND4_X1 port map( A1 => n34636, A2 => n34637, A3 => n34638, A4 => 
                           n34639, ZN => n34626);
   U35243 : OAI22_X1 port map( A1 => n16944, A2 => n39544, B1 => n35899, B2 => 
                           n39538, ZN => n7205);
   U35244 : NOR2_X1 port map( A1 => n35900, A2 => n35901, ZN => n35899);
   U35245 : NAND4_X1 port map( A1 => n35902, A2 => n35903, A3 => n35904, A4 => 
                           n35905, ZN => n35901);
   U35246 : NAND4_X1 port map( A1 => n35910, A2 => n35911, A3 => n35912, A4 => 
                           n35913, ZN => n35900);
   U35247 : OAI22_X1 port map( A1 => n17007, A2 => n39796, B1 => n34644, B2 => 
                           n39790, ZN => n7268);
   U35248 : NOR2_X1 port map( A1 => n34645, A2 => n34646, ZN => n34644);
   U35249 : NAND4_X1 port map( A1 => n34647, A2 => n34648, A3 => n34649, A4 => 
                           n34650, ZN => n34646);
   U35250 : NAND4_X1 port map( A1 => n34655, A2 => n34656, A3 => n34657, A4 => 
                           n34658, ZN => n34645);
   U35251 : OAI22_X1 port map( A1 => n16943, A2 => n39544, B1 => n35918, B2 => 
                           n39538, ZN => n7204);
   U35252 : NOR2_X1 port map( A1 => n35919, A2 => n35920, ZN => n35918);
   U35253 : NAND4_X1 port map( A1 => n35921, A2 => n35922, A3 => n35923, A4 => 
                           n35924, ZN => n35920);
   U35254 : NAND4_X1 port map( A1 => n35929, A2 => n35930, A3 => n35931, A4 => 
                           n35932, ZN => n35919);
   U35255 : OAI22_X1 port map( A1 => n17006, A2 => n39796, B1 => n34663, B2 => 
                           n39790, ZN => n7267);
   U35256 : NOR2_X1 port map( A1 => n34664, A2 => n34665, ZN => n34663);
   U35257 : NAND4_X1 port map( A1 => n34666, A2 => n34667, A3 => n34668, A4 => 
                           n34669, ZN => n34665);
   U35258 : NAND4_X1 port map( A1 => n34685, A2 => n34686, A3 => n34687, A4 => 
                           n34688, ZN => n34664);
   U35259 : OAI22_X1 port map( A1 => n16942, A2 => n39544, B1 => n35937, B2 => 
                           n39538, ZN => n7203);
   U35260 : NOR2_X1 port map( A1 => n35938, A2 => n35939, ZN => n35937);
   U35261 : NAND4_X1 port map( A1 => n35940, A2 => n35941, A3 => n35942, A4 => 
                           n35943, ZN => n35939);
   U35262 : NAND4_X1 port map( A1 => n35959, A2 => n35960, A3 => n35961, A4 => 
                           n35962, ZN => n35938);
   U35263 : NOR2_X1 port map( A1 => n2699, A2 => n2710, ZN => n12791);
   U35264 : NOR2_X1 port map( A1 => n2695, A2 => n32167, ZN => U3_U194_Z_4);
   U35265 : NOR2_X1 port map( A1 => n2695, A2 => n32172, ZN => U3_U195_Z_4);
   U35266 : AND2_X1 port map( A1 => n33301, A2 => WR, ZN => n33330);
   U35267 : NOR2_X1 port map( A1 => n2698, A2 => n32167, ZN => U3_U194_Z_1);
   U35268 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n32253, A3 => n33208, ZN 
                           => r504_n3);
   U35269 : NOR2_X1 port map( A1 => n2698, A2 => n32172, ZN => U3_U195_Z_1);
   U35270 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n32253, A3 => n33207, ZN 
                           => r510_n3);
   U35271 : NOR2_X1 port map( A1 => n2697, A2 => n32167, ZN => U3_U194_Z_2);
   U35272 : NOR2_X1 port map( A1 => n2697, A2 => n32172, ZN => U3_U195_Z_2);
   U35273 : NOR2_X1 port map( A1 => n2698, A2 => n32162, ZN => U3_U193_Z_1);
   U35274 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n32253, A3 => n33209, ZN 
                           => r498_n1);
   U35275 : NAND2_X1 port map( A1 => n2696, A2 => n33208, ZN => U3_U194_Z_3);
   U35276 : NAND2_X1 port map( A1 => n2696, A2 => n33207, ZN => U3_U195_Z_3);
   U35277 : NOR2_X1 port map( A1 => n2697, A2 => n32162, ZN => U3_U193_Z_2);
   U35278 : NAND2_X1 port map( A1 => n2696, A2 => n33209, ZN => U3_U193_Z_3);
   U35279 : NOR3_X1 port map( A1 => n32075, A2 => RESET, A3 => n33227, ZN => 
                           n33223);
   U35280 : OAI222_X1 port map( A1 => n32240, A2 => n33211, B1 => n33215, B2 =>
                           n33213, C1 => n2683, C2 => n33212, ZN => n9902);
   U35281 : INV_X1 port map( A => n33215, ZN => n32240);
   U35282 : OAI22_X1 port map( A1 => n33250, A2 => i_2_port, B1 => n2707, B2 =>
                           n33251, ZN => n9891);
   U35283 : AOI211_X1 port map( C1 => n2709, C2 => n33249, A => n32077, B => 
                           n32076, ZN => n33251);
   U35284 : NAND4_X1 port map( A1 => n2699, A2 => n2698, A3 => n35979, A4 => 
                           n2697, ZN => n33218);
   U35285 : NOR2_X1 port map( A1 => n2695, A2 => N661, ZN => n35979);
   U35286 : XNOR2_X1 port map( A => n32244, B => n2695, ZN => n33215);
   U35287 : OAI21_X1 port map( B1 => n23853, B2 => n32081, A => n39297, ZN => 
                           n33233);
   U35288 : NAND4_X1 port map( A1 => n33238, A2 => n33239, A3 => n32238, A4 => 
                           n33240, ZN => n33227);
   U35289 : NOR4_X1 port map( A1 => n33241, A2 => n32083, A3 => n33242, A4 => 
                           n33243, ZN => n33240);
   U35290 : INV_X1 port map( A => n33244, ZN => n32238);
   U35291 : OAI211_X1 port map( C1 => n35974, C2 => n35975, A => ENABLE, B => 
                           CALL, ZN => n33232);
   U35292 : NOR4_X1 port map( A1 => n35976, A2 => n33218, A3 => n32259, A4 => 
                           n32261, ZN => n35975);
   U35293 : NOR4_X1 port map( A1 => n35977, A2 => n35978, A3 => n33242, A4 => 
                           n33243, ZN => n35974);
   U35294 : NAND4_X1 port map( A1 => n2695, A2 => n2683, A3 => n33246, A4 => 
                           n2699, ZN => n33216);
   U35295 : AND2_X1 port map( A1 => n2696, A2 => n2697, ZN => n33246);
   U35296 : XNOR2_X1 port map( A => n32322, B => n2695, ZN => n33238);
   U35297 : OAI211_X1 port map( C1 => N659, C2 => n33216, A => RETRN, B => 
                           n33217, ZN => n33213);
   U35298 : AND2_X1 port map( A1 => n41370, A2 => n33212, ZN => n33217);
   U35299 : OAI22_X1 port map( A1 => n33220, A2 => n32323, B1 => n27870, B2 => 
                           n33221, ZN => n9901);
   U35300 : AOI221_X1 port map( B1 => n33223, B2 => n27872, C1 => n33222, C2 =>
                           n32322, A => n32075, ZN => n33220);
   U35301 : AOI22_X1 port map( A1 => n33222, A2 => n27872, B1 => n33223, B2 => 
                           n32322, ZN => n33221);
   U35302 : OAI22_X1 port map( A1 => n2707, A2 => n33250, B1 => n2706, B2 => 
                           n37252, ZN => n25394);
   U35303 : NOR2_X1 port map( A1 => n33249, A2 => n32077, ZN => n37252);
   U35304 : OR4_X1 port map( A1 => n2706, A2 => n2707, A3 => n2709, A4 => n2710
                           , ZN => n33237);
   U35305 : OAI21_X1 port map( B1 => n2695, B2 => n33212, A => n33214, ZN => 
                           n9903);
   U35306 : NAND2_X1 port map( A1 => n33247, A2 => n33248, ZN => n9892);
   U35307 : OAI21_X1 port map( B1 => n32076, B2 => n32077, A => i_1_port, ZN =>
                           n33247);
   U35308 : OAI21_X1 port map( B1 => n23853, B2 => n33235, A => n33236, ZN => 
                           n9893);
   U35309 : OAI211_X1 port map( C1 => n23853, C2 => n33237, A => n33235, B => 
                           n41368, ZN => n33236);
   U35310 : OAI22_X1 port map( A1 => n23853, A2 => n32081, B1 => n33231, B2 => 
                           n33230, ZN => n33235);
   U35311 : OAI21_X1 port map( B1 => n2700, B2 => n39296, A => n35973, ZN => 
                           n7202);
   U35312 : OAI221_X1 port map( B1 => n32080, B2 => n39294, C1 => n2700, C2 => 
                           n33237, A => n41364, ZN => n35973);
   U35313 : INV_X1 port map( A => n33232, ZN => n32080);
   U35314 : NAND2_X1 port map( A1 => n2710, A2 => n33249, ZN => n33234);
   U35315 : INV_X1 port map( A => n35972, ZN => n39297);
   U35316 : OAI21_X1 port map( B1 => n2700, B2 => n33231, A => n41370, ZN => 
                           n35972);
   U35317 : OAI21_X1 port map( B1 => n2710, B2 => n33233, A => n33234, ZN => 
                           n9895);
   U35318 : AND4_X1 port map( A1 => n33228, A2 => n33227, A3 => n33225, A4 => 
                           n41364, ZN => n33222);
   U35319 : NAND4_X1 port map( A1 => n27872, A2 => n27871, A3 => n33229, A4 => 
                           n27874, ZN => n33228);
   U35320 : NOR2_X1 port map( A1 => n38789, A2 => n38790, ZN => n33229);
   U35321 : NOR2_X1 port map( A1 => n2699, A2 => n33210, ZN => n9907);
   U35322 : NOR2_X1 port map( A1 => n2698, A2 => n33210, ZN => n9906);
   U35323 : NOR2_X1 port map( A1 => n2697, A2 => n33210, ZN => n9905);
   U35324 : NOR2_X1 port map( A1 => n2696, A2 => n33210, ZN => n9904);
   U35325 : NOR2_X1 port map( A1 => n27871, A2 => n33224, ZN => n9900);
   U35326 : NOR2_X1 port map( A1 => n27874, A2 => n33224, ZN => n9898);
   U35327 : NOR2_X1 port map( A1 => n32082, A2 => RESET, ZN => n33230);
   U35328 : INV_X1 port map( A => n33227, ZN => n32082);
   U35329 : OAI21_X1 port map( B1 => n33231, B2 => n32148, A => n41370, ZN => 
                           n33424);
   U35330 : INV_X1 port map( A => RD1, ZN => n32148);
   U35331 : OAI21_X1 port map( B1 => n33231, B2 => n32149, A => n41370, ZN => 
                           n34698);
   U35332 : INV_X1 port map( A => RD2, ZN => n32149);
   U35333 : NOR2_X1 port map( A1 => ENABLE, A2 => RESET, ZN => n33231);
   U35334 : NAND2_X1 port map( A1 => n41370, A2 => n33219, ZN => n33212);
   U35335 : OAI21_X1 port map( B1 => CALL, B2 => RETRN, A => ENABLE, ZN => 
                           n33219);
   U35336 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n33208
                           );
   U35337 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n33207
                           );
   U35338 : NAND2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n33209);
   U35339 : INV_X1 port map( A => RESET, ZN => n32079);
   U35340 : INV_X1 port map( A => ENABLE, ZN => n32081);
   U35341 : INV_X1 port map( A => RETRN, ZN => n32083);
   U35342 : AND2_X1 port map( A1 => WR, A2 => n41370, ZN => n33300);
   U35343 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n33299);
   U35344 : INV_X1 port map( A => BUSin(23), ZN => n32124);
   U35345 : INV_X1 port map( A => DATAIN(23), ZN => n32214);
   U35346 : INV_X1 port map( A => BUSin(24), ZN => n32123);
   U35347 : INV_X1 port map( A => DATAIN(24), ZN => n32213);
   U35348 : INV_X1 port map( A => BUSin(25), ZN => n32122);
   U35349 : INV_X1 port map( A => DATAIN(25), ZN => n32212);
   U35350 : INV_X1 port map( A => BUSin(26), ZN => n32121);
   U35351 : INV_X1 port map( A => DATAIN(26), ZN => n32211);
   U35352 : INV_X1 port map( A => BUSin(27), ZN => n32120);
   U35353 : INV_X1 port map( A => DATAIN(27), ZN => n32210);
   U35354 : INV_X1 port map( A => BUSin(28), ZN => n32119);
   U35355 : INV_X1 port map( A => DATAIN(28), ZN => n32209);
   U35356 : INV_X1 port map( A => BUSin(29), ZN => n32118);
   U35357 : INV_X1 port map( A => DATAIN(29), ZN => n32208);
   U35358 : INV_X1 port map( A => BUSin(30), ZN => n32117);
   U35359 : INV_X1 port map( A => DATAIN(30), ZN => n32207);
   U35360 : INV_X1 port map( A => BUSin(31), ZN => n32116);
   U35361 : INV_X1 port map( A => DATAIN(31), ZN => n32206);
   U35362 : INV_X1 port map( A => BUSin(32), ZN => n32115);
   U35363 : INV_X1 port map( A => DATAIN(32), ZN => n32205);
   U35364 : INV_X1 port map( A => BUSin(33), ZN => n32114);
   U35365 : INV_X1 port map( A => DATAIN(33), ZN => n32204);
   U35366 : INV_X1 port map( A => BUSin(34), ZN => n32113);
   U35367 : INV_X1 port map( A => DATAIN(34), ZN => n32203);
   U35368 : INV_X1 port map( A => BUSin(35), ZN => n32112);
   U35369 : INV_X1 port map( A => DATAIN(35), ZN => n32202);
   U35370 : INV_X1 port map( A => BUSin(36), ZN => n32111);
   U35371 : INV_X1 port map( A => DATAIN(36), ZN => n32201);
   U35372 : INV_X1 port map( A => BUSin(37), ZN => n32110);
   U35373 : INV_X1 port map( A => DATAIN(37), ZN => n32200);
   U35374 : INV_X1 port map( A => BUSin(38), ZN => n32109);
   U35375 : INV_X1 port map( A => DATAIN(38), ZN => n32199);
   U35376 : INV_X1 port map( A => BUSin(39), ZN => n32108);
   U35377 : INV_X1 port map( A => DATAIN(39), ZN => n32198);
   U35378 : INV_X1 port map( A => BUSin(40), ZN => n32107);
   U35379 : INV_X1 port map( A => DATAIN(40), ZN => n32197);
   U35380 : INV_X1 port map( A => BUSin(41), ZN => n32106);
   U35381 : INV_X1 port map( A => DATAIN(41), ZN => n32196);
   U35382 : INV_X1 port map( A => BUSin(42), ZN => n32105);
   U35383 : INV_X1 port map( A => DATAIN(42), ZN => n32195);
   U35384 : INV_X1 port map( A => BUSin(43), ZN => n32104);
   U35385 : INV_X1 port map( A => DATAIN(43), ZN => n32194);
   U35386 : INV_X1 port map( A => BUSin(44), ZN => n32103);
   U35387 : INV_X1 port map( A => DATAIN(44), ZN => n32193);
   U35388 : INV_X1 port map( A => BUSin(45), ZN => n32102);
   U35389 : INV_X1 port map( A => DATAIN(45), ZN => n32192);
   U35390 : INV_X1 port map( A => BUSin(46), ZN => n32101);
   U35391 : INV_X1 port map( A => DATAIN(46), ZN => n32191);
   U35392 : INV_X1 port map( A => BUSin(47), ZN => n32100);
   U35393 : INV_X1 port map( A => DATAIN(47), ZN => n32190);
   U35394 : INV_X1 port map( A => BUSin(48), ZN => n32099);
   U35395 : INV_X1 port map( A => DATAIN(48), ZN => n32189);
   U35396 : INV_X1 port map( A => BUSin(49), ZN => n32098);
   U35397 : INV_X1 port map( A => DATAIN(49), ZN => n32188);
   U35398 : INV_X1 port map( A => BUSin(50), ZN => n32097);
   U35399 : INV_X1 port map( A => DATAIN(50), ZN => n32187);
   U35400 : INV_X1 port map( A => BUSin(51), ZN => n32096);
   U35401 : INV_X1 port map( A => DATAIN(51), ZN => n32186);
   U35402 : INV_X1 port map( A => BUSin(52), ZN => n32095);
   U35403 : INV_X1 port map( A => DATAIN(52), ZN => n32185);
   U35404 : INV_X1 port map( A => BUSin(53), ZN => n32094);
   U35405 : INV_X1 port map( A => DATAIN(53), ZN => n32184);
   U35406 : INV_X1 port map( A => BUSin(54), ZN => n32093);
   U35407 : INV_X1 port map( A => DATAIN(54), ZN => n32183);
   U35408 : INV_X1 port map( A => BUSin(55), ZN => n32092);
   U35409 : INV_X1 port map( A => DATAIN(55), ZN => n32182);
   U35410 : INV_X1 port map( A => BUSin(56), ZN => n32091);
   U35411 : INV_X1 port map( A => DATAIN(56), ZN => n32181);
   U35412 : INV_X1 port map( A => BUSin(57), ZN => n32090);
   U35413 : INV_X1 port map( A => DATAIN(57), ZN => n32180);
   U35414 : INV_X1 port map( A => BUSin(58), ZN => n32089);
   U35415 : INV_X1 port map( A => DATAIN(58), ZN => n32179);
   U35416 : INV_X1 port map( A => BUSin(59), ZN => n32088);
   U35417 : INV_X1 port map( A => DATAIN(59), ZN => n32178);
   U35418 : INV_X1 port map( A => BUSin(60), ZN => n32087);
   U35419 : INV_X1 port map( A => DATAIN(60), ZN => n32177);
   U35420 : INV_X1 port map( A => BUSin(61), ZN => n32086);
   U35421 : INV_X1 port map( A => DATAIN(61), ZN => n32176);
   U35422 : INV_X1 port map( A => BUSin(62), ZN => n32085);
   U35423 : INV_X1 port map( A => DATAIN(62), ZN => n32175);
   U35424 : INV_X1 port map( A => BUSin(63), ZN => n32084);
   U35425 : INV_X1 port map( A => DATAIN(63), ZN => n32174);
   U35426 : INV_X1 port map( A => BUSin(0), ZN => n32147);
   U35427 : INV_X1 port map( A => DATAIN(0), ZN => n32237);
   U35428 : INV_X1 port map( A => BUSin(1), ZN => n32146);
   U35429 : INV_X1 port map( A => DATAIN(1), ZN => n32236);
   U35430 : INV_X1 port map( A => BUSin(2), ZN => n32145);
   U35431 : INV_X1 port map( A => DATAIN(2), ZN => n32235);
   U35432 : INV_X1 port map( A => BUSin(3), ZN => n32144);
   U35433 : INV_X1 port map( A => DATAIN(3), ZN => n32234);
   U35434 : INV_X1 port map( A => BUSin(4), ZN => n32143);
   U35435 : INV_X1 port map( A => DATAIN(4), ZN => n32233);
   U35436 : INV_X1 port map( A => BUSin(5), ZN => n32142);
   U35437 : INV_X1 port map( A => DATAIN(5), ZN => n32232);
   U35438 : INV_X1 port map( A => BUSin(6), ZN => n32141);
   U35439 : INV_X1 port map( A => DATAIN(6), ZN => n32231);
   U35440 : INV_X1 port map( A => BUSin(7), ZN => n32140);
   U35441 : INV_X1 port map( A => DATAIN(7), ZN => n32230);
   U35442 : INV_X1 port map( A => BUSin(8), ZN => n32139);
   U35443 : INV_X1 port map( A => DATAIN(8), ZN => n32229);
   U35444 : INV_X1 port map( A => BUSin(9), ZN => n32138);
   U35445 : INV_X1 port map( A => DATAIN(9), ZN => n32228);
   U35446 : INV_X1 port map( A => BUSin(10), ZN => n32137);
   U35447 : INV_X1 port map( A => DATAIN(10), ZN => n32227);
   U35448 : INV_X1 port map( A => BUSin(11), ZN => n32136);
   U35449 : INV_X1 port map( A => DATAIN(11), ZN => n32226);
   U35450 : INV_X1 port map( A => BUSin(12), ZN => n32135);
   U35451 : INV_X1 port map( A => DATAIN(12), ZN => n32225);
   U35452 : INV_X1 port map( A => BUSin(13), ZN => n32134);
   U35453 : INV_X1 port map( A => DATAIN(13), ZN => n32224);
   U35454 : INV_X1 port map( A => BUSin(14), ZN => n32133);
   U35455 : INV_X1 port map( A => DATAIN(14), ZN => n32223);
   U35456 : INV_X1 port map( A => BUSin(15), ZN => n32132);
   U35457 : INV_X1 port map( A => DATAIN(15), ZN => n32222);
   U35458 : INV_X1 port map( A => BUSin(16), ZN => n32131);
   U35459 : INV_X1 port map( A => DATAIN(16), ZN => n32221);
   U35460 : INV_X1 port map( A => BUSin(17), ZN => n32130);
   U35461 : INV_X1 port map( A => DATAIN(17), ZN => n32220);
   U35462 : INV_X1 port map( A => BUSin(18), ZN => n32129);
   U35463 : INV_X1 port map( A => DATAIN(18), ZN => n32219);
   U35464 : INV_X1 port map( A => BUSin(19), ZN => n32128);
   U35465 : INV_X1 port map( A => DATAIN(19), ZN => n32218);
   U35466 : INV_X1 port map( A => BUSin(20), ZN => n32127);
   U35467 : INV_X1 port map( A => DATAIN(20), ZN => n32217);
   U35468 : INV_X1 port map( A => BUSin(21), ZN => n32126);
   U35469 : INV_X1 port map( A => DATAIN(21), ZN => n32216);
   U35470 : INV_X1 port map( A => BUSin(22), ZN => n32125);
   U35471 : INV_X1 port map( A => DATAIN(22), ZN => n32215);
   U35472 : CLKBUF_X1 port map( A => n36039, Z => n39053);
   U35473 : CLKBUF_X1 port map( A => n36038, Z => n39059);
   U35474 : CLKBUF_X1 port map( A => n36037, Z => n39065);
   U35475 : CLKBUF_X1 port map( A => n36035, Z => n39071);
   U35476 : CLKBUF_X1 port map( A => n36034, Z => n39077);
   U35477 : CLKBUF_X1 port map( A => n36033, Z => n39083);
   U35478 : CLKBUF_X1 port map( A => n36032, Z => n39089);
   U35479 : CLKBUF_X1 port map( A => n36031, Z => n39095);
   U35480 : CLKBUF_X1 port map( A => n36029, Z => n39101);
   U35481 : CLKBUF_X1 port map( A => n36028, Z => n39107);
   U35482 : CLKBUF_X1 port map( A => n36027, Z => n39113);
   U35483 : CLKBUF_X1 port map( A => n36026, Z => n39119);
   U35484 : CLKBUF_X1 port map( A => n36025, Z => n39125);
   U35485 : CLKBUF_X1 port map( A => n36023, Z => n39131);
   U35486 : CLKBUF_X1 port map( A => n36022, Z => n39137);
   U35487 : CLKBUF_X1 port map( A => n36021, Z => n39143);
   U35488 : CLKBUF_X1 port map( A => n36020, Z => n39149);
   U35489 : CLKBUF_X1 port map( A => n36019, Z => n39155);
   U35490 : CLKBUF_X1 port map( A => n36017, Z => n39161);
   U35491 : CLKBUF_X1 port map( A => n36016, Z => n39167);
   U35492 : CLKBUF_X1 port map( A => n36011, Z => n39173);
   U35493 : CLKBUF_X1 port map( A => n36010, Z => n39179);
   U35494 : CLKBUF_X1 port map( A => n36009, Z => n39185);
   U35495 : CLKBUF_X1 port map( A => n36007, Z => n39191);
   U35496 : CLKBUF_X1 port map( A => n36006, Z => n39197);
   U35497 : CLKBUF_X1 port map( A => n36005, Z => n39203);
   U35498 : CLKBUF_X1 port map( A => n36004, Z => n39209);
   U35499 : CLKBUF_X1 port map( A => n36003, Z => n39215);
   U35500 : CLKBUF_X1 port map( A => n36001, Z => n39221);
   U35501 : CLKBUF_X1 port map( A => n36000, Z => n39227);
   U35502 : CLKBUF_X1 port map( A => n35999, Z => n39233);
   U35503 : CLKBUF_X1 port map( A => n35998, Z => n39239);
   U35504 : CLKBUF_X1 port map( A => n35997, Z => n39245);
   U35505 : CLKBUF_X1 port map( A => n35995, Z => n39251);
   U35506 : CLKBUF_X1 port map( A => n35994, Z => n39257);
   U35507 : CLKBUF_X1 port map( A => n35993, Z => n39263);
   U35508 : CLKBUF_X1 port map( A => n35992, Z => n39269);
   U35509 : CLKBUF_X1 port map( A => n35991, Z => n39275);
   U35510 : CLKBUF_X1 port map( A => n35989, Z => n39281);
   U35511 : CLKBUF_X1 port map( A => n35988, Z => n39287);
   U35512 : CLKBUF_X1 port map( A => n35981, Z => n39293);
   U35513 : CLKBUF_X1 port map( A => n34758, Z => n39303);
   U35514 : CLKBUF_X1 port map( A => n34757, Z => n39309);
   U35515 : CLKBUF_X1 port map( A => n34756, Z => n39315);
   U35516 : CLKBUF_X1 port map( A => n34754, Z => n39321);
   U35517 : CLKBUF_X1 port map( A => n34753, Z => n39327);
   U35518 : CLKBUF_X1 port map( A => n34752, Z => n39333);
   U35519 : CLKBUF_X1 port map( A => n34751, Z => n39339);
   U35520 : CLKBUF_X1 port map( A => n34750, Z => n39345);
   U35521 : CLKBUF_X1 port map( A => n34748, Z => n39351);
   U35522 : CLKBUF_X1 port map( A => n34747, Z => n39357);
   U35523 : CLKBUF_X1 port map( A => n34746, Z => n39363);
   U35524 : CLKBUF_X1 port map( A => n34745, Z => n39369);
   U35525 : CLKBUF_X1 port map( A => n34744, Z => n39375);
   U35526 : CLKBUF_X1 port map( A => n34742, Z => n39381);
   U35527 : CLKBUF_X1 port map( A => n34741, Z => n39387);
   U35528 : CLKBUF_X1 port map( A => n34740, Z => n39393);
   U35529 : CLKBUF_X1 port map( A => n34739, Z => n39399);
   U35530 : CLKBUF_X1 port map( A => n34738, Z => n39405);
   U35531 : CLKBUF_X1 port map( A => n34736, Z => n39411);
   U35532 : CLKBUF_X1 port map( A => n34735, Z => n39417);
   U35533 : CLKBUF_X1 port map( A => n34730, Z => n39423);
   U35534 : CLKBUF_X1 port map( A => n34729, Z => n39429);
   U35535 : CLKBUF_X1 port map( A => n34728, Z => n39435);
   U35536 : CLKBUF_X1 port map( A => n34726, Z => n39441);
   U35537 : CLKBUF_X1 port map( A => n34725, Z => n39447);
   U35538 : CLKBUF_X1 port map( A => n34724, Z => n39453);
   U35539 : CLKBUF_X1 port map( A => n34723, Z => n39459);
   U35540 : CLKBUF_X1 port map( A => n34722, Z => n39465);
   U35541 : CLKBUF_X1 port map( A => n34720, Z => n39471);
   U35542 : CLKBUF_X1 port map( A => n34719, Z => n39477);
   U35543 : CLKBUF_X1 port map( A => n34718, Z => n39483);
   U35544 : CLKBUF_X1 port map( A => n34717, Z => n39489);
   U35545 : CLKBUF_X1 port map( A => n34716, Z => n39495);
   U35546 : CLKBUF_X1 port map( A => n34714, Z => n39501);
   U35547 : CLKBUF_X1 port map( A => n34713, Z => n39507);
   U35548 : CLKBUF_X1 port map( A => n34712, Z => n39513);
   U35549 : CLKBUF_X1 port map( A => n34711, Z => n39519);
   U35550 : CLKBUF_X1 port map( A => n34710, Z => n39525);
   U35551 : CLKBUF_X1 port map( A => n34708, Z => n39531);
   U35552 : CLKBUF_X1 port map( A => n34707, Z => n39537);
   U35553 : CLKBUF_X1 port map( A => n34700, Z => n39543);
   U35554 : CLKBUF_X1 port map( A => n34698, Z => n39549);
   U35555 : CLKBUF_X1 port map( A => n33484, Z => n39555);
   U35556 : CLKBUF_X1 port map( A => n33483, Z => n39561);
   U35557 : CLKBUF_X1 port map( A => n33482, Z => n39567);
   U35558 : CLKBUF_X1 port map( A => n33480, Z => n39573);
   U35559 : CLKBUF_X1 port map( A => n33479, Z => n39579);
   U35560 : CLKBUF_X1 port map( A => n33478, Z => n39585);
   U35561 : CLKBUF_X1 port map( A => n33477, Z => n39591);
   U35562 : CLKBUF_X1 port map( A => n33476, Z => n39597);
   U35563 : CLKBUF_X1 port map( A => n33474, Z => n39603);
   U35564 : CLKBUF_X1 port map( A => n33473, Z => n39609);
   U35565 : CLKBUF_X1 port map( A => n33472, Z => n39615);
   U35566 : CLKBUF_X1 port map( A => n33471, Z => n39621);
   U35567 : CLKBUF_X1 port map( A => n33470, Z => n39627);
   U35568 : CLKBUF_X1 port map( A => n33468, Z => n39633);
   U35569 : CLKBUF_X1 port map( A => n33467, Z => n39639);
   U35570 : CLKBUF_X1 port map( A => n33466, Z => n39645);
   U35571 : CLKBUF_X1 port map( A => n33465, Z => n39651);
   U35572 : CLKBUF_X1 port map( A => n33464, Z => n39657);
   U35573 : CLKBUF_X1 port map( A => n33462, Z => n39663);
   U35574 : CLKBUF_X1 port map( A => n33461, Z => n39669);
   U35575 : CLKBUF_X1 port map( A => n33456, Z => n39675);
   U35576 : CLKBUF_X1 port map( A => n33455, Z => n39681);
   U35577 : CLKBUF_X1 port map( A => n33454, Z => n39687);
   U35578 : CLKBUF_X1 port map( A => n33452, Z => n39693);
   U35579 : CLKBUF_X1 port map( A => n33451, Z => n39699);
   U35580 : CLKBUF_X1 port map( A => n33450, Z => n39705);
   U35581 : CLKBUF_X1 port map( A => n33449, Z => n39711);
   U35582 : CLKBUF_X1 port map( A => n33448, Z => n39717);
   U35583 : CLKBUF_X1 port map( A => n33446, Z => n39723);
   U35584 : CLKBUF_X1 port map( A => n33445, Z => n39729);
   U35585 : CLKBUF_X1 port map( A => n33444, Z => n39735);
   U35586 : CLKBUF_X1 port map( A => n33443, Z => n39741);
   U35587 : CLKBUF_X1 port map( A => n33442, Z => n39747);
   U35588 : CLKBUF_X1 port map( A => n33440, Z => n39753);
   U35589 : CLKBUF_X1 port map( A => n33439, Z => n39759);
   U35590 : CLKBUF_X1 port map( A => n33438, Z => n39765);
   U35591 : CLKBUF_X1 port map( A => n33437, Z => n39771);
   U35592 : CLKBUF_X1 port map( A => n33436, Z => n39777);
   U35593 : CLKBUF_X1 port map( A => n33434, Z => n39783);
   U35594 : CLKBUF_X1 port map( A => n33433, Z => n39789);
   U35595 : CLKBUF_X1 port map( A => n33426, Z => n39795);
   U35596 : CLKBUF_X1 port map( A => n33424, Z => n39801);
   U35597 : CLKBUF_X1 port map( A => n39807, Z => n39813);
   U35598 : CLKBUF_X1 port map( A => n39814, Z => n39820);
   U35599 : CLKBUF_X1 port map( A => n33417, Z => n39826);
   U35600 : CLKBUF_X1 port map( A => n39827, Z => n39833);
   U35601 : CLKBUF_X1 port map( A => n39834, Z => n39840);
   U35602 : CLKBUF_X1 port map( A => n33414, Z => n39846);
   U35603 : CLKBUF_X1 port map( A => n39847, Z => n39853);
   U35604 : CLKBUF_X1 port map( A => n39854, Z => n39860);
   U35605 : CLKBUF_X1 port map( A => n33411, Z => n39866);
   U35606 : CLKBUF_X1 port map( A => n39867, Z => n39873);
   U35607 : CLKBUF_X1 port map( A => n39874, Z => n39880);
   U35608 : CLKBUF_X1 port map( A => n33408, Z => n39886);
   U35609 : CLKBUF_X1 port map( A => n39887, Z => n39893);
   U35610 : CLKBUF_X1 port map( A => n39894, Z => n39900);
   U35611 : CLKBUF_X1 port map( A => n39906, Z => n39912);
   U35612 : CLKBUF_X1 port map( A => n39913, Z => n39919);
   U35613 : CLKBUF_X1 port map( A => n39925, Z => n39931);
   U35614 : CLKBUF_X1 port map( A => n39932, Z => n39938);
   U35615 : CLKBUF_X1 port map( A => n33393, Z => n39944);
   U35616 : CLKBUF_X1 port map( A => n39945, Z => n39951);
   U35617 : CLKBUF_X1 port map( A => n39952, Z => n39958);
   U35618 : CLKBUF_X1 port map( A => n33390, Z => n39964);
   U35619 : CLKBUF_X1 port map( A => n39965, Z => n39971);
   U35620 : CLKBUF_X1 port map( A => n39972, Z => n39978);
   U35621 : CLKBUF_X1 port map( A => n33387, Z => n39984);
   U35622 : CLKBUF_X1 port map( A => n39985, Z => n39991);
   U35623 : CLKBUF_X1 port map( A => n39992, Z => n39998);
   U35624 : CLKBUF_X1 port map( A => n40004, Z => n40010);
   U35625 : CLKBUF_X1 port map( A => n40011, Z => n40017);
   U35626 : CLKBUF_X1 port map( A => n40023, Z => n40029);
   U35627 : CLKBUF_X1 port map( A => n40030, Z => n40036);
   U35628 : CLKBUF_X1 port map( A => n33378, Z => n40042);
   U35629 : CLKBUF_X1 port map( A => n40043, Z => n40049);
   U35630 : CLKBUF_X1 port map( A => n40050, Z => n40056);
   U35631 : CLKBUF_X1 port map( A => n33375, Z => n40062);
   U35632 : CLKBUF_X1 port map( A => n40063, Z => n40069);
   U35633 : CLKBUF_X1 port map( A => n40070, Z => n40076);
   U35634 : CLKBUF_X1 port map( A => n33372, Z => n40082);
   U35635 : CLKBUF_X1 port map( A => n40083, Z => n40089);
   U35636 : CLKBUF_X1 port map( A => n40090, Z => n40096);
   U35637 : CLKBUF_X1 port map( A => n40102, Z => n40108);
   U35638 : CLKBUF_X1 port map( A => n40109, Z => n40115);
   U35639 : CLKBUF_X1 port map( A => n33361, Z => n40121);
   U35640 : CLKBUF_X1 port map( A => n40122, Z => n40128);
   U35641 : CLKBUF_X1 port map( A => n40129, Z => n40135);
   U35642 : CLKBUF_X1 port map( A => n33358, Z => n40141);
   U35643 : CLKBUF_X1 port map( A => n40142, Z => n40148);
   U35644 : CLKBUF_X1 port map( A => n40149, Z => n40155);
   U35645 : CLKBUF_X1 port map( A => n33355, Z => n40161);
   U35646 : CLKBUF_X1 port map( A => n40162, Z => n40168);
   U35647 : CLKBUF_X1 port map( A => n40169, Z => n40175);
   U35648 : CLKBUF_X1 port map( A => n33352, Z => n40181);
   U35649 : CLKBUF_X1 port map( A => n40182, Z => n40188);
   U35650 : CLKBUF_X1 port map( A => n40189, Z => n40195);
   U35651 : CLKBUF_X1 port map( A => n33349, Z => n40201);
   U35652 : CLKBUF_X1 port map( A => n40202, Z => n40208);
   U35653 : CLKBUF_X1 port map( A => n40209, Z => n40215);
   U35654 : CLKBUF_X1 port map( A => n33346, Z => n40221);
   U35655 : CLKBUF_X1 port map( A => n40222, Z => n40228);
   U35656 : CLKBUF_X1 port map( A => n40229, Z => n40235);
   U35657 : CLKBUF_X1 port map( A => n33343, Z => n40241);
   U35658 : CLKBUF_X1 port map( A => n40242, Z => n40248);
   U35659 : CLKBUF_X1 port map( A => n40249, Z => n40255);
   U35660 : CLKBUF_X1 port map( A => n33336, Z => n40261);
   U35661 : CLKBUF_X1 port map( A => n40262, Z => n40268);
   U35662 : CLKBUF_X1 port map( A => n40269, Z => n40275);
   U35663 : CLKBUF_X1 port map( A => n33329, Z => n40281);
   U35664 : CLKBUF_X1 port map( A => n40282, Z => n40288);
   U35665 : CLKBUF_X1 port map( A => n40289, Z => n40295);
   U35666 : CLKBUF_X1 port map( A => n33326, Z => n40301);
   U35667 : CLKBUF_X1 port map( A => n40302, Z => n40308);
   U35668 : CLKBUF_X1 port map( A => n40309, Z => n40315);
   U35669 : CLKBUF_X1 port map( A => n33323, Z => n40321);
   U35670 : CLKBUF_X1 port map( A => n40322, Z => n40328);
   U35671 : CLKBUF_X1 port map( A => n40329, Z => n40335);
   U35672 : CLKBUF_X1 port map( A => n33320, Z => n40341);
   U35673 : CLKBUF_X1 port map( A => n40342, Z => n40348);
   U35674 : CLKBUF_X1 port map( A => n40349, Z => n40355);
   U35675 : CLKBUF_X1 port map( A => n33317, Z => n40361);
   U35676 : CLKBUF_X1 port map( A => n40362, Z => n40368);
   U35677 : CLKBUF_X1 port map( A => n40369, Z => n40375);
   U35678 : CLKBUF_X1 port map( A => n33314, Z => n40381);
   U35679 : CLKBUF_X1 port map( A => n40382, Z => n40388);
   U35680 : CLKBUF_X1 port map( A => n40389, Z => n40395);
   U35681 : CLKBUF_X1 port map( A => n33311, Z => n40401);
   U35682 : CLKBUF_X1 port map( A => n40402, Z => n40408);
   U35683 : CLKBUF_X1 port map( A => n40409, Z => n40415);
   U35684 : CLKBUF_X1 port map( A => n33304, Z => n40421);
   U35685 : CLKBUF_X1 port map( A => n40422, Z => n40428);
   U35686 : CLKBUF_X1 port map( A => n40429, Z => n40435);
   U35687 : CLKBUF_X1 port map( A => n33293, Z => n40441);
   U35688 : CLKBUF_X1 port map( A => n40442, Z => n40448);
   U35689 : CLKBUF_X1 port map( A => n40449, Z => n40455);
   U35690 : CLKBUF_X1 port map( A => n33288, Z => n40461);
   U35691 : CLKBUF_X1 port map( A => n40462, Z => n40468);
   U35692 : CLKBUF_X1 port map( A => n40469, Z => n40475);
   U35693 : CLKBUF_X1 port map( A => n33283, Z => n40481);
   U35694 : CLKBUF_X1 port map( A => n40482, Z => n40488);
   U35695 : CLKBUF_X1 port map( A => n40489, Z => n40495);
   U35696 : CLKBUF_X1 port map( A => n33278, Z => n40501);
   U35697 : CLKBUF_X1 port map( A => n40502, Z => n40508);
   U35698 : CLKBUF_X1 port map( A => n40509, Z => n40515);
   U35699 : CLKBUF_X1 port map( A => n33273, Z => n40521);
   U35700 : CLKBUF_X1 port map( A => n40522, Z => n40528);
   U35701 : CLKBUF_X1 port map( A => n40529, Z => n40535);
   U35702 : CLKBUF_X1 port map( A => n33268, Z => n40541);
   U35703 : CLKBUF_X1 port map( A => n40542, Z => n40548);
   U35704 : CLKBUF_X1 port map( A => n40549, Z => n40555);
   U35705 : CLKBUF_X1 port map( A => n33263, Z => n40561);
   U35706 : CLKBUF_X1 port map( A => n40562, Z => n40568);
   U35707 : CLKBUF_X1 port map( A => n40569, Z => n40575);
   U35708 : CLKBUF_X1 port map( A => n33254, Z => n40581);
   U35709 : CLKBUF_X1 port map( A => n40582, Z => n40588);
   U35710 : CLKBUF_X1 port map( A => n40589, Z => n40595);

end SYN_bhv;
